.model nch_ss_1 nmos (
+ level = 54
+ fprout = 300
+ xrcrg1 = 12
+ xrcrg2 = 1
+ ags = 0.9375
+ wtvoff = 0
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ tvoff = 0.0019109629
+ keta = -0.06
+ cjd = 0.00145199
+ cit = 0.0001
+ cjs = 0.00145199
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 9.8024918e-9
+ xjbvd = 1
+ k3b = 1.9326
+ xjbvs = 1
+ lk2we = -1.5e-12
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ tvfbsdoff = 0.022
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 4e-12
+ capmod = 2
+ la0 = 0
+ kt1l = 0
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = 0.0004
+ kt1 = -0.200226
+ kt2 = -0.05325
+ wku0we = 2e-11
+ wkvth0we = 2e-12
+ llc = 0
+ ku0we = -0.0007
+ lln = 1
+ lu0 = -6e-12
+ mjd = 0.26
+ mjs = 0.26
+ beta0 = 13
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ leta0 = 0
+ njs = 1.02
+ pa0 = 0
+ mobmod = 0
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 6e-11
+ pbs = 0.52
+ lint = 6.5375218e-9
+ trnqsmod = 0
+ pu0 = 0
+ prt = 0
+ pud = 0
+ lkt1 = 0
+ lmax = 2.001e-5
+ lmin = 8.99743e-6
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 1.2299687e-9
+ ub1 = -7.2455506e-19
+ uc1 = 3.028e-11
+ dlcig = 2.5e-9
+ tpb = 0.0014
+ lpe0 = 9.2e-8
+ njtsswg = 9
+ bgidl = 2320000000.0
+ lpeb = 2.5e-7
+ wa0 = 0
+ ute = -1.007
+ wat = 0
+ web = 6843.8
+ wec = -25529.0
+ wlc = 0
+ wln = 1
+ wu0 = 2e-11
+ xgl = -1.09e-8
+ xgw = 0
+ wud = 0
+ wwc = 0
+ minv = -0.3
+ wwl = 0
+ wwn = 1
+ xtsswgd = 0.18
+ wvfbsdoff = 0
+ xtsswgs = 0.18
+ lvfbsdoff = 0
+ lub1 = 0
+ ndep = 1e+18
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.018555248
+ lwlc = 0
+ rgatemod = 0
+ dmcgt = 0
+ pdiblcb = -0.3
+ moin = 5.1
+ tcjsw = 0.000357
+ tnjtsswg = 1
+ nigc = 3.083
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ bigsd = 0.00125
+ bigbacc = 0.002588
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ wvoff = 0
+ ntox = -0.31099999999999994
+ pcit = 0
+ kvth0we = 0.00018
+ pclm = 1.4
+ wvsat = 0
+ wvth0 = 2.6e-9
+ lintnoi = -1.5e-8
+ bigbinv = 0.004953
+ phin = 0.15
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ pkt1 = 0
+ a0 = 3.25
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 72000
+ cf = 7.5795e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.026601253999999998
+ k3 = -1.8419
+ em = 1000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.01607
+ w0 = 0
+ ua = -1.8237726e-9
+ ub = 2.103696e-18
+ xpart = 1
+ uc = 7.33e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 5.6700000000000005e-9
+ ww = 0
+ xw = 3.4e-9
+ toxref = 3e-9
+ rbdb = 50
+ prwb = 0
+ prwg = 0
+ pub1 = 0
+ egidl = 0.29734
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ rdsw = 100
+ ijthsfwd = 0.01
+ ltvoff = 0
+ nfactor = 1
+ rshg = 15.6
+ ijthsrev = 0.01
+ pvoff = -7e-17
+ lku0we = 2.5e-11
+ cdscb = 0
+ cdscd = 0
+ epsrox = 3.9
+ pvsat = 0
+ wk2we = 5e-12
+ pvth0 = 2.3e-16
+ drout = 0.56
+ nigbacc = 10
+ rdsmod = 0
+ igbmod = 1
+ voffl = 0
+ tnom = 25
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ toxe = 2.47e-9
+ toxm = 2.43e-9
+ weta0 = 0
+ pbswgd = 0.95
+ pbswgs = 0.95
+ nigbinv = 10
+ igcmod = 1
+ cgidl = 0.22
+ wags = 1e-8
+ wcit = 0
+ voff = -0.1128204
+ fnoimod = 1
+ pbswd = 0.8
+ pbsws = 0.8
+ acde = 0.4
+ pkvth0we = -1.3e-19
+ eigbinv = 1.1
+ vsat = 102860
+ wint = 0
+ vth0 = 0.37711089000000003
+ wkt1 = 1.2e-9
+ pvfbsdoff = 0
+ wmax = 0.00090001
+ aigc = 0.011769394
+ wmin = 9.0026e-6
+ pdits = 0
+ vfbsdoff = 0.02
+ permod = 1
+ cigsd = 0.069865
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ bigc = 0.001442
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ paramchk = 1
+ wwlc = 0
+ cigbacc = 0.32875
+ voffcv = -0.16942
+ wpemod = 1
+ cdsc = 0
+ tnoia = 0
+ tnoimod = 0
+ cgbo = 0
+ cgdl = 3.0874977e-12
+ cgdo = 4.5622265999999996e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.0874977e-12
+ cgso = 4.5622265999999996e-11
+ cigc = 0.000625
+ peta0 = 0
+ cigbinv = 0.006
+ tpbsw = 0.0019
+ ijthdfwd = 0.01
+ cjswd = 8.774000000000001e-11
+ cjsws = 8.774000000000001e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ version = 4.5
+ tempmod = 0
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ tpbswg = 0.0009
+ ijthdrev = 0.01
+ aigbacc = 0.02
+ k2we = 5e-5
+ dsub = 0.75
+ dtox = 2.7e-10
+ scref = 1e-6
+ ptvoff = 0
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ pigcd = 2.621
+ aigsd = 0.01077322
+ lvoff = 0
+ eta0 = 0.3
+ aigbinv = 0.0163
+ diomod = 1
+ etab = -0.25
+ wtvfbsdoff = 0
+ lvsat = 0.0003
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 3.0174000000000004e-10
+ pku0we = -1.5e-18
+ lvth0 = 0
+ cjswgs = 3.0174000000000004e-10
+ lkvth0we = -2e-12
+ delta = 0.007595625
+ ltvfbsdoff = 0
+ rnoia = 0
+ rnoib = 0
+ mjswgd = 0.85
+ mjswgs = 0.85
+ acnqsmod = 0
+ ngate = 8e+20
+ tcjswg = 0.001
+ ngcon = 1
+ poxedge = 1
+ rbodymod = 0
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ binunit = 2
+ ptvfbsdoff = 0
+ )

.model nch_ss_2 nmos (
+ level = 54
+ wtvoff = 0
+ cgidl = 0.22
+ ijthdfwd = 0.01
+ capmod = 2
+ pbswd = 0.8
+ pbsws = 0.8
+ wku0we = 2e-11
+ rshg = 15.6
+ cigbacc = 0.32875
+ mobmod = 0
+ pvfbsdoff = 0
+ ijthdrev = 0.01
+ tnoimod = 0
+ pdits = 0
+ lpdiblc2 = -5.8501673e-10
+ cigsd = 0.069865
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ cigbinv = 0.006
+ tnom = 25
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ toxe = 2.47e-9
+ toxm = 2.43e-9
+ version = 4.5
+ tnoia = 0
+ tempmod = 0
+ lkvth0we = -2e-12
+ peta0 = 0
+ tpbsw = 0.0019
+ aigbacc = 0.02
+ wags = 1e-8
+ cjswd = 8.774000000000001e-11
+ cjsws = 8.774000000000001e-11
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ wcit = 0
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ acnqsmod = 0
+ voff = -0.11120139
+ acde = 0.4
+ vsat = 102860
+ wint = 0
+ rbodymod = 0
+ aigbinv = 0.0163
+ vth0 = 0.37136703000000004
+ wkt1 = 1.2e-9
+ wmax = 0.00090001
+ aigc = 0.01178613
+ wmin = 9.0026e-6
+ scref = 1e-6
+ pigcd = 2.621
+ toxref = 3e-9
+ aigsd = 0.01077322
+ bigc = 0.001442
+ wwlc = 0
+ lvoff = -1.4554874e-8
+ poxedge = 1
+ cdsc = 0
+ lvsat = 0.0003
+ cgbo = 0
+ cgdl = 3.0874977e-12
+ cgdo = 4.5622265999999996e-11
+ xtid = 3
+ xtis = 3
+ lvth0 = 5.1637332e-8
+ cgsl = 3.0874977e-12
+ cgso = 4.5622265999999996e-11
+ cigc = 0.000625
+ delta = 0.007595625
+ binunit = 2
+ laigc = -1.5044982e-10
+ rnoia = 0
+ rnoib = 0
+ ltvoff = -1.4627394e-10
+ a0 = 3.4752469
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ ngate = 8e+20
+ at = 61592.494
+ cf = 7.5795e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.028088843000000002
+ k3 = -1.8419
+ em = 1000000.0
+ ngcon = 1
+ ll = 0
+ lw = 0
+ u0 = 0.016291951000000002
+ w0 = 0
+ ua = -1.7995884e-9
+ ub = 2.1046515e-18
+ uc = 7.3387901e-11
+ ud = 0
+ wkvth0we = 2e-12
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 5.6700000000000005e-9
+ ww = 0
+ xw = 3.4e-9
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ lku0we = 2.5e-11
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ trnqsmod = 0
+ epsrox = 3.9
+ k2we = 5e-5
+ rdsmod = 0
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ dsub = 0.75
+ dtox = 2.7e-10
+ igbmod = 1
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ ags = 0.94104901
+ pbswgd = 0.95
+ pbswgs = 0.95
+ eta0 = 0.3
+ cjd = 0.00145199
+ rgatemod = 0
+ etab = -0.25
+ cit = -2.3830864e-5
+ cjs = 0.00145199
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 9.8024918e-9
+ tnjtsswg = 1
+ k3b = 1.9326
+ igcmod = 1
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ tvoff = 0.0019272336
+ la0 = -2.0249698e-6
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = 0.093963481
+ kt1 = -0.19577666
+ lk2 = -1.337342e-8
+ kt2 = -0.051823539
+ xjbvd = 1
+ llc = 0
+ xjbvs = 1
+ lln = 1
+ tvfbsdoff = 0.022
+ lk2we = -1.5e-12
+ lu0 = -2.0013361e-9
+ mjd = 0.26
+ lua = -2.1741579e-16
+ mjs = 0.26
+ lub = -8.5898229e-27
+ luc = -7.902321e-19
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njtsswg = 9
+ njd = 1.02
+ njs = 1.02
+ pa0 = 0
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 6e-11
+ pbs = 0.52
+ pu0 = 0
+ xtsswgd = 0.18
+ prt = 0
+ pud = 0
+ xtsswgs = 0.18
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 1.2713861e-9
+ ub1 = -7.4616446e-19
+ ku0we = -0.0007
+ uc1 = 2.5703642e-11
+ ckappad = 0.6
+ ckappas = 0.6
+ beta0 = 13
+ tpb = 0.0014
+ wa0 = 0
+ leta0 = 0
+ pdiblc1 = 0
+ pdiblc2 = 0.018620322
+ pdiblcb = -0.3
+ ute = -1.0077691
+ wat = 0
+ web = 6843.8
+ wec = -25529.0
+ wlc = 0
+ wln = 1
+ wu0 = 2e-11
+ xgl = -1.09e-8
+ xgw = 0
+ permod = 1
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ bigbacc = 0.002588
+ voffcv = -0.16942
+ wpemod = 1
+ dmcgt = 0
+ tcjsw = 0.000357
+ kvth0we = 0.00018
+ lintnoi = -1.5e-8
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ keta = -0.059896633
+ ijthsfwd = 0.01
+ bigsd = 0.00125
+ lags = -3.1905621e-8
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 1.1172395e-9
+ wvoff = 0
+ kt1l = 0
+ tpbswg = 0.0009
+ wvsat = 0
+ wvth0 = 2.6e-9
+ ijthsrev = 0.01
+ lint = 6.5375218e-9
+ lkt1 = -3.9999573e-8
+ lkt2 = -1.2823887e-8
+ wtvfbsdoff = 0
+ lmax = 8.99743e-6
+ lmin = 8.974099999999999e-7
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ ptvoff = 0
+ lketa = -9.2926692e-10
+ xpart = 1
+ ltvfbsdoff = 0
+ minv = -0.3
+ lua1 = -3.7234224e-16
+ lub1 = 1.9426851e-25
+ luc1 = 4.1141459e-17
+ nfactor = 1
+ diomod = 1
+ ndep = 1e+18
+ lute = 6.9145309e-9
+ egidl = 0.29734
+ lwlc = 0
+ moin = 5.1
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 3.0174000000000004e-10
+ pku0we = -1.5e-18
+ cjswgs = 3.0174000000000004e-10
+ nigc = 3.083
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ mjswgd = 0.85
+ mjswgs = 0.85
+ nigbacc = 10
+ ptvfbsdoff = 0
+ tcjswg = 0.001
+ ntox = -0.31099999999999994
+ pkvth0we = -1.3e-19
+ pcit = 0
+ pclm = 1.4
+ pvoff = -7e-17
+ nigbinv = 10
+ phin = 0.15
+ cdscb = 0
+ cdscd = 0
+ vfbsdoff = 0.02
+ pvsat = 0
+ wk2we = 5e-12
+ pkt1 = 0
+ pvth0 = 2.3e-16
+ drout = 0.56
+ voffl = 0
+ fprout = 300
+ paramchk = 1
+ rbdb = 50
+ prwb = 0
+ prwg = 0
+ pub1 = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ fnoimod = 1
+ weta0 = 0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ eigbinv = 1.1
+ rdsw = 100
+ )

.model nch_ss_3 nmos (
+ level = 54
+ ku0we = -0.0007
+ beta0 = 13
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ leta0 = 0
+ ijthsrev = 0.01
+ kvth0we = 0.00018
+ lintnoi = -1.5e-8
+ k2we = 5e-5
+ bigbinv = 0.004953
+ dlcig = 2.5e-9
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ bgidl = 2320000000.0
+ dsub = 0.75
+ wvfbsdoff = 0
+ dtox = 2.7e-10
+ lvfbsdoff = 0
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ eta0 = 0.3
+ dmcgt = 0
+ etab = -0.25
+ tcjsw = 0.000357
+ bigsd = 0.00125
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ wvoff = 0
+ pkvth0we = -1.3e-19
+ nfactor = 1
+ wvsat = 0
+ wvth0 = 2.6e-9
+ vfbsdoff = 0.02
+ lketa = -2.6515603e-8
+ toxref = 3e-9
+ xpart = 1
+ nigbacc = 10
+ paramchk = 1
+ egidl = 0.29734
+ nigbinv = 10
+ keta = -0.031147941
+ ltvoff = -6.4393769e-10
+ ijthdfwd = 0.01
+ lags = 4.0889306e-7
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = -1.0651822e-10
+ kt1l = 0
+ lku0we = 2.5e-11
+ fnoimod = 1
+ ijthdrev = 0.01
+ epsrox = 3.9
+ eigbinv = 1.1
+ pvoff = -7e-17
+ lint = 6.5375218e-9
+ cdscb = 0
+ cdscd = 0
+ lkt1 = -1.7764368e-8
+ lkt2 = -1.1493547e-8
+ lmax = 8.974099999999999e-7
+ lpdiblc2 = 3.0380287e-9
+ pvsat = 0
+ lmin = 4.4741e-7
+ rdsmod = 0
+ wk2we = 5e-12
+ pvth0 = 2.3e-16
+ drout = 0.56
+ igbmod = 1
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ minv = -0.3
+ voffl = 0
+ lua1 = -1.0281867e-16
+ lub1 = 1.8552992e-26
+ luc1 = 3.7680622e-18
+ pbswgd = 0.95
+ pbswgs = 0.95
+ ndep = 1e+18
+ weta0 = 0
+ lwlc = 0
+ igcmod = 1
+ moin = 5.1
+ a0 = 1.288
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ cigbacc = 0.32875
+ at = 219598.22
+ cf = 7.5795e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.027010322000000003
+ k3 = -1.8419
+ em = 1000000.0
+ ll = 0
+ nigc = 3.083
+ lw = 0
+ u0 = 0.015790444
+ w0 = 0
+ ua = -1.9429424e-9
+ ub = 2.1566e-18
+ uc = 9.3717778e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 5.6700000000000005e-9
+ ww = 0
+ xw = 3.4e-9
+ lkvth0we = -2e-12
+ cgidl = 0.22
+ tnoimod = 0
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ cigbinv = 0.006
+ acnqsmod = 0
+ pbswd = 0.8
+ pbsws = 0.8
+ ntox = -0.31099999999999994
+ pcit = 0
+ pclm = 1.4
+ pvfbsdoff = 0
+ rbodymod = 0
+ version = 4.5
+ permod = 1
+ phin = 0.15
+ tempmod = 0
+ pdits = 0
+ cigsd = 0.069865
+ pkt1 = 0
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ aigbacc = 0.02
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ voffcv = -0.16942
+ wpemod = 1
+ rbdb = 50
+ prwb = 0
+ pub1 = 0
+ prwg = 0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ tnoia = 0
+ rdsw = 100
+ aigbinv = 0.0163
+ peta0 = 0
+ tpbsw = 0.0019
+ wtvfbsdoff = 0
+ cjswd = 8.774000000000001e-11
+ cjsws = 8.774000000000001e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ tpbswg = 0.0009
+ rshg = 15.6
+ ltvfbsdoff = 0
+ wkvth0we = 2e-12
+ poxedge = 1
+ trnqsmod = 0
+ ptvoff = 0
+ binunit = 2
+ scref = 1e-6
+ pigcd = 2.621
+ aigsd = 0.01077322
+ tnom = 25
+ diomod = 1
+ toxe = 2.47e-9
+ toxm = 2.43e-9
+ ptvfbsdoff = 0
+ lvoff = -1.3768912e-8
+ pditsd = 0
+ rgatemod = 0
+ pditsl = 0
+ cjswgd = 3.0174000000000004e-10
+ pku0we = -1.5e-18
+ cjswgs = 3.0174000000000004e-10
+ tnjtsswg = 1
+ lvsat = 0.0003
+ lvth0 = 7.4115504e-9
+ delta = 0.007595625
+ laigc = -5.5724245e-11
+ rnoia = 0
+ rnoib = 0
+ mjswgd = 0.85
+ mjswgs = 0.85
+ wags = 1e-8
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ wcit = 0
+ tcjswg = 0.001
+ ngate = 8e+20
+ voff = -0.1120845
+ acde = 0.4
+ ngcon = 1
+ vsat = 102860
+ wint = 0
+ vth0 = 0.42105892
+ gbmin = 1e-12
+ wkt1 = 1.2e-9
+ jswgd = 1.28e-13
+ wmax = 0.00090001
+ jswgs = 1.28e-13
+ aigc = 0.011679696
+ wmin = 9.0026e-6
+ ags = 0.4457696
+ cjd = 0.00145199
+ cit = 0.0013511778
+ cjs = 0.00145199
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 9.8024918e-9
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ fprout = 300
+ dwg = 0
+ dwj = 0
+ njtsswg = 9
+ bigc = 0.001442
+ xrcrg1 = 12
+ xrcrg2 = 1
+ wwlc = 0
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ la0 = -7.832e-8
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.046661618
+ kt1 = -0.22076004
+ kt2 = -0.053318302
+ lk2 = -1.2413537e-8
+ llc = 0
+ cdsc = 0
+ lln = 1
+ lu0 = -1.5549956e-9
+ ckappad = 0.6
+ ckappas = 0.6
+ mjd = 0.26
+ mjs = 0.26
+ lua = -8.9830708e-17
+ lub = -5.4824e-26
+ luc = -1.8883822e-17
+ lud = 0
+ lwc = 0
+ cgbo = 0
+ wtvoff = 0
+ lwl = 0
+ lwn = 1
+ cgdl = 3.0874977e-12
+ cgdo = 4.5622265999999996e-11
+ xtid = 3
+ pdiblc1 = 0
+ pdiblc2 = 0.014549485
+ njd = 1.02
+ xtis = 3
+ njs = 1.02
+ pa0 = 0
+ pdiblcb = -0.3
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 6e-11
+ pbs = 0.52
+ cgsl = 3.0874977e-12
+ cgso = 4.5622265999999996e-11
+ cigc = 0.000625
+ pu0 = 0
+ tvoff = 0.0024864064
+ prt = 0
+ pud = 0
+ tvfbsdoff = 0.022
+ rsh = 17.5
+ tcj = 0.00076
+ ijthsfwd = 0.01
+ xjbvd = 1
+ ua1 = 9.685506e-10
+ ub1 = -5.4873129e-19
+ xjbvs = 1
+ uc1 = 6.7696222e-11
+ lk2we = -1.5e-12
+ tpb = 0.0014
+ capmod = 2
+ wa0 = 0
+ ute = -1
+ wat = 0
+ web = 6843.8
+ wec = -25529.0
+ wlc = 0
+ wln = 1
+ wku0we = 2e-11
+ wu0 = 2e-11
+ xgl = -1.09e-8
+ xgw = 0
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ bigbacc = 0.002588
+ mobmod = 0
+ )

.model nch_ss_4 nmos (
+ level = 54
+ minv = -0.3
+ lua1 = -3.0475764e-17
+ pk2we = -1e-19
+ lub1 = -2.9971927e-26
+ luc1 = -4.3987511e-18
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ ndep = 1e+18
+ rgatemod = 0
+ lwlc = 0
+ moin = 5.1
+ tnjtsswg = 1
+ tnoia = 0
+ nigc = 3.083
+ peta0 = 0
+ poxedge = 1
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ tpbsw = 0.0019
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ binunit = 2
+ cjswd = 8.774000000000001e-11
+ cjsws = 8.774000000000001e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ ntox = -0.31099999999999994
+ pcit = 0
+ pclm = 1.5439223
+ phin = 0.15
+ pkt1 = 0
+ toxref = 3e-9
+ scref = 1e-6
+ jtsswgd = 2.3e-7
+ pigcd = 2.621
+ jtsswgs = 2.3e-7
+ aigsd = 0.01077322
+ rbdb = 50
+ prwb = 0
+ pub1 = 0
+ prwg = 0
+ lvoff = -6.3216134e-9
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ rdsw = 100
+ lvsat = 0.0003
+ lvth0 = -4.690878e-9
+ delta = 0.007595625
+ ltvoff = -1.206053e-10
+ laigc = -1.9935708e-11
+ rnoia = 0
+ rnoib = 0
+ ijthsfwd = 0.01
+ ngate = 8e+20
+ njtsswg = 9
+ ngcon = 1
+ rshg = 15.6
+ lku0we = 2.5e-11
+ ags = 0.124315598
+ epsrox = 3.9
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ cjd = 0.00145199
+ cit = 0.00073144105
+ ijthsrev = 0.01
+ cjs = 0.00145199
+ clc = 1e-7
+ cle = 0.6
+ gbmin = 1e-12
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 1.30529375e-8
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ k3b = 1.9326
+ ckappad = 0.6
+ ckappas = 0.6
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ rdsmod = 0
+ pdiblc1 = 0
+ pdiblc2 = 0.027331777
+ pdiblcb = -0.3
+ igbmod = 1
+ la0 = -2.4730306e-7
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.016465258
+ kt1 = -0.23920434
+ kt2 = -0.070668297
+ lk2 = -9.6174482e-9
+ llc = -1.18e-13
+ lln = 0.7
+ lu0 = -6.303388699999999e-10
+ mjd = 0.26
+ mjs = 0.26
+ lua = -1.0757894e-17
+ lub = -4.7838952e-26
+ luc = -6.6488035e-18
+ lud = 0
+ pbswgd = 0.95
+ pbswgs = 0.95
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ tnom = 25
+ njd = 1.02
+ njs = 1.02
+ pa0 = 0
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 6e-11
+ pbs = 0.52
+ toxe = 2.47e-9
+ toxm = 2.43e-9
+ pu0 = 0
+ igcmod = 1
+ prt = 0
+ pud = 0
+ bigbacc = 0.002588
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 8.041349e-10
+ ub1 = -4.3844738e-19
+ uc1 = 8.6257162e-11
+ tpb = 0.0014
+ wa0 = 0
+ ute = -1
+ wat = 0
+ web = 6843.8
+ wec = -25529.0
+ kvth0we = 0.00018
+ wlc = 0
+ wln = 1
+ wu0 = 2e-11
+ xgl = -1.09e-8
+ xgw = 0
+ tvoff = 0.0012970146
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ tvfbsdoff = 0.022
+ lintnoi = -1.5e-8
+ xjbvd = 1
+ xjbvs = 1
+ wags = 1e-8
+ lk2we = -1.5e-12
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ wcit = 0
+ voff = -0.12901018
+ acde = 0.4
+ pkvth0we = -1.3e-19
+ ku0we = -0.0007
+ beta0 = 13
+ vsat = 102860
+ wint = 0
+ permod = 1
+ leta0 = 0
+ vth0 = 0.44856443
+ wkt1 = 1.2e-9
+ wmax = 0.00090001
+ aigc = 0.011598359
+ wmin = 9.0026e-6
+ vfbsdoff = 0.02
+ a0 = 1.6720524
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 150970.13
+ cf = 7.5795e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.020655575000000002
+ k3 = -1.8419
+ em = 1000000.0
+ dlcig = 2.5e-9
+ ll = -1.18e-13
+ wvfbsdoff = 0
+ lw = 0
+ u0 = 0.013688951999999999
+ bgidl = 2320000000.0
+ w0 = 0
+ lvfbsdoff = 0
+ ua = -2.1226533e-9
+ ub = 2.1407249e-18
+ uc = 6.5910917e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 5.6700000000000005e-9
+ ww = 0
+ xw = 3.4e-9
+ voffcv = -0.16942
+ wpemod = 1
+ bigc = 0.001442
+ paramchk = 1
+ wwlc = 0
+ wtvfbsdoff = 0
+ dmcgt = 0
+ tcjsw = 0.000357
+ nfactor = 1
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.0874977e-12
+ cgdo = 4.5622265999999996e-11
+ xtid = 3
+ xtis = 3
+ ltvfbsdoff = 0
+ cgsl = 3.0874977e-12
+ cgso = 4.5622265999999996e-11
+ cigc = 0.000625
+ ijthdfwd = 0.01
+ bigsd = 0.00125
+ tpbswg = 0.0009
+ wvoff = 0
+ nigbacc = 10
+ wvsat = 0
+ wvth0 = 2.6e-9
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ ijthdrev = 0.01
+ ptvfbsdoff = 0
+ lpdiblc2 = -2.58618e-9
+ ptvoff = 0
+ nigbinv = 10
+ k2we = 5e-5
+ dsub = 0.75
+ lketa = -2.2644187e-8
+ dtox = 2.7e-10
+ xpart = 1
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ diomod = 1
+ pditsd = 0
+ pditsl = 0
+ egidl = 0.29734
+ cjswgd = 3.0174000000000004e-10
+ pku0we = -1.5e-18
+ cjswgs = 3.0174000000000004e-10
+ eta0 = 0.3
+ etab = -0.25
+ fnoimod = 1
+ eigbinv = 1.1
+ lkvth0we = -2e-12
+ mjswgd = 0.85
+ mjswgs = 0.85
+ tcjswg = 0.001
+ acnqsmod = 0
+ rbodymod = 0
+ pvoff = -7e-17
+ cigbacc = 0.32875
+ cdscb = 0
+ cdscd = 0
+ pvsat = 0
+ wk2we = 5e-12
+ pvth0 = 2.3e-16
+ drout = 0.56
+ tnoimod = 0
+ fprout = 300
+ voffl = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ cigbinv = 0.006
+ weta0 = 0
+ lpclm = -6.3325799e-8
+ wtvoff = 0
+ version = 4.5
+ cgidl = 0.22
+ tempmod = 0
+ keta = -0.039946614
+ capmod = 2
+ lags = 5.5033282e-7
+ wku0we = 2e-11
+ aigbacc = 0.02
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 1.6616594000000001e-10
+ pbswd = 0.8
+ mobmod = 0
+ pbsws = 0.8
+ kt1l = 0
+ wkvth0we = 2e-12
+ pvfbsdoff = 0
+ lint = 9.7879675e-9
+ trnqsmod = 0
+ pdits = 0
+ lkt1 = -9.6488734e-9
+ lkt2 = -3.8595493e-9
+ aigbinv = 0.0163
+ lmax = 4.4741e-7
+ cigsd = 0.069865
+ lmin = 2.1410000000000002e-7
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ laigsd = -8.1082969e-17
+ )

.model nch_ss_5 nmos (
+ level = 54
+ nigbinv = 10
+ bigsd = 0.00125
+ wags = 1e-8
+ wcit = 0
+ acnqsmod = 0
+ wvoff = 0
+ voff = -0.15746310460000001
+ acde = 0.4
+ wvsat = 0
+ vsat = 102521.2852
+ wvth0 = 2.6e-9
+ rbodymod = 0
+ wint = 0
+ vth0 = 0.46456137420000004
+ wkt1 = 1.2e-9
+ wmax = 0.00090001
+ aigc = 0.011526753
+ wmin = 9.0026e-6
+ fnoimod = 1
+ eigbinv = 1.1
+ toxref = 3e-9
+ lketa = -1.1430034e-8
+ xpart = 1
+ bigc = 0.001442
+ wwlc = 0
+ egidl = 0.29734
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.0874977e-12
+ cgdo = 4.5622265999999996e-11
+ xtid = 3
+ xtis = 3
+ ltvoff = 1.4850105e-11
+ cgsl = 3.0874977e-12
+ cgso = 4.5622265999999996e-11
+ cigc = 0.000625
+ cigbacc = 0.32875
+ tnoimod = 0
+ lku0we = 2.5e-11
+ cigbinv = 0.006
+ epsrox = 3.9
+ wkvth0we = 2e-12
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ pvoff = -7e-17
+ rdsmod = 0
+ trnqsmod = 0
+ cdscb = 0
+ cdscd = 0
+ igbmod = 1
+ pvsat = 0
+ version = 4.5
+ wk2we = 5e-12
+ pvth0 = 2.3e-16
+ k2we = 5e-5
+ drout = 0.56
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ tempmod = 0
+ dsub = 0.75
+ dtox = 2.7e-10
+ pbswgd = 0.95
+ pbswgs = 0.95
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ voffl = 0
+ igcmod = 1
+ aigbacc = 0.02
+ weta0 = 0
+ eta0 = 0.3
+ rgatemod = 0
+ etab = -0.25
+ lpclm = -2.4377173e-8
+ tnjtsswg = 1
+ cgidl = 0.22
+ aigbinv = 0.0163
+ pbswd = 0.8
+ pbsws = 0.8
+ pvfbsdoff = 0
+ permod = 1
+ wtvfbsdoff = 0
+ pdits = 0
+ cigsd = 0.069865
+ dvt0w = 0
+ dvt1w = 0
+ poxedge = 1
+ dvt2w = 0
+ ltvfbsdoff = 0
+ voffcv = -0.16942
+ wpemod = 1
+ binunit = 2
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ tnoia = 0
+ peta0 = 0
+ wketa = 0
+ keta = -0.093093889
+ ptvfbsdoff = 0
+ tpbsw = 0.0019
+ ijthsfwd = 0.01
+ cjswd = 8.774000000000001e-11
+ cjsws = 8.774000000000001e-11
+ a0 = 0.66068814
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ mjswd = 0.11
+ lags = 3.3904274e-13
+ mjsws = 0.11
+ agidl = 9.41e-8
+ tpbswg = 0.0009
+ at = 79499.116
+ cf = 7.5795e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = -0.014112077999999998
+ k3 = -1.8419
+ em = 1000000.0
+ jswd = 1.28e-13
+ ll = -1.18e-13
+ jsws = 1.28e-13
+ lw = 0
+ u0 = 0.011686872
+ w0 = 0
+ lcit = 8.8591162e-11
+ ua = -2.2893587e-9
+ ub = 2.089788886e-18
+ uc = 4.5969231e-11
+ ud = 0
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 5.6700000000000005e-9
+ ww = 0
+ xw = 3.4e-9
+ kt1l = 0
+ ijthsrev = 0.01
+ lint = 9.7879675e-9
+ ptvoff = 0
+ lkt1 = -3.3075226e-9
+ lkt2 = -6.0180086e-10
+ lmax = 2.1410000000000002e-7
+ lmin = 8.833e-8
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ scref = 1e-6
+ diomod = 1
+ pigcd = 2.621
+ minv = -0.3
+ aigsd = 0.01077322
+ lua1 = 7.6861327e-18
+ lub1 = -5.2342256e-26
+ luc1 = -4.2210821e-18
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 3.0174000000000004e-10
+ pku0we = -1.5e-18
+ cjswgs = 3.0174000000000004e-10
+ ndep = 1e+18
+ lvoff = -3.1806260000000004e-10
+ njtsswg = 9
+ lwlc = 0
+ moin = 5.1
+ lvsat = 0.00037148429999999994
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ lvth0 = -8.0662159e-9
+ nigc = 3.083
+ delta = 0.007595625
+ mjswgd = 0.85
+ mjswgs = 0.85
+ laigc = -4.8268328e-12
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.02163037
+ pdiblcb = -0.3
+ tcjswg = 0.001
+ rnoia = 0
+ rnoib = 0
+ ags = 2.7325264
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ cjd = 0.00145199
+ cit = 0.001099094
+ cjs = 0.00145199
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 1.30529375e-8
+ pketa = 0
+ ngate = 8e+20
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ ngcon = 1
+ pkvth0we = -1.3e-19
+ ntox = -0.31099999999999994
+ pcit = 0
+ pclm = 1.3593316
+ bigbacc = 0.002588
+ la0 = -3.3904685e-8
+ gbmin = 1e-12
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.0013848735
+ kt1 = -0.26925814
+ kt2 = -0.086107863
+ lk2 = -2.2814734e-9
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ llc = -1.18e-13
+ lln = 0.7
+ phin = 0.15
+ lu0 = -2.0789995e-10
+ mjd = 0.26
+ mjs = 0.26
+ lua = 2.4416942e-17
+ lub = -3.7091512499999996e-26
+ luc = -2.4411077e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ vfbsdoff = 0.02
+ njd = 1.02
+ njs = 1.02
+ pa0 = 0
+ nsd = 1e+20
+ kvth0we = 0.00018
+ pbd = 0.52
+ pat = 6e-11
+ pbs = 0.52
+ pkt1 = 0
+ pu0 = 0
+ prt = 0
+ fprout = 300
+ pub = 0
+ pud = 0
+ lintnoi = -1.5e-8
+ rsh = 17.5
+ xrcrg1 = 12
+ xrcrg2 = 1
+ tcj = 0.00076
+ ua1 = 6.2327283e-10
+ ub1 = -3.3242687e-19
+ uc1 = 8.5415128e-11
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ tpb = 0.0014
+ wa0 = 0
+ ute = -1
+ paramchk = 1
+ wat = 0
+ web = 6843.8
+ wec = -25529.0
+ wlc = 0
+ wln = 1
+ wu0 = 2e-11
+ rbdb = 50
+ xgl = -1.09e-8
+ prwb = 0
+ pub1 = 0
+ prwg = 0
+ xgw = 0
+ wub = 0
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ rbpb = 50
+ rbpd = 50
+ wtvoff = 0
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ rdsw = 100
+ tvfbsdoff = 0.022
+ tvoff = 0.00065504585
+ capmod = 2
+ ijthdfwd = 0.01
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ wku0we = 2e-11
+ mobmod = 0
+ rshg = 15.6
+ ku0we = -0.0007
+ beta0 = 13
+ leta0 = 0
+ ijthdrev = 0.01
+ nfactor = 1
+ lpdiblc2 = -1.3831831e-9
+ wvfbsdoff = 0
+ dlcig = 2.5e-9
+ lvfbsdoff = 0
+ bgidl = 2320000000.0
+ laigsd = 3.3904273e-17
+ tnom = 25
+ toxe = 2.47e-9
+ toxm = 2.43e-9
+ nigbacc = 10
+ dmcgt = 0
+ tcjsw = 0.000357
+ lkvth0we = -2e-12
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ )

.model nch_ss_6 nmos (
+ level = 54
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ vfbsdoff = 0.02
+ toxref = 3e-9
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.0069155858
+ scref = 1e-6
+ pdiblcb = -0.3
+ pigcd = 2.621
+ aigsd = 0.01077322
+ paramchk = 1
+ lvoff = -2.06441089e-9
+ ags = 2.7325299999999997
+ lvsat = 0.0024722048699999995
+ ltvoff = 1.0839662e-10
+ lvth0 = 2.2492931699999996e-9
+ bigbacc = 0.002588
+ cjd = 0.00145199
+ cit = -3.6108899999999955e-6
+ cjs = 0.00145199
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ delta = 0.007595625
+ dlc = 3.26497e-9
+ k3b = 1.9326
+ laigc = -2.2427226e-11
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ keta = -0.52835722
+ rnoia = 0
+ rnoib = 0
+ ijthdfwd = 0.01
+ kvth0we = 0.00018
+ la0 = 3.0288889e-8
+ jsd = 6.11e-7
+ lintnoi = -1.5e-8
+ jss = 6.11e-7
+ lat = 1.9707860000000026e-5
+ kt1 = -0.40872879
+ kt2 = -0.10088778
+ lk2 = -4.8654938e-10
+ lku0we = 2.5e-11
+ pketa = 0
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ ngate = 8e+20
+ bigbinv = 0.004953
+ llc = 0
+ lln = 1
+ lu0 = 9.683078e-11
+ lcit = 1.9224546e-10
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ mjd = 0.26
+ mjs = 0.26
+ lua = 3.5218789e-17
+ lub = -1.9869262700000004e-26
+ luc = 2.2716666e-18
+ lud = 0
+ epsrox = 3.9
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ ngcon = 1
+ njd = 1.02
+ njs = 1.02
+ kt1l = 0
+ pa0 = 0
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 6e-11
+ pbs = 0.52
+ pu0 = 0.0
+ prt = 0
+ pub = 0
+ puc = 0
+ pud = 0
+ rdsmod = 0
+ ijthdrev = 0.01
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ rsh = 17.5
+ jswgs = 1.28e-13
+ lint = 0
+ tcj = 0.00076
+ igbmod = 1
+ ua1 = 8.897383e-10
+ ub1 = -8.0235504e-19
+ uc1 = -6.3390556e-11
+ tpb = 0.0014
+ lkt1 = 9.8027184e-9
+ lkt2 = 7.8751111e-10
+ wa0 = 0
+ lpdiblc2 = 6.6256944e-15
+ lmax = 8.833e-8
+ ute = -1
+ wat = 0
+ web = 6843.8
+ pscbe1 = 1000000000.0
+ wec = -25529.0
+ pscbe2 = 1e-20
+ lmin = 5.233e-8
+ wlc = 0
+ wln = 1
+ wu0 = 2e-11
+ xgl = -1.09e-8
+ xgw = 0
+ wub = 0
+ wuc = 0
+ wud = 0
+ lpe0 = 9.2e-8
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ pbswgd = 0.95
+ lpeb = 2.5e-7
+ pbswgs = 0.95
+ minv = -0.3
+ igcmod = 1
+ lua1 = -1.7361621e-17
+ lub1 = -8.1690078e-27
+ luc1 = 9.7666522e-18
+ ndep = 1e+18
+ lwlc = 0
+ moin = 5.1
+ nigc = 3.083
+ tvfbsdoff = 0.022
+ nfactor = 1
+ lkvth0we = -2e-12
+ tvoff = -0.00034012981
+ wtvfbsdoff = 0
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ acnqsmod = 0
+ ltvfbsdoff = 0
+ permod = 1
+ ntox = -0.31099999999999994
+ pcit = 0.0
+ ku0we = -0.0007
+ pclm = 1.2209944
+ beta0 = 13
+ rbodymod = 0
+ leta0 = 3.0288889e-9
+ nigbacc = 10
+ letab = -2.2684433e-8
+ phin = 0.15
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ pkt1 = 0
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ voffcv = -0.16942
+ wpemod = 1
+ nigbinv = 10
+ ptvfbsdoff = 0
+ rbdb = 50
+ prwb = 0
+ pub1 = 0
+ prwg = 0
+ dmcgt = 0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ tcjsw = 0.000357
+ rdsw = 100
+ fnoimod = 1
+ eigbinv = 1.1
+ bigsd = 0.00125
+ tpbswg = 0.0009
+ wvoff = 0
+ rshg = 15.6
+ wkvth0we = 2e-12
+ wvsat = 0.0
+ wvth0 = 2.6e-9
+ ptvoff = 0
+ trnqsmod = 0
+ cigbacc = 0.32875
+ diomod = 1
+ lketa = 2.9484719e-8
+ xpart = 1
+ pditsd = 0
+ pditsl = 0
+ tnoimod = 0
+ cjswgd = 3.0174000000000004e-10
+ pku0we = -1.5e-18
+ cjswgs = 3.0174000000000004e-10
+ tnom = 25
+ toxe = 2.47e-9
+ toxm = 2.43e-9
+ egidl = 0.29734
+ a0 = -0.02222221999999996
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ rgatemod = 0
+ at = 64556.761
+ cf = 7.5795e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = -0.033207015
+ k3 = -1.8419
+ em = 1000000.0
+ cigbinv = 0.006
+ ll = 0
+ lw = 0
+ u0 = 0.0084450556
+ tnjtsswg = 1
+ w0 = 0
+ ua = -2.404272e-9
+ ub = 1.906573466e-18
+ uc = -4.166667e-12
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 5.6700000000000005e-9
+ ww = 0
+ xw = 3.4e-9
+ mjswgd = 0.85
+ mjswgs = 0.85
+ tcjswg = 0.001
+ version = 4.5
+ wags = 1e-8
+ tempmod = 0
+ wcit = 0.0
+ voff = -0.138884931
+ acde = 0.4
+ aigbacc = 0.02
+ vsat = 80173.2
+ wint = 0
+ vth0 = 0.354821916
+ pvoff = -7e-17
+ wkt1 = 1.2e-9
+ wmax = 0.00090001
+ aigc = 0.011713991
+ wmin = 9.0026e-6
+ cdscb = 0
+ cdscd = 0
+ pvsat = 0.0
+ wk2we = 5e-12
+ pvth0 = 2.3e-16
+ fprout = 300
+ drout = 0.56
+ xrcrg1 = 12
+ xrcrg2 = 1
+ aigbinv = 0.0163
+ voffl = 0
+ bigc = 0.001442
+ wwlc = 0
+ wtvoff = 0
+ weta0 = 0
+ lpclm = -1.1373478e-8
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.0874977e-12
+ cgdo = 4.5622265999999996e-11
+ xtid = 3
+ xtis = 3
+ cgidl = 0.22
+ cgsl = 3.0874977e-12
+ cgso = 4.5622265999999996e-11
+ cigc = 0.000625
+ capmod = 2
+ wku0we = 2e-11
+ ijthsfwd = 0.01
+ poxedge = 1
+ mobmod = 0
+ pbswd = 0.8
+ pvfbsdoff = 0
+ pbsws = 0.8
+ binunit = 2
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ ijthsrev = 0.01
+ pdits = 0
+ cigsd = 0.069865
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ k2we = 5e-5
+ dsub = 0.75
+ dtox = 2.7e-10
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ eta0 = 0.26777778
+ etab = -0.0086762422
+ tnoia = 0
+ peta0 = 0
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ wketa = 0
+ tpbsw = 0.0019
+ cjswd = 8.774000000000001e-11
+ cjsws = 8.774000000000001e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ pkvth0we = -1.3e-19
+ njtsswg = 9
+ )

.model nch_ss_7 nmos (
+ level = 54
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ ltvoff = -2.4740506e-10
+ aigbacc = 0.02
+ rdsw = 100
+ ijthsfwd = 0.01
+ lku0we = 2.5e-11
+ aigbinv = 0.0163
+ epsrox = 3.9
+ rshg = 15.6
+ rdsmod = 0
+ igbmod = 1
+ ijthsrev = 0.01
+ pvoff = -7e-17
+ cdscb = 0
+ cdscd = 0
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ pvsat = 0.0
+ wk2we = 5e-12
+ pvth0 = 2.3e-16
+ drout = 0.56
+ pbswgd = 0.95
+ pbswgs = 0.95
+ igcmod = 1
+ poxedge = 1
+ wtvfbsdoff = 0
+ voffl = 0
+ tnom = 25
+ toxe = 2.47e-9
+ toxm = 2.43e-9
+ weta0 = 0
+ binunit = 2
+ lpclm = -7.2871722e-8
+ ltvfbsdoff = 0
+ cgidl = 0.22
+ wags = 1e-8
+ wcit = 0.0
+ pvfbsdoff = 0
+ permod = 1
+ pbswd = 0.8
+ pbsws = 0.8
+ voff = -0.112415764
+ pkvth0we = -1.3e-19
+ acde = 0.4
+ ptvfbsdoff = 0
+ vsat = 88037.262
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ wint = 0
+ vth0 = 0.35271759700000005
+ wkt1 = 1.2e-9
+ wmax = 0.00090001
+ aigc = 0.011692671
+ pdits = 0
+ wmin = 9.0026e-6
+ vfbsdoff = 0.02
+ cigsd = 0.069865
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ voffcv = -0.16942
+ wpemod = 1
+ wub1 = 0.0
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ bigc = 0.001442
+ paramchk = 1
+ wwlc = 0
+ tnoia = 0
+ cdsc = 0
+ cgbo = 0
+ njtsswg = 9
+ cgdl = 3.0874977e-12
+ cgdo = 4.5622265999999996e-11
+ xtid = 3
+ xtis = 3
+ peta0 = 0
+ cgsl = 3.0874977e-12
+ cgso = 4.5622265999999996e-11
+ cigc = 0.000625
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ tpbsw = 0.0019
+ ijthdfwd = 0.01
+ tpbswg = 0.0009
+ ckappad = 0.6
+ cjswd = 8.774000000000001e-11
+ ckappas = 0.6
+ cjsws = 8.774000000000001e-11
+ mjswd = 0.11
+ pdiblc1 = 0
+ pdiblc2 = 0.0069157
+ mjsws = 0.11
+ agidl = 9.41e-8
+ pdiblcb = -0.3
+ ptvoff = 0
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ ijthdrev = 0.01
+ bigbacc = 0.002588
+ diomod = 1
+ k2we = 5e-5
+ dsub = 0.75
+ scref = 1e-6
+ dtox = 2.7e-10
+ pditsd = 0
+ pditsl = 0
+ kvth0we = 0.00018
+ cjswgd = 3.0174000000000004e-10
+ pku0we = -1.5e-18
+ cjswgs = 3.0174000000000004e-10
+ ags = 2.7325299999999997
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ pigcd = 2.621
+ aigsd = 0.01077322
+ cjd = 0.00145199
+ cit = -0.0036312757
+ cjs = 0.00145199
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ lintnoi = -1.5e-8
+ dlc = 3.26497e-9
+ bigbinv = 0.004953
+ k3b = 1.9326
+ lvoff = -3.599622200000001e-9
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ eta0 = 0.35179556
+ etab = -1.0973583
+ lvsat = 0.0020160890999999996
+ mjswgd = 0.85
+ mjswgs = 0.85
+ lvth0 = 2.3713433000000004e-9
+ la0 = -3.1577778e-7
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = 0.009241776699999999
+ lkvth0we = -2e-12
+ kt1 = 0.010917511
+ kt2 = -0.10990444
+ lk2 = -1.5787889e-9
+ delta = 0.007595625
+ tcjswg = 0.001
+ llc = 0
+ laigc = -2.1190647e-11
+ lln = 1
+ lu0 = 5.409271100000001e-10
+ mjd = 0.26
+ mjs = 0.26
+ lua = 7.8730998e-17
+ lub = -4.3148946000000005e-26
+ luc = 1.578889e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 0
+ rnoia = 0
+ rnoib = 0
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 6e-11
+ pbs = 0.52
+ pu0 = 0.0
+ prt = 0
+ pub = 0
+ puc = 0
+ pud = 0
+ acnqsmod = 0
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 3.744227e-10
+ ngate = 8e+20
+ ub1 = -1.5595112e-18
+ uc1 = -1.6722222e-10
+ tpb = 0.0014
+ ngcon = 1
+ wa0 = 0
+ ute = -1
+ wat = 0.0
+ web = 6843.8
+ wec = -25529.0
+ wlc = 0
+ wln = 1
+ wu0 = 2e-11
+ xgl = -1.09e-8
+ xgw = 0
+ wub = 0
+ wuc = 0
+ wud = 0
+ rbodymod = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ a0 = 5.9444444
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = -94444.467
+ cf = 7.5795e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = -0.014375299
+ k3 = -1.8419
+ em = 1000000.0
+ fprout = 300
+ ll = 0
+ lw = 0
+ u0 = 0.0007882222200000001
+ nfactor = 1
+ w0 = 0
+ ua = -3.1544825e-9
+ ub = 2.30794738e-18
+ uc = 7.77778e-12
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 5.6700000000000005e-9
+ ww = 0
+ xw = 3.4e-9
+ xrcrg1 = 12
+ xrcrg2 = 1
+ wtvoff = 0
+ tvfbsdoff = 0.022
+ nigbacc = 10
+ capmod = 2
+ tvoff = 0.0057943818
+ wku0we = 2e-11
+ keta = 0.088888889
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ mobmod = 0
+ nigbinv = 10
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 4.0264971e-10
+ kt1l = 0
+ ku0we = -0.0007
+ wkvth0we = 2e-12
+ beta0 = 13
+ leta0 = -1.8441422e-9
+ letab = 4.0459126e-8
+ lint = 0
+ trnqsmod = 0
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ lkt1 = -1.4536767e-8
+ lkt2 = 1.3104778e-9
+ lmax = 5.233e-8
+ lmin = 4.333e-8
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ lpe0 = 9.2e-8
+ fnoimod = 1
+ lpeb = 2.5e-7
+ eigbinv = 1.1
+ minv = -0.3
+ lua1 = 1.2526683e-17
+ lub1 = 3.5746048999999995e-26
+ luc1 = 1.5788889e-17
+ ndep = 1e+18
+ dmcgt = 0
+ rgatemod = 0
+ lwlc = 0
+ tcjsw = 0.000357
+ moin = 5.1
+ tnjtsswg = 1
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ nigc = 3.083
+ bigsd = 0.00125
+ noff = 2.7195
+ cigbacc = 0.32875
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ wvoff = 0
+ tnoimod = 0
+ ntox = -0.31099999999999994
+ pcit = 0.0
+ pclm = 2.281309
+ wvsat = 0.0
+ wvth0 = 2.6e-9
+ cigbinv = 0.006
+ phin = 0.15
+ toxref = 3e-9
+ pkt1 = 0
+ lketa = -6.3155556e-9
+ version = 4.5
+ xpart = 1
+ tempmod = 0
+ egidl = 0.29734
+ rbdb = 50
+ prwb = 0
+ pub1 = 0.0
+ prwg = 0
+ )

.model nch_ss_8 nmos (
+ level = 54
+ ngate = 8e+20
+ ngcon = 1
+ wpclm = 0
+ rdsmod = 0
+ wkvth0we = 2e-12
+ wtvfbsdoff = 0
+ igbmod = 1
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ trnqsmod = 0
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ nigbacc = 10
+ ltvfbsdoff = 0
+ pbswgd = 0.95
+ pbswgs = 0.95
+ k2we = 5e-5
+ igcmod = 1
+ dsub = 0.75
+ dtox = 2.7e-10
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ nigbinv = 10
+ rgatemod = 0
+ eta0 = -0.001232
+ etab = -0.88502038
+ tnjtsswg = 1
+ tvfbsdoff = 0.022
+ ptvfbsdoff = 0
+ tvoff = 0.0030235155
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ fnoimod = 1
+ permod = 1
+ eigbinv = 1.1
+ ku0we = -0.0007
+ beta0 = 13
+ leta0 = 1.5454208e-8
+ letab = 3.0054568e-8
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ ppclm = 0
+ voffcv = -0.16942
+ wpemod = 1
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ cigbacc = 0.32875
+ dmcgt = 0
+ tnoimod = 0
+ tcjsw = 0.000357
+ cigbinv = 0.006
+ tpbswg = 0.0009
+ keta = 0.44888889
+ ijthsfwd = 0.01
+ bigsd = 0.00125
+ version = 4.5
+ wvoff = 0
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 2.8614459e-10
+ tempmod = 0
+ kt1l = 0
+ ptvoff = 0
+ wvsat = 0.0
+ wvth0 = 2.6e-9
+ ijthsrev = 0.01
+ lint = 0
+ aigbacc = 0.02
+ lkt1 = -3.9088498e-9
+ lkt2 = 1.6072e-9
+ diomod = 1
+ lmax = 4.333e-8
+ lmin = 3.6e-8
+ lpe0 = 9.2e-8
+ pditsd = 0
+ pditsl = 0
+ lketa = -2.3955556e-8
+ lpeb = 2.5e-7
+ cjswgd = 3.0174000000000004e-10
+ pku0we = -1.5e-18
+ cjswgs = 3.0174000000000004e-10
+ xpart = 1
+ minv = -0.3
+ aigbinv = 0.0163
+ lua1 = 7.1708778e-18
+ lub1 = -2.8298559e-26
+ luc1 = -1.63268e-17
+ egidl = 0.29734
+ ndep = 1e+18
+ lwlc = 0
+ mjswgd = 0.85
+ mjswgs = 0.85
+ moin = 5.1
+ nigc = 3.083
+ tcjswg = 0.001
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ poxedge = 1
+ pkvth0we = -1.3e-19
+ ntox = -0.31099999999999994
+ pcit = 0.0
+ pclm = 2.10165423
+ binunit = 2
+ pvoff = -7e-17
+ fprout = 300
+ phin = 0.15
+ cdscb = 0
+ cdscd = 0
+ vfbsdoff = 0.02
+ pvsat = 0.0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ wk2we = 5e-12
+ pvth0 = 2.3e-16
+ drout = 0.56
+ pkt1 = 0
+ voffl = 0
+ wtvoff = 0
+ paramchk = 1
+ weta0 = 0
+ rbdb = 50
+ prwb = 0
+ pub1 = 0.0
+ prwg = 0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ lpclm = -6.406864000000001e-8
+ rdsw = 100
+ capmod = 2
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ cgidl = 0.22
+ wku0we = 2e-11
+ mobmod = 0
+ ijthdfwd = 0.01
+ a0 = 3.6555556
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 149459.93
+ cf = 7.5795e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.026156861000000003
+ k3 = -1.8419
+ em = 1000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.0039055553
+ pvfbsdoff = 0
+ w0 = 0
+ ua = -2.2580401200000003e-9
+ ub = 1.5627388499999998e-18
+ uc = 2.4e-10
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 5.6700000000000005e-9
+ ww = 0
+ xw = 3.4e-9
+ pbswd = 0.8
+ pbsws = 0.8
+ rshg = 15.6
+ ijthdrev = 0.01
+ pdits = 0
+ njtsswg = 9
+ cigsd = 0.069865
+ laigsd = -2.1777778e-17
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ ckappad = 0.6
+ ckappas = 0.6
+ pk2we = -1e-19
+ tnom = 25
+ pdiblc1 = 0
+ pdiblc2 = 0.0069157
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ pdiblcb = -0.3
+ toxe = 2.47e-9
+ toxm = 2.43e-9
+ tnoia = 0
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ peta0 = 0
+ lkvth0we = -2e-12
+ bigbacc = 0.002588
+ tpbsw = 0.0019
+ wags = 1e-8
+ cjswd = 8.774000000000001e-11
+ cjsws = 8.774000000000001e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ wcit = 0.0
+ kvth0we = 0.00018
+ acnqsmod = 0
+ voff = -0.039834349000000005
+ acde = 0.4
+ lintnoi = -1.5e-8
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ vsat = 101093.02200000003
+ rbodymod = 0
+ vtsswgs = 4.2
+ wint = 0
+ vth0 = 0.343205703
+ toxref = 3e-9
+ wkt1 = 1.2e-9
+ ags = 2.7325299999999997
+ wmax = 0.00090001
+ aigc = 0.011387162
+ wmin = 9.0026e-6
+ cjd = 0.00145199
+ cit = -0.0012536118
+ cjs = 0.00145199
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 3.26497e-9
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ scref = 1e-6
+ wub1 = 0.0
+ pigcd = 2.621
+ aigsd = 0.010773221
+ la0 = -2.0362223e-7
+ bigc = 0.001442
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.0027095388000000003
+ kt1 = -0.20597876
+ kt2 = -0.11596
+ lk2 = -3.5648647e-9
+ wwlc = 0
+ llc = 0
+ lvoff = -7.156111900000001e-9
+ lln = 1
+ lu0 = 3.8817777e-10
+ mjd = 0.26
+ mjs = 0.26
+ lua = 3.4805321000000004e-17
+ lub = -6.633731000000002e-27
+ luc = -9.7999999e-18
+ lud = 0
+ ltvoff = -1.1163261e-10
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 0
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 6e-11
+ pbs = 0.52
+ pk2 = 0
+ lvsat = 0.0013763563899999998
+ cdsc = 0
+ pu0 = 0.0
+ lvth0 = 2.8374218800000004e-9
+ prt = 0
+ cgbo = 0
+ pua = 0
+ pub = 0
+ puc = 0
+ pud = 0
+ cgdl = 3.0874977e-12
+ cgdo = 4.5622265999999996e-11
+ xtid = 3
+ xtis = 3
+ delta = 0.007595625
+ cgsl = 3.0874977e-12
+ cgso = 4.5622265999999996e-11
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 4.8372486e-10
+ ub1 = -2.5247838e-19
+ cigc = 0.000625
+ laigc = -6.2207351e-12
+ uc1 = 4.882e-10
+ tpb = 0.0014
+ wa0 = 0
+ rnoia = 0
+ rnoib = 0
+ nfactor = 1
+ ute = -1
+ wat = 0.0
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 0
+ wlc = 0
+ lku0we = 2.5e-11
+ wln = 1
+ wu0 = 2e-11
+ xgl = -1.09e-8
+ xgw = 0
+ wua = 0
+ wub = 0
+ wuc = 0
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ epsrox = 3.9
+ )

.model nch_ss_9 nmos (
+ level = 54
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ ptvfbsdoff = 0
+ voffl = 0
+ minv = -0.3
+ lub1 = 0
+ weta0 = 0
+ ndep = 1e+18
+ wetab = -1.0073378e-8
+ lwlc = 0
+ moin = 5.1
+ nigc = 3.083
+ cgidl = 0.22
+ lkvth0we = -2e-12
+ njtsswg = 9
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ pvfbsdoff = 0
+ noic = 45200000.0
+ permod = 1
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ acnqsmod = 0
+ pbswd = 0.8
+ pbsws = 0.8
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.018557155
+ pdiblcb = -0.3
+ ntox = -0.31099999999999994
+ pcit = 0
+ pclm = 1.4152454
+ rbodymod = 0
+ phin = 0.15
+ voffcv = -0.16942
+ wpemod = 1
+ pdits = 0
+ cigsd = 0.069865
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ pkt1 = 0
+ bigbacc = 0.002588
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ kvth0we = 0.00018
+ rbdb = 50
+ prwb = 0
+ pub1 = 0
+ prwg = 0
+ wpdiblc2 = -1.7177628e-11
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ lintnoi = -1.5e-8
+ tnoia = 0
+ bigbinv = 0.004953
+ rdsw = 100
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ peta0 = 0
+ tpbswg = 0.0009
+ wketa = 3.3422159e-8
+ tpbsw = 0.0019
+ cjswd = 8.774000000000001e-11
+ cjsws = 8.774000000000001e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ ags = 0.9468331400000001
+ ptvoff = 0
+ cjd = 0.00145199
+ cit = 4.8708935e-5
+ cjs = 0.00145199
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ wkvth0we = 2e-12
+ bvs = 8.7
+ rshg = 15.6
+ waigsd = 3.0716751e-12
+ dlc = 9.8024918e-9
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ trnqsmod = 0
+ diomod = 1
+ la0 = 0
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = 0.0004
+ kt1 = -0.19515831
+ kt2 = -0.052853133
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 3.0174000000000004e-10
+ llc = 0
+ pku0we = -1.5e-18
+ lln = 1
+ cjswgs = 3.0174000000000004e-10
+ lu0 = -6e-12
+ mjd = 0.26
+ mjs = 0.26
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ scref = 1e-6
+ njd = 1.02
+ njs = 1.02
+ pa0 = 0
+ nfactor = 1
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 6e-11
+ pbs = 0.52
+ pigcd = 2.621
+ aigsd = 0.010772879
+ pu0 = 0
+ prt = 0
+ pud = 0
+ tnom = 25
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 1.311952e-9
+ toxe = 2.47e-9
+ ub1 = -8.0649865e-19
+ toxm = 2.43e-9
+ lvoff = 0
+ uc1 = 3.0375074e-11
+ mjswgd = 0.85
+ mjswgs = 0.85
+ tpb = 0.0014
+ rgatemod = 0
+ wa0 = -2.5183444e-7
+ ute = -0.96248296
+ wat = 0
+ tnjtsswg = 1
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -3.7920026e-9
+ lvsat = 0.0003
+ wlc = 0
+ tcjswg = 0.001
+ wln = 1
+ wu0 = -2.4190782e-10
+ xgl = -1.09e-8
+ xgw = 0
+ lvth0 = 0
+ wua = -4.0765791e-17
+ wub = 4.0599742e-26
+ wuc = -7.8572347e-18
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ delta = 0.007595625
+ nigbacc = 10
+ rnoia = 0
+ rnoib = 0
+ wags = -7.4054279e-8
+ wcit = 4.6192733e-10
+ ngate = 8e+20
+ voff = -0.11308442
+ ngcon = 1
+ wpclm = -1.3730014e-7
+ acde = 0.4
+ nigbinv = 10
+ vsat = 103058.98
+ wint = 0
+ gbmin = 1e-12
+ vth0 = 0.37834845
+ fprout = 300
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ wkt1 = -4.4439654e-8
+ wkt2 = -3.5741805e-9
+ wmax = 9.0026e-6
+ xrcrg1 = 12
+ xrcrg2 = 1
+ aigc = 0.011766468
+ wmin = 9.025999999999999e-7
+ wtvoff = -8.3463378e-10
+ wua1 = -7.3834184e-16
+ wub1 = 7.3798399e-25
+ wuc1 = -8.5623711e-19
+ fnoimod = 1
+ bigc = 0.001442
+ wute = -4.0092044e-7
+ eigbinv = 1.1
+ wwlc = 0
+ tvfbsdoff = 0.022
+ capmod = 2
+ cdsc = 0
+ cgbo = 0
+ wku0we = 2e-11
+ cgdl = 3.0874977e-12
+ cgdo = 4.5622265999999996e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.0874977e-12
+ cgso = 4.5622265999999996e-11
+ tvoff = 0.0020036382
+ cigc = 0.000625
+ mobmod = 0
+ xjbvd = 1
+ ijthsfwd = 0.01
+ xjbvs = 1
+ lk2we = -1.5e-12
+ cigbacc = 0.32875
+ ku0we = -0.0007
+ beta0 = 13
+ leta0 = 0
+ tnoimod = 0
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ ijthsrev = 0.01
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ cigbinv = 0.006
+ dlcig = 2.5e-9
+ k2we = 5e-5
+ bgidl = 2320000000.0
+ dsub = 0.75
+ dtox = 2.7e-10
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ a0 = 3.277963
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ version = 4.5
+ at = 72000
+ cf = 7.5795e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.027022307000000002
+ k3 = -1.8419
+ em = 1000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.016099082
+ dmcgt = 0
+ w0 = 0
+ tempmod = 0
+ ua = -1.8192461e-9
+ ub = 2.0991879e-18
+ uc = 7.4172444e-11
+ ud = 0
+ eta0 = 0.3
+ tcjsw = 0.000357
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 5.6700000000000005e-9
+ alpha0 = 2e-10
+ ww = 0
+ alpha1 = 3.6
+ xw = 3.4e-9
+ etab = -0.24888148
+ aigbacc = 0.02
+ bigsd = 0.00125
+ wvoff = 2.3777201e-9
+ pkvth0we = -1.3e-19
+ aigbinv = 0.0163
+ wvsat = -0.0017920539
+ wvth0 = -8.545485e-9
+ toxref = 3e-9
+ waigc = 2.6350949e-11
+ vfbsdoff = 0.02
+ xpart = 1
+ paramchk = 1
+ ltvoff = 0
+ egidl = 0.29734
+ poxedge = 1
+ binunit = 2
+ wtvfbsdoff = 0
+ keta = -0.063711099
+ lku0we = 2.5e-11
+ ijthdfwd = 0.01
+ epsrox = 3.9
+ ltvfbsdoff = 0
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 4e-12
+ rdsmod = 0
+ kt1l = 0
+ igbmod = 1
+ ijthdrev = 0.01
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ pvoff = -7e-17
+ lint = 6.5375218e-9
+ pbswgd = 0.95
+ cdscb = 0
+ cdscd = 0
+ pbswgs = 0.95
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ lkt1 = 0
+ pvsat = 0
+ lmax = 2.001e-5
+ wk2we = 5e-12
+ pvth0 = 2.3e-16
+ lmin = 8.99743e-6
+ drout = 0.56
+ igcmod = 1
+ )

.model nch_ss_10 nmos (
+ level = 54
+ xrcrg1 = 12
+ xrcrg2 = 1
+ cgidl = 0.22
+ vfbsdoff = 0.02
+ wtvoff = -8.9580408e-10
+ nfactor = 1
+ pbswd = 0.8
+ pbsws = 0.8
+ paramchk = 1
+ capmod = 2
+ wku0we = 2e-11
+ mobmod = 0
+ pdits = 0
+ cigsd = 0.069865
+ nigbacc = 10
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ ijthdfwd = 0.01
+ keta = -0.064075044
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ nigbinv = 10
+ lags = -6.3328546e-8
+ wtvfbsdoff = 0
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 1.1377416e-9
+ tnoia = 0
+ laigsd = 1.1048614e-17
+ ijthdrev = 0.01
+ kt1l = 0
+ peta0 = 0
+ ltvfbsdoff = 0
+ lpdiblc2 = -6.1589259e-10
+ wketa = 3.7630763e-8
+ lint = 6.5375218e-9
+ tpbsw = 0.0019
+ lkt1 = -4.5537316e-8
+ lkt2 = -1.2972142e-8
+ cjswd = 8.774000000000001e-11
+ lmax = 8.99743e-6
+ cjsws = 8.774000000000001e-11
+ lmin = 8.974099999999999e-7
+ fnoimod = 1
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ lpe0 = 9.2e-8
+ eigbinv = 1.1
+ lpeb = 2.5e-7
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ minv = -0.3
+ lua1 = -4.3996966e-16
+ lub1 = 2.6060002e-25
+ luc1 = 3.9191378e-17
+ ndep = 1e+18
+ lute = -3.7058959e-8
+ lwlc = 0
+ ptvfbsdoff = 0
+ moin = 5.1
+ lkvth0we = -2e-12
+ nigc = 3.083
+ scref = 1e-6
+ pigcd = 2.621
+ aigsd = 0.010772879
+ cigbacc = 0.32875
+ acnqsmod = 0
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ lvoff = -1.4242682e-8
+ toxref = 3e-9
+ tnoimod = 0
+ pags = 2.8299487e-13
+ rbodymod = 0
+ lvsat = 0.0003
+ lvth0 = 5.1255324e-8
+ ntox = -0.31099999999999994
+ pcit = -1.846418e-16
+ pclm = 1.4152454
+ cigbinv = 0.006
+ delta = 0.007595625
+ laigc = -1.4938914e-10
+ tvfbsdoff = 0.022
+ rnoia = 0
+ rnoib = 0
+ phin = 0.15
+ pkt1 = 4.9872912e-14
+ pkt2 = 1.3351872e-15
+ pketa = -3.7835355e-14
+ version = 4.5
+ ngate = 8e+20
+ ltvoff = -2.0733557e-10
+ ngcon = 1
+ tempmod = 0
+ wpclm = -1.3730014e-7
+ wpdiblc2 = -4.8108443e-11
+ gbmin = 1e-12
+ rbdb = 50
+ pua1 = 6.0905252e-22
+ prwb = 0
+ prwg = 0
+ pub1 = -5.9738158e-31
+ jswgd = 1.28e-13
+ puc1 = 1.7562426e-23
+ jswgs = 1.28e-13
+ rbpb = 50
+ rbpd = 50
+ aigbacc = 0.02
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ pute = 3.9602525e-13
+ lku0we = 2.5e-11
+ rdsw = 100
+ wvfbsdoff = 0
+ epsrox = 3.9
+ lvfbsdoff = 0
+ rdsmod = 0
+ aigbinv = 0.0163
+ igbmod = 1
+ wkvth0we = 2e-12
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ pbswgd = 0.95
+ pbswgs = 0.95
+ rshg = 15.6
+ trnqsmod = 0
+ tvoff = 0.0020267011
+ igcmod = 1
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ poxedge = 1
+ ku0we = -0.0007
+ beta0 = 13
+ tnom = 25
+ rgatemod = 0
+ leta0 = 0
+ binunit = 2
+ tnjtsswg = 1
+ toxe = 2.47e-9
+ paigsd = -9.9503825e-23
+ toxm = 2.43e-9
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ permod = 1
+ wags = -1.0553313e-7
+ wcit = 4.8246591e-10
+ dmcgt = 0
+ tcjsw = 0.000357
+ voff = -0.11150014
+ acde = 0.4
+ voffcv = -0.16942
+ wpemod = 1
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ vsat = 103058.98
+ wint = 0
+ vth0 = 0.37264708
+ wkt1 = -4.9987253e-8
+ wkt2 = -3.7226997e-9
+ wmax = 9.0026e-6
+ aigc = 0.011783086
+ bigsd = 0.00125
+ wmin = 9.025999999999999e-7
+ wvoff = 2.6904676e-9
+ wua1 = -8.0608962e-16
+ wub1 = 8.0443355e-25
+ wuc1 = -2.8097884e-18
+ wvsat = -0.0017920539
+ wvth0 = -8.928173e-9
+ bigc = 0.001442
+ wute = -4.4497219e-7
+ wwlc = 0
+ waigc = 2.7413515e-11
+ tpbswg = 0.0009
+ njtsswg = 9
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.0874977e-12
+ cgdo = 4.5622265999999996e-11
+ xtid = 3
+ xtis = 3
+ lketa = 3.2718606e-9
+ xtsswgd = 0.18
+ cgsl = 3.0874977e-12
+ ijthsfwd = 0.01
+ cgso = 4.5622265999999996e-11
+ xtsswgs = 0.18
+ cigc = 0.000625
+ xpart = 1
+ ckappad = 0.6
+ ckappas = 0.6
+ ptvoff = 5.4992103e-16
+ pdiblc1 = 0
+ pdiblc2 = 0.018625664
+ pdiblcb = -0.3
+ waigsd = 3.0716862e-12
+ egidl = 0.29734
+ diomod = 1
+ ijthsrev = 0.01
+ pditsd = 0
+ pditsl = 0
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ cjswgd = 3.0174000000000004e-10
+ pku0we = -1.5e-18
+ cjswgs = 3.0174000000000004e-10
+ ags = 0.9538774700000001
+ bigbacc = 0.002588
+ cjd = 0.00145199
+ cit = -7.7402473e-5
+ cjs = 0.00145199
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 9.8024918e-9
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ k2we = 5e-5
+ kvth0we = 0.00018
+ dsub = 0.75
+ dtox = 2.7e-10
+ mjswgd = 0.85
+ mjswgs = 0.85
+ pvfbsdoff = 0
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ la0 = -2.0592205e-6
+ lintnoi = -1.5e-8
+ ppdiblc2 = 2.7806803e-16
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = 0.094882725
+ tcjswg = 0.001
+ kt1 = -0.19009298
+ lk2 = -1.3154073e-8
+ kt2 = -0.051410181
+ bigbinv = 0.004953
+ llc = 0
+ vtsswgd = 4.2
+ lln = 1
+ vtsswgs = 4.2
+ lu0 = -2.0024409000000003e-9
+ mjd = 0.26
+ lua = -2.2049077e-16
+ mjs = 0.26
+ lub = -1.5408759e-27
+ luc = 1.1211784e-18
+ lud = 0
+ pvoff = -2.8816001e-15
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 3.0846188e-13
+ eta0 = 0.3
+ nsd = 1e+20
+ pbd = 0.52
+ pat = -8.2187187e-9
+ pbs = 0.52
+ pk2 = -1.9754424e-15
+ cdscb = 0
+ cdscd = 0
+ etab = -0.24888148
+ pu0 = 9.9503831e-18
+ pvsat = 0
+ prt = 0
+ pua = 2.7693259e-23
+ pub = -6.3482817e-32
+ puc = -1.7214163e-23
+ pud = 0
+ wk2we = 5e-12
+ pvth0 = 3.6703639e-15
+ drout = 0.56
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 1.3608919e-9
+ ub1 = -8.3548641e-19
+ uc1 = 2.6015633e-11
+ paigc = -9.5524673e-18
+ tpb = 0.0014
+ wa0 = -2.8614611e-7
+ ute = -0.95836072
+ wat = 0.00092088084
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -3.5722648e-9
+ voffl = 0
+ wlc = 0
+ wln = 1
+ wu0 = -2.4301465e-10
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -4.3846243e-17
+ wub = 4.7661234e-26
+ wuc = -5.9424224e-18
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ a0 = 3.5070197
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ weta0 = 0
+ pkvth0we = -1.3e-19
+ at = 61490.242
+ cf = 7.5795e-11
+ wetab = -1.0073378e-8
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.028485497
+ k3 = -1.8419
+ em = 1000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.016321155
+ fprout = 300
+ w0 = 0
+ ua = -1.7947198e-9
+ ub = 2.0993593e-18
+ uc = 7.4047731e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 5.6700000000000005e-9
+ ww = 0
+ xw = 3.4e-9
+ )

.model nch_ss_11 nmos (
+ level = 54
+ ku0we = -0.0007
+ beta0 = 13
+ wku0we = 2e-11
+ leta0 = 0
+ rbdb = 50
+ mobmod = 0
+ pua1 = 9.7840116e-23
+ prwb = 0
+ prwg = 0
+ pub1 = -1.2240721e-31
+ puc1 = -3.5940917e-24
+ a0 = 1.2386098
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ wtvfbsdoff = 0
+ at = 220073.87
+ cf = 7.5795e-11
+ rbpb = 50
+ rbpd = 50
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.027732723
+ k3 = -1.8419
+ rbps = 50
+ em = 1000000.0
+ rbsb = 50
+ pvag = 1.2
+ ll = 0
+ lw = 0
+ u0 = 0.015821688
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ w0 = 0
+ ua = -1.9419497e-9
+ ub = 2.1613601e-18
+ uc = 9.7509556e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 5.6700000000000005e-9
+ ww = 0
+ xw = 3.4e-9
+ rdsw = 100
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ ijthsfwd = 0.01
+ ltvfbsdoff = 0
+ dmcgt = 0
+ tcjsw = 0.000357
+ laigsd = -9.7335958e-18
+ ijthsrev = 0.01
+ rshg = 15.6
+ njtsswg = 9
+ bigsd = 0.00125
+ ptvfbsdoff = 0
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ wvoff = -7.7864574e-9
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.014827337
+ pdiblcb = -0.3
+ wvsat = -0.0017920539
+ ppdiblc2 = 2.4623293e-15
+ tnom = 25
+ wvth0 = 1.3738106e-9
+ toxe = 2.47e-9
+ toxm = 2.43e-9
+ waigc = -9.5733062e-12
+ lketa = -3.0044615e-8
+ bigbacc = 0.002588
+ xpart = 1
+ wags = 1.2560313e-6
+ kvth0we = 0.00018
+ toxref = 3e-9
+ egidl = 0.29734
+ pkvth0we = -1.3e-19
+ wcit = 1.5976377e-10
+ ags = 0.30741392
+ cjd = 0.00145199
+ cit = 0.0013334381
+ voff = -0.11121991
+ lintnoi = -1.5e-8
+ cjs = 0.00145199
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ acde = 0.4
+ dlc = 9.8024918e-9
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ k3b = 1.9326
+ vtsswgs = 4.2
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ vsat = 103058.98
+ wint = 0
+ vfbsdoff = 0.02
+ vth0 = 0.42119507
+ wkt1 = 1.9028643e-8
+ wkt2 = -3.7425887e-9
+ wmax = 9.0026e-6
+ la0 = -4.0335612e-8
+ aigc = 0.011680759
+ wmin = 9.025999999999999e-7
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.046256700000000005
+ kt1 = -0.22273968
+ lk2 = -1.2484105e-8
+ kt2 = -0.052902736
+ llc = 0
+ lln = 1
+ lu0 = -1.5579156e-9
+ mjd = 0.26
+ ltvoff = -6.7137092e-10
+ lua = -8.9456155e-17
+ mjs = 0.26
+ lub = -5.6721601e-26
+ luc = -1.9759846e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = -3.420874e-13
+ nsd = 1e+20
+ pbd = 0.52
+ pat = -3.5866881e-9
+ pbs = 0.52
+ pk2 = 6.3553328e-16
+ pvfbsdoff = 0
+ paramchk = 1
+ pu0 = 2.6298232e-17
+ wua1 = -2.3169366e-16
+ wub1 = 2.7075449e-25
+ prt = 0
+ wuc1 = 2.096158e-17
+ pua = -3.3732216e-24
+ pub = 1.7089792e-32
+ puc = 7.8894695e-24
+ pud = 0
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 9.9427719e-10
+ bigc = 0.001442
+ ub1 = -5.7879508e-19
+ uc1 = 6.536871e-11
+ pvoff = 6.4428631e-15
+ tpb = 0.0014
+ wwlc = 0
+ wa0 = 4.4480813e-7
+ ute = -1
+ wat = -0.0042836479
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -6.5059453e-9
+ cdscb = 0
+ cdscd = 0
+ lku0we = 2.5e-11
+ wlc = 0
+ wln = 1
+ wu0 = -2.6138302e-10
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -8.9400845e-18
+ wub = -4.2869787e-26
+ pvsat = 0
+ wuc = -3.4148751e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ epsrox = 3.9
+ cdsc = 0
+ wk2we = 5e-12
+ pvth0 = -5.4984018e-15
+ drout = 0.56
+ cgbo = 0
+ cgdl = 3.0874977e-12
+ cgdo = 4.5622265999999996e-11
+ xtid = 3
+ xtis = 3
+ ijthdfwd = 0.01
+ cgsl = 3.0874977e-12
+ paigc = 2.3365803e-17
+ cgso = 4.5622265999999996e-11
+ cigc = 0.000625
+ rdsmod = 0
+ nfactor = 1
+ voffl = 0
+ igbmod = 1
+ weta0 = 0
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ wetab = -1.0073378e-8
+ pbswgd = 0.95
+ pbswgs = 0.95
+ ijthdrev = 0.01
+ igcmod = 1
+ cgidl = 0.22
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ lpdiblc2 = 2.7646188e-9
+ nigbacc = 10
+ k2we = 5e-5
+ pbswd = 0.8
+ pbsws = 0.8
+ dsub = 0.75
+ dtox = 2.7e-10
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ nigbinv = 10
+ paigsd = 8.7660773e-23
+ eta0 = 0.3
+ pdits = 0
+ etab = -0.24888148
+ cigsd = 0.069865
+ lkvth0we = -2e-12
+ permod = 1
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ pk2we = -1e-19
+ fnoimod = 1
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ acnqsmod = 0
+ eigbinv = 1.1
+ voffcv = -0.16942
+ wpemod = 1
+ tnoia = 0
+ rbodymod = 0
+ peta0 = 0
+ wketa = -4.0591301e-8
+ tpbsw = 0.0019
+ cjswd = 8.774000000000001e-11
+ cjsws = 8.774000000000001e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ cigbacc = 0.32875
+ wpdiblc2 = -2.5023346e-9
+ tnoimod = 0
+ tpbswg = 0.0009
+ cigbinv = 0.006
+ scref = 1e-6
+ ptvoff = 2.4706364e-16
+ pigcd = 2.621
+ keta = -0.026640801
+ aigsd = 0.010772879
+ waigsd = 3.0714759e-12
+ version = 4.5
+ lvoff = -1.4492081e-8
+ lags = 5.1202402e-7
+ wkvth0we = 2e-12
+ tempmod = 0
+ jswd = 1.28e-13
+ diomod = 1
+ jsws = 1.28e-13
+ lcit = -1.1790652999999998e-10
+ lvsat = 0.0003
+ kt1l = 0
+ lvth0 = 8.0476154e-9
+ pditsd = 0
+ pditsl = 0
+ trnqsmod = 0
+ cjswgd = 3.0174000000000004e-10
+ tvfbsdoff = 0.022
+ pku0we = -1.5e-18
+ cjswgs = 3.0174000000000004e-10
+ delta = 0.007595625
+ laigc = -5.8318716e-11
+ aigbacc = 0.02
+ lint = 6.5375218e-9
+ rnoia = 0
+ rnoib = 0
+ lkt1 = -1.6481753e-8
+ lkt2 = -1.1643768e-8
+ lmax = 8.974099999999999e-7
+ lmin = 4.4741e-7
+ pketa = 3.1782283e-14
+ mjswgd = 0.85
+ lpe0 = 9.2e-8
+ ngate = 8e+20
+ mjswgs = 0.85
+ lpeb = 2.5e-7
+ ngcon = 1
+ wpclm = -1.3730014e-7
+ aigbinv = 0.0163
+ tcjswg = 0.001
+ minv = -0.3
+ rgatemod = 0
+ lua1 = -1.1368255e-16
+ lub1 = 3.2144732e-26
+ luc1 = 4.1671397e-18
+ gbmin = 1e-12
+ tnjtsswg = 1
+ ndep = 1e+18
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ lwlc = 0
+ moin = 5.1
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ nigc = 3.083
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ poxedge = 1
+ fprout = 300
+ xrcrg1 = 12
+ xrcrg2 = 1
+ pags = -9.2879744e-13
+ ntox = -0.31099999999999994
+ pcit = 1.025631e-16
+ binunit = 2
+ pclm = 1.4152454
+ tvoff = 0.0025480892
+ wtvoff = -5.5551488e-10
+ xjbvd = 1
+ phin = 0.15
+ xjbvs = 1
+ lk2we = -1.5e-12
+ pkt1 = -1.1551235e-14
+ pkt2 = 1.3528884e-15
+ capmod = 2
+ )

.model nch_ss_12 nmos (
+ level = 54
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ ptvfbsdoff = 0
+ cigbacc = 0.32875
+ laigsd = -9.015225e-17
+ wkvth0we = 2e-12
+ tnoia = 0
+ tnoimod = 0
+ trnqsmod = 0
+ peta0 = 0
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ wketa = 1.7936379e-8
+ tpbsw = 0.0019
+ a0 = 1.7327189
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ cigbinv = 0.006
+ at = 153009.14
+ cf = 7.5795e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.021241707
+ k3 = -1.8419
+ em = 1000000.0
+ cjswd = 8.774000000000001e-11
+ ll = -1.18e-13
+ cjsws = 8.774000000000001e-11
+ lw = 0
+ u0 = 0.013715620999999999
+ w0 = 0
+ mjswd = 0.11
+ ua = -2.1226101e-9
+ ub = 2.1428106e-18
+ uc = 6.8443458e-11
+ ud = 0
+ mjsws = 0.11
+ agidl = 9.41e-8
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 5.6700000000000005e-9
+ ww = 0
+ xw = 3.4e-9
+ k2we = 5e-5
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ dsub = 0.75
+ dtox = 2.7e-10
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ version = 4.5
+ rgatemod = 0
+ tnjtsswg = 1
+ tempmod = 0
+ eta0 = 0.3
+ etab = -0.24888148
+ aigbacc = 0.02
+ scref = 1e-6
+ pigcd = 2.621
+ aigsd = 0.010772879
+ toxref = 3e-9
+ lvoff = -6.0911145e-9
+ aigbinv = 0.0163
+ lvsat = 0.0003
+ lvth0 = -4.941492e-9
+ tvfbsdoff = 0.022
+ delta = 0.007595625
+ laigc = -1.9233809e-11
+ rnoia = 0
+ rnoib = 0
+ ltvoff = -1.0250882e-10
+ pketa = 6.0301037e-15
+ ngate = 8e+20
+ ngcon = 1
+ wpclm = -2.8227848e-7
+ poxedge = 1
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ lku0we = 2.5e-11
+ wvfbsdoff = 0
+ epsrox = 3.9
+ lvfbsdoff = 0
+ binunit = 2
+ rdsmod = 0
+ ijthsfwd = 0.01
+ igbmod = 1
+ keta = -0.041938217
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ lags = 4.5664516e-7
+ pbswgd = 0.95
+ pbswgs = 0.95
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 1.7314929e-10
+ ijthsrev = 0.01
+ igcmod = 1
+ kt1l = 0
+ tvoff = 0.0012552207
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ lint = 9.7879675e-9
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ lkt1 = -9.5958544e-9
+ lkt2 = -3.7159363e-9
+ lmax = 4.4741e-7
+ lmin = 2.1410000000000002e-7
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ ku0we = -0.0007
+ paigsd = 8.167794e-23
+ ppdiblc2 = -2.773275e-15
+ beta0 = 13
+ minv = -0.3
+ lua1 = -3.2594611e-17
+ lub1 = -2.740043e-26
+ leta0 = 0
+ luc1 = -3.5163101e-18
+ ndep = 1e+18
+ ppclm = 6.379047e-14
+ lwlc = 0
+ permod = 1
+ moin = 5.1
+ dlcig = 2.5e-9
+ nigc = 3.083
+ bgidl = 2320000000.0
+ njtsswg = 9
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ pkvth0we = -1.3e-19
+ dmcgt = 0
+ voffcv = -0.16942
+ ckappad = 0.6
+ wpemod = 1
+ ckappas = 0.6
+ tcjsw = 0.000357
+ pdiblc1 = 0
+ pdiblc2 = 0.026288388
+ pags = 8.4375107e-13
+ pdiblcb = -0.3
+ ntox = -0.31099999999999994
+ pcit = -6.2892012e-17
+ pclm = 1.5752657
+ vfbsdoff = 0.02
+ phin = 0.15
+ bigsd = 0.00125
+ pkt1 = -4.7748923e-16
+ pkt2 = -1.2933793e-15
+ bigbacc = 0.002588
+ wvoff = 1.1733398e-8
+ paramchk = 1
+ wvsat = -0.0017920539
+ kvth0we = 0.00018
+ wvth0 = -1.6774896e-8
+ tpbswg = 0.0009
+ rbdb = 50
+ pua1 = 1.9082335e-23
+ prwb = 0
+ prwg = 0
+ pub1 = -2.3158905e-32
+ puc1 = -7.9472634e-24
+ waigc = 5.7897385e-11
+ lintnoi = -1.5e-8
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ rdsw = 100
+ ags = 0.43327497
+ lketa = -2.3313752e-8
+ ijthdfwd = 0.01
+ ptvoff = -1.6297696e-16
+ xpart = 1
+ cjd = 0.00145199
+ cit = 0.00067194759
+ cjs = 0.00145199
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ waigsd = 3.0714895e-12
+ dlc = 1.30529375e-8
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ egidl = 0.29734
+ diomod = 1
+ la0 = -2.5774361e-7
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.016748218999999998
+ pditsd = 0
+ pditsl = 0
+ kt1 = -0.23838945
+ ijthdrev = 0.01
+ lk2 = -9.6280577e-9
+ kt2 = -0.070920535
+ cjswgd = 3.0174000000000004e-10
+ pku0we = -1.5e-18
+ cjswgs = 3.0174000000000004e-10
+ llc = -1.18e-13
+ lln = 0.7
+ rshg = 15.6
+ lu0 = -6.3124579e-10
+ mjd = 0.26
+ lua = -9.9655811e-18
+ mjs = 0.26
+ lub = -4.8559819e-26
+ luc = -6.9707629e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 9.4027643e-14
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 2.6083516999999997e-9
+ lpdiblc2 = -2.2782436e-9
+ pbs = 0.52
+ pk2 = 9.5548939e-17
+ pu0 = 8.1677938e-18
+ prt = 0
+ pua = -7.1355685e-24
+ pub = 6.4921301e-33
+ puc = 2.8995668e-24
+ pud = 0
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 8.0998641e-10
+ ub1 = -4.4346517e-19
+ uc1 = 8.2831095e-11
+ mjswgd = 0.85
+ mjswgs = 0.85
+ tpb = 0.0014
+ wa0 = -5.4636242e-7
+ nfactor = 1
+ pvfbsdoff = 0
+ ute = -1
+ wat = -0.018363284
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -5.2787082e-9
+ tcjswg = 0.001
+ wlc = 0
+ wln = 1
+ wu0 = -2.2017747999999998e-10
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -3.8929611e-19
+ wub = -1.8784192e-26
+ wuc = -2.2808063e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ tnom = 25
+ pvoff = -2.1458734e-15
+ toxe = 2.47e-9
+ toxm = 2.43e-9
+ cdscb = 0
+ cdscd = 0
+ lkvth0we = -2e-12
+ pvsat = 0
+ wk2we = 5e-12
+ pvth0 = 2.4870293e-15
+ drout = 0.56
+ paigc = -6.3213007e-18
+ nigbacc = 10
+ voffl = 0
+ acnqsmod = 0
+ wags = -2.7724881e-6
+ fprout = 300
+ weta0 = 0
+ wetab = -1.0073378e-8
+ wcit = 5.3579813e-10
+ xrcrg1 = 12
+ xrcrg2 = 1
+ lpclm = -7.0408907e-8
+ voff = -0.13031302
+ rbodymod = 0
+ nigbinv = 10
+ acde = 0.4
+ cgidl = 0.22
+ vsat = 103058.98
+ wtvoff = 3.7639557e-10
+ wint = 0
+ vth0 = 0.45071577
+ wkt1 = -6.1389616e-9
+ wkt2 = 2.2716562e-9
+ wmax = 9.0026e-6
+ wtvfbsdoff = 0
+ aigc = 0.01159193
+ wmin = 9.025999999999999e-7
+ capmod = 2
+ pbswd = 0.8
+ pbsws = 0.8
+ ltvfbsdoff = 0
+ fnoimod = 1
+ wua1 = -5.2698704e-17
+ wub1 = 4.5190152e-26
+ wku0we = 2e-11
+ wuc1 = 3.0855152e-17
+ eigbinv = 1.1
+ wpdiblc2 = 9.3967661e-9
+ bigc = 0.001442
+ mobmod = 0
+ wwlc = 0
+ pdits = 0
+ cigsd = 0.069865
+ cdsc = 0
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ cgbo = 0
+ cgdl = 3.0874977e-12
+ cgdo = 4.5622265999999996e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.0874977e-12
+ cgso = 4.5622265999999996e-11
+ cigc = 0.000625
+ )

.model nch_ss_13 nmos (
+ level = 54
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ lint = 9.7879675e-9
+ bigsd = 0.00125
+ lkt1 = -3.621126e-9
+ lkt2 = -5.6046527e-10
+ lmax = 2.1410000000000002e-7
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ lmin = 8.833e-8
+ wvoff = -2.233608000000001e-9
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ wvsat = -0.00035982647999999954
+ minv = -0.3
+ wvth0 = -3.2626169999999995e-9
+ lua1 = 8.0644671e-18
+ lub1 = -5.2760301e-26
+ luc1 = -4.6427809e-18
+ ags = 2.5974682
+ ndep = 1e+18
+ waigc = 3.6164887e-11
+ cjd = 0.00145199
+ cit = 0.0010410649
+ cjs = 0.00145199
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ lwlc = 0
+ dlc = 1.30529375e-8
+ k3b = 1.9326
+ moin = 5.1
+ lkvth0we = -2e-12
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ nigc = 3.083
+ lketa = -1.0074554e-8
+ xpart = 1
+ la0 = -3.95931149e-8
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.0014760989
+ toxref = 3e-9
+ kt1 = -0.26670569
+ lk2 = -2.2996724e-9
+ kt2 = -0.085875374
+ llc = -1.18e-13
+ lln = 0.7
+ a0 = 0.69883298
+ a1 = 0
+ a2 = 1
+ lu0 = -2.0539706e-10
+ b0 = 0
+ b1 = 0
+ acnqsmod = 0
+ mjd = 0.26
+ lua = 2.3685126e-17
+ mjs = 0.26
+ lub = -3.581049857e-26
+ luc = -1.971816e-18
+ lud = 0
+ at = 80629.42
+ cf = 7.5795e-11
+ lwc = 0
+ noff = 2.7195
+ lwl = 0
+ lwn = 1
+ ef = 1.0
+ k1 = 0.274
+ k2 = -0.013489977
+ k3 = -1.8419
+ em = 1000000.0
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ njd = 1.02
+ njs = 1.02
+ nfactor = 1
+ pa0 = 5.1229998e-14
+ egidl = 0.29734
+ ll = -1.18e-13
+ lw = 0
+ u0 = 0.011697379999999999
+ w0 = 0
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 8.8157566e-10
+ pbs = 0.52
+ ua = -2.2820921e-9
+ ub = 2.0823870489000003e-18
+ uc = 4.4751766e-11
+ ud = 0
+ pk2 = 1.6389978e-16
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 5.6700000000000005e-9
+ ww = 0
+ xw = 3.4e-9
+ pu0 = -2.2541017e-17
+ prt = 0
+ pua = 6.5907354e-24
+ pub = -1.1536808500000001e-32
+ puc = -4.2264406e-24
+ pud = 0
+ pags = -3.4153056e-19
+ rbodymod = 0
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 6.1728936e-10
+ ub1 = -3.2327621e-19
+ uc1 = 8.8169819e-11
+ ntox = -0.31099999999999994
+ pcit = -6.0109378e-17
+ pclm = 1.3619854
+ tpb = 0.0014
+ wa0 = -3.4353242e-7
+ ute = -1
+ wat = -0.010179511
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -5.6026458e-9
+ wlc = 0
+ wln = 1
+ wu0 = -7.4638093e-11
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -6.5442869e-17
+ wub = 6.6660889e-26
+ wuc = 1.0964484e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ ltvoff = 4.8985213e-12
+ phin = 0.15
+ pvfbsdoff = 0
+ nigbacc = 10
+ pkt1 = 2.8243122e-15
+ pkt2 = -3.7226831e-16
+ wpdiblc2 = -7.3538749e-9
+ lku0we = 2.5e-11
+ pvoff = 8.011494700000001e-16
+ rbdb = 50
+ pua1 = -3.4072796e-24
+ prwb = 0
+ prwg = 0
+ pub1 = 3.7649133e-33
+ epsrox = 3.9
+ puc1 = 3.7978198e-24
+ cdscb = 0
+ cdscd = 0
+ rbpb = 50
+ rbpd = 50
+ nigbinv = 10
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ pvsat = -3.0219949000000006e-10
+ wk2we = 5e-12
+ pvth0 = -3.6404360000000004e-16
+ rdsw = 100
+ drout = 0.56
+ rdsmod = 0
+ igbmod = 1
+ paigc = -1.7357437e-18
+ voffl = 0
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ pbswgd = 0.95
+ pbswgs = 0.95
+ weta0 = 0
+ wetab = -1.0073378e-8
+ wkvth0we = 2e-12
+ fnoimod = 1
+ lpclm = -2.540677e-8
+ igcmod = 1
+ eigbinv = 1.1
+ rshg = 15.6
+ trnqsmod = 0
+ cgidl = 0.22
+ pbswd = 0.8
+ pbsws = 0.8
+ paigsd = -5.1229584e-23
+ rgatemod = 0
+ tnom = 25
+ cigbacc = 0.32875
+ tnjtsswg = 1
+ toxe = 2.47e-9
+ toxm = 2.43e-9
+ permod = 1
+ pdits = 0
+ cigsd = 0.069865
+ tnoimod = 0
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ cigbinv = 0.006
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ wags = 1.2263337999999998e-6
+ voffcv = -0.16942
+ wpemod = 1
+ wcit = 5.2261028e-10
+ tnoia = 0
+ voff = -0.1572150866
+ version = 4.5
+ acde = 0.4
+ tempmod = 0
+ peta0 = 0
+ vsat = 102561.23895
+ wint = 0
+ vth0 = 0.46521233990000005
+ wketa = 1.0437078e-7
+ wkt1 = -2.1787309999999998e-8
+ wkt2 = -2.0937989e-9
+ tpbsw = 0.0019
+ wmax = 9.0026e-6
+ aigc = 0.011522737
+ wmin = 9.025999999999999e-7
+ cjswd = 8.774000000000001e-11
+ aigbacc = 0.02
+ cjsws = 8.774000000000001e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ wua1 = 5.3887147e-17
+ wub1 = -8.2410881e-26
+ wuc1 = -2.4808749e-17
+ tpbswg = 0.0009
+ bigc = 0.001442
+ wwlc = 0
+ aigbinv = 0.0163
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.0874977e-12
+ cgdo = 4.5622265999999996e-11
+ xtid = 3
+ xtis = 3
+ ptvoff = 8.9623963e-17
+ ijthsfwd = 0.01
+ scref = 1e-6
+ cgsl = 3.0874977e-12
+ cgso = 4.5622265999999996e-11
+ cigc = 0.000625
+ waigsd = 3.0721194e-12
+ pigcd = 2.621
+ aigsd = 0.010772879
+ diomod = 1
+ lvoff = -4.1479246e-10
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 3.0174000000000004e-10
+ pku0we = -1.5e-18
+ cjswgs = 3.0174000000000004e-10
+ lvsat = 0.00040503965999999996
+ tvfbsdoff = 0.022
+ ijthsrev = 0.01
+ lvth0 = -8.000254980000001e-9
+ poxedge = 1
+ delta = 0.007595625
+ laigc = -4.6341008e-12
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ binunit = 2
+ rnoia = 0
+ rnoib = 0
+ mjswgd = 0.85
+ mjswgs = 0.85
+ k2we = 5e-5
+ pketa = -1.2207451e-14
+ tcjswg = 0.001
+ ngate = 8e+20
+ dsub = 0.75
+ ngcon = 1
+ dtox = 2.7e-10
+ wpclm = -2.3899735e-8
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ ppdiblc2 = 7.6111026e-16
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ eta0 = 0.3
+ etab = -0.24888148
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ fprout = 300
+ wtvfbsdoff = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ pkvth0we = -1.3e-19
+ ltvfbsdoff = 0
+ wtvoff = -8.2076521e-10
+ tvoff = 0.00074618122
+ vfbsdoff = 0.02
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ capmod = 2
+ njtsswg = 9
+ wku0we = 2e-11
+ paramchk = 1
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ ku0we = -0.0007
+ mobmod = 0
+ beta0 = 13
+ leta0 = 0
+ ckappad = 0.6
+ ptvfbsdoff = 0
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.022446923
+ pdiblcb = -0.3
+ ppclm = 9.2725546e-15
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ ijthdfwd = 0.01
+ keta = -0.10468292
+ bigbacc = 0.002588
+ laigsd = 3.9592657e-17
+ lags = 3.7696529e-13
+ dmcgt = 0
+ tcjsw = 0.000357
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 9.5265533e-11
+ kvth0we = 0.00018
+ ijthdrev = 0.01
+ kt1l = 0
+ lintnoi = -1.5e-8
+ lpdiblc2 = -1.4676946e-9
+ bigbinv = 0.004953
+ )

.model nch_ss_14 nmos (
+ level = 54
+ poxedge = 1
+ binunit = 2
+ scref = 1e-6
+ toxref = 3e-9
+ pigcd = 2.621
+ aigsd = 0.010772879
+ wags = 1.2263301999999999e-6
+ lvoff = -2.0518068800000008e-9
+ pkvth0we = -1.3e-19
+ wcit = -1.7332863999999998e-10
+ tvfbsdoff = 0.022
+ voff = -0.13980004150000003
+ lvsat = 0.0024133598900000003
+ lvth0 = 2.23756691e-9
+ acde = 0.4
+ delta = 0.007595625
+ vsat = 81196.12610000001
+ laigc = -2.2637509e-11
+ wint = 0
+ vfbsdoff = 0.02
+ vth0 = 0.3562993353
+ ltvoff = 1.2509019e-10
+ wkt1 = 8.5030806e-8
+ wkt2 = 1.6147625e-8
+ rnoia = 0
+ rnoib = 0
+ wmax = 9.0026e-6
+ aigc = 0.011714263
+ wmin = 9.025999999999999e-7
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ pketa = 8.4378567e-15
+ ngate = 8e+20
+ paramchk = 1
+ ngcon = 1
+ wpclm = 3.4675908e-7
+ wua1 = -1.154179e-16
+ wub1 = 3.1505286e-27
+ wuc1 = 9.7519251e-17
+ lku0we = 2.5e-11
+ a0 = -0.035582299999999956
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ bigc = 0.001442
+ gbmin = 1e-12
+ epsrox = 3.9
+ at = 65883.509
+ cf = 7.5795e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = -0.032587969
+ k3 = -1.8419
+ wvfbsdoff = 0
+ em = 1000000.0
+ wwlc = 0
+ jswgd = 1.28e-13
+ lvfbsdoff = 0
+ jswgs = 1.28e-13
+ ll = 0
+ lw = 0
+ u0 = 0.008294596199999999
+ w0 = 0
+ ua = -2.421907e-9
+ ub = 1.9130826320999997e-18
+ uc = 4.338735e-12
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 5.6700000000000005e-9
+ ww = 0
+ xw = 3.4e-9
+ rdsmod = 0
+ cdsc = 0
+ igbmod = 1
+ cgbo = 0
+ cgdl = 3.0874977e-12
+ cgdo = 4.5622265999999996e-11
+ xtid = 3
+ xtis = 3
+ ijthdfwd = 0.01
+ cgsl = 3.0874977e-12
+ cgso = 4.5622265999999996e-11
+ cigc = 0.000625
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ pbswgd = 0.95
+ pbswgs = 0.95
+ njtsswg = 9
+ igcmod = 1
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ ijthdrev = 0.01
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.006833075
+ pdiblcb = -0.3
+ tvoff = -0.00053245355
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ lpdiblc2 = 7.1362462e-15
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ k2we = 5e-5
+ paigsd = 1.5255572e-23
+ dsub = 0.75
+ dtox = 2.7e-10
+ ku0we = -0.0007
+ bigbacc = 0.002588
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ beta0 = 13
+ leta0 = 2.6128654e-9
+ letab = -2.2297043e-8
+ permod = 1
+ kvth0we = 0.00018
+ ppclm = -2.5569374e-14
+ eta0 = 0.27220356
+ etab = -0.011678893
+ lkvth0we = -2e-12
+ dlcig = 2.5e-9
+ lintnoi = -1.5e-8
+ bgidl = 2320000000.0
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ acnqsmod = 0
+ voffcv = -0.16942
+ wpemod = 1
+ dmcgt = 0
+ tcjsw = 0.000357
+ rbodymod = 0
+ bigsd = 0.00125
+ ags = 2.5974722
+ wvoff = 8.241506600000007e-9
+ cjd = 0.00145199
+ cit = 1.5634930000000017e-5
+ cjs = 0.00145199
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 3.26497e-9
+ tpbswg = 0.0009
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ wvsat = -0.009212557199999995
+ nfactor = 1
+ wvth0 = -1.0705709100000002e-8
+ wpdiblc2 = 7.4309162e-10
+ waigc = -2.4473999e-12
+ la0 = 2.94419216e-8
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -8.998333e-5
+ kt1 = -0.41803712
+ lk2 = -5.0446112e-10
+ kt2 = -0.10268076
+ llc = 0
+ lln = 1
+ lu0 = 1.1446464e-10
+ mjd = 0.26
+ lua = 3.6827721e-17
+ mjs = 0.26
+ lub = -1.9895881809999996e-26
+ luc = 1.827009e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ ptvoff = -1.5034232e-16
+ njd = 1.02
+ njs = 1.02
+ pa0 = 7.627786000000002e-15
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 1.04787885e-9
+ pbs = 0.52
+ pk2 = 1.6131306e-16
+ waigsd = 3.0714121e-12
+ lketa = 2.8547804e-8
+ pu0 = -1.5881047e-16
+ prt = 0
+ pua = -1.4490045e-23
+ xpart = 1
+ pub = 2.3973370000000036e-34
+ puc = 4.0045874e-24
+ pud = 0
+ rsh = 17.5
+ keta = -0.51555907
+ tcj = 0.00076
+ ua1 = 9.0255397e-10
+ ub1 = -8.0270486e-19
+ uc1 = -7.4218809e-11
+ diomod = 1
+ tpb = 0.0014
+ nigbacc = 10
+ wa0 = 1.203209e-7
+ egidl = 0.29734
+ ute = -1
+ wat = -0.011948694
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -5.5751276e-9
+ pditsd = 0
+ pditsl = 0
+ wlc = 0
+ wln = 1
+ wkvth0we = 2e-12
+ wu0 = 1.3750374999999999e-9
+ cjswgd = 3.0174000000000004e-10
+ pku0we = -1.5e-18
+ xgl = -1.09e-8
+ cjswgs = 3.0174000000000004e-10
+ xgw = 0
+ wua = 1.5882075e-16
+ wub = -5.862147e-26
+ wuc = -7.6599643e-17
+ wud = 0
+ wwc = 0
+ jswd = 1.28e-13
+ wwl = 0
+ wwn = 1
+ jsws = 1.28e-13
+ lcit = 1.9165604e-10
+ kt1l = 0
+ trnqsmod = 0
+ nigbinv = 10
+ lint = 0
+ mjswgd = 0.85
+ mjswgs = 0.85
+ lkt1 = 1.0604028e-8
+ lkt2 = 1.0192413e-9
+ pvfbsdoff = 0
+ lmax = 8.833e-8
+ tcjswg = 0.001
+ lmin = 5.233e-8
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ minv = -0.3
+ rgatemod = 0
+ lua1 = -1.8750406e-17
+ wtvfbsdoff = 0
+ lub1 = -7.6940068e-27
+ luc1 = 1.062175e-17
+ pvoff = -1.8351133999999986e-16
+ tnjtsswg = 1
+ fnoimod = 1
+ ndep = 1e+18
+ eigbinv = 1.1
+ cdscb = 0
+ cdscd = 0
+ lwlc = 0
+ moin = 5.1
+ pvsat = 5.2995686e-10
+ wk2we = 5e-12
+ pvth0 = 3.3560707800000023e-16
+ ltvfbsdoff = 0
+ drout = 0.56
+ nigc = 3.083
+ paigc = 1.8938113e-18
+ fprout = 300
+ voffl = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ weta0 = -3.9858587e-8
+ wetab = 2.7041872e-8
+ lpclm = -8.5343289e-9
+ wtvoff = 1.7320676e-9
+ cigbacc = 0.32875
+ ntox = -0.31099999999999994
+ pcit = 5.3089970000000015e-18
+ pclm = 1.1824913
+ cgidl = 0.22
+ ptvfbsdoff = 0
+ tnoimod = 0
+ phin = 0.15
+ capmod = 2
+ pkt1 = -7.2165907e-15
+ pkt2 = -2.0869621e-15
+ wku0we = 2e-11
+ cigbinv = 0.006
+ pbswd = 0.8
+ pbsws = 0.8
+ mobmod = 0
+ rbdb = 50
+ pua1 = 1.2507395e-23
+ prwb = 0
+ prwg = 0
+ pub1 = -4.2778592e-33
+ puc1 = -7.7010123e-24
+ version = 4.5
+ pdits = 0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ cigsd = 0.069865
+ tempmod = 0
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ rdsw = 100
+ ijthsfwd = 0.01
+ aigbacc = 0.02
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ laigsd = -1.6939346e-18
+ tnoia = 0
+ ijthsrev = 0.01
+ rshg = 15.6
+ peta0 = 3.7467072e-15
+ aigbinv = 0.0163
+ petab = -3.4888335e-15
+ wketa = -1.1526014e-7
+ tpbsw = 0.0019
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ cjswd = 8.774000000000001e-11
+ cjsws = 8.774000000000001e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ ppdiblc2 = -4.5980291e-21
+ tnom = 25
+ toxe = 2.47e-9
+ toxm = 2.43e-9
+ )

.model nch_ss_15 nmos (
+ level = 54
+ fnoimod = 1
+ ltvoff = -2.8596488e-10
+ eigbinv = 1.1
+ pvfbsdoff = 0
+ lku0we = 2.5e-11
+ epsrox = 3.9
+ pvoff = 8.15540199999999e-16
+ cdscb = 0
+ cdscd = 0
+ rdsmod = 0
+ cigbacc = 0.32875
+ pvsat = -3.6390273e-9
+ igbmod = 1
+ wk2we = 5e-12
+ pvth0 = -5.048169999999999e-16
+ drout = 0.56
+ ijthsfwd = 0.01
+ paigc = 1.0773556e-18
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ tnoimod = 0
+ voffl = 0
+ pbswgd = 0.95
+ pbswgs = 0.95
+ keta = 0.067264197
+ cigbinv = 0.006
+ weta0 = 3.2678994e-7
+ igcmod = 1
+ wetab = -1.4667966e-7
+ lpclm = -8.0899178e-8
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 4.0133514e-10
+ ijthsrev = 0.01
+ kt1l = 0
+ cgidl = 0.22
+ version = 4.5
+ a0 = 5.6809619
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = -112965.493
+ cf = 7.5795e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = -0.012951152
+ k3 = -1.8419
+ em = 1000000.0
+ ll = 0
+ tempmod = 0
+ lw = 0
+ lint = 0
+ u0 = 0.0008145198599999999
+ w0 = 0
+ ua = -3.0786989e-9
+ ub = 2.197681248e-18
+ uc = -5.08518e-12
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 5.6700000000000005e-9
+ ww = 0
+ xw = 3.4e-9
+ lkt1 = -1.5973163e-8
+ lkt2 = 1.223943e-9
+ lmax = 5.233e-8
+ lmin = 4.333e-8
+ paigsd = -3.180948e-23
+ pbswd = 0.8
+ lpe0 = 9.2e-8
+ pbsws = 0.8
+ lpeb = 2.5e-7
+ aigbacc = 0.02
+ minv = -0.3
+ permod = 1
+ lua1 = 1.293984e-17
+ lub1 = 4.41313939e-26
+ luc1 = 1.702510023e-17
+ ndep = 1e+18
+ pdits = 0
+ lwlc = 0
+ cigsd = 0.069865
+ moin = 5.1
+ aigbinv = 0.0163
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ nigc = 3.083
+ voffcv = -0.16942
+ wpemod = 1
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ pkvth0we = -1.3e-19
+ tnoia = 0
+ ntox = -0.31099999999999994
+ pcit = 1.1838403e-17
+ pclm = 2.4301611
+ peta0 = -1.7518907e-14
+ petab = 6.5870154e-15
+ vfbsdoff = 0.02
+ wketa = 1.9475197e-7
+ poxedge = 1
+ tpbsw = 0.0019
+ phin = 0.15
+ cjswd = 8.774000000000001e-11
+ cjsws = 8.774000000000001e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ binunit = 2
+ pkt1 = 1.293618e-14
+ pkt2 = 7.7933247e-16
+ tpbswg = 0.0009
+ paramchk = 1
+ rbdb = 50
+ pua1 = -3.7208869e-24
+ prwb = 0
+ prwg = 0
+ pub1 = -7.551847900000001e-32
+ puc1 = -1.1133321e-23
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ ptvoff = 3.472697e-16
+ waigsd = 3.0722235e-12
+ rdsw = 100
+ ijthdfwd = 0.01
+ scref = 1e-6
+ diomod = 1
+ pigcd = 2.621
+ aigsd = 0.010772879
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ pditsd = 0
+ pditsl = 0
+ lvoff = -3.6979500799999987e-9
+ cjswgd = 3.0174000000000004e-10
+ pku0we = -1.5e-18
+ cjswgs = 3.0174000000000004e-10
+ tvfbsdoff = 0.022
+ lvsat = 0.0024201537900000003
+ ijthdrev = 0.01
+ lvth0 = 2.4529352400000003e-9
+ rshg = 15.6
+ delta = 0.007595625
+ laigc = -2.1310273e-11
+ wtvfbsdoff = 0
+ mjswgd = 0.85
+ mjswgs = 0.85
+ rnoia = 0
+ rnoib = 0
+ tcjswg = 0.001
+ ltvfbsdoff = 0
+ pketa = -9.5428465e-15
+ ngate = 8e+20
+ ngcon = 1
+ wpclm = -1.3405624e-6
+ njtsswg = 9
+ tnom = 25
+ wvfbsdoff = 0
+ gbmin = 1e-12
+ lvfbsdoff = 0
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ jswgd = 1.28e-13
+ toxe = 2.47e-9
+ jswgs = 1.28e-13
+ toxm = 2.43e-9
+ ckappad = 0.6
+ lkvth0we = -2e-12
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.0068331981
+ pdiblcb = -0.3
+ fprout = 300
+ ptvfbsdoff = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ acnqsmod = 0
+ wags = 1.2263301999999999e-6
+ wcit = -2.8590309999999997e-10
+ wtvoff = -6.84745e-9
+ bigbacc = 0.002588
+ rbodymod = 0
+ voff = -0.111418263
+ acde = 0.4
+ vsat = 81078.93740000001
+ tvoff = 0.0065547027
+ kvth0we = 0.00018
+ wint = 0
+ vth0 = 0.352586088
+ wkt1 = -2.6243076e-7
+ wkt2 = -3.3271248e-8
+ xjbvd = 1
+ xjbvs = 1
+ wmax = 9.0026e-6
+ lk2we = -1.5e-12
+ capmod = 2
+ aigc = 0.011691379
+ wmin = 9.025999999999999e-7
+ lintnoi = -1.5e-8
+ bigbinv = 0.004953
+ wku0we = 2e-11
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ mobmod = 0
+ ku0we = -0.0007
+ wua1 = 1.6438006e-16
+ wub1 = 1.23143716e-24
+ wuc1 = 1.56696984e-16
+ beta0 = 13
+ wpdiblc2 = 7.4301235e-10
+ leta0 = 1.0110619e-10
+ letab = 3.9727723e-8
+ bigc = 0.001442
+ wwlc = 0
+ ppclm = 7.229527e-14
+ cdsc = 0
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ cgbo = 0
+ cgdl = 3.0874977e-12
+ cgdo = 4.5622265999999996e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.0874977e-12
+ cgso = 4.5622265999999996e-11
+ cigc = 0.000625
+ laigsd = 3.532034e-18
+ dmcgt = 0
+ wkvth0we = 2e-12
+ tcjsw = 0.000357
+ nfactor = 1
+ ags = 2.5974722
+ trnqsmod = 0
+ cjd = 0.00145199
+ cit = -0.0035995337999999997
+ cjs = 0.00145199
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ dlc = 3.26497e-9
+ k3b = 1.9326
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ bigsd = 0.00125
+ k2we = 5e-5
+ wvoff = -8.983524000000003e-9
+ la0 = -3.0211764e-7
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = 0.0102832542
+ dsub = 0.75
+ kt1 = 0.040190302
+ lk2 = -1.6433965e-9
+ kt2 = -0.1062101
+ dtox = 2.7e-10
+ llc = 0
+ lln = 1
+ lu0 = 5.4830906e-10
+ mjd = 0.26
+ nigbacc = 10
+ lua = 7.492165e-17
+ mjs = 0.26
+ lub = -3.6402602300000003e-26
+ luc = 2.373596e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ wvsat = 0.062666402
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ njd = 1.02
+ njs = 1.02
+ pa0 = -1.230232e-13
+ rgatemod = 0
+ wvth0 = 3.784367999999988e-9
+ nsd = 1e+20
+ pbd = 0.52
+ pat = -9.3195589e-9
+ pbs = 0.52
+ pk2 = 5.8185614e-16
+ tnjtsswg = 1
+ pu0 = -6.648187499999999e-17
+ prt = 0
+ pua = 3.4306982e-23
+ pub = -6.0757564e-32
+ puc = -7.1571349e-24
+ pud = 0
+ waigc = 1.1629424e-11
+ eta0 = 0.31550975
+ rsh = 17.5
+ etab = -1.0810714
+ tcj = 0.00076
+ ua1 = 3.5617042e-10
+ ub1 = -1.696246019e-18
+ uc1 = -1.8462139999999999e-10
+ tpb = 0.0014
+ wa0 = 2.372924e-6
+ ute = -1
+ wat = 0.16680025
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -1.282587e-8
+ nigbinv = 10
+ lketa = -5.2559457e-9
+ toxref = 3e-9
+ wlc = 0
+ wln = 1
+ wu0 = -2.16836354e-10
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -6.825073e-16
+ wub = 9.9305604e-25
+ wuc = 1.1584384e-16
+ wud = 0
+ wwc = 0
+ xpart = 1
+ wwl = 0
+ wwn = 1
+ egidl = 0.29734
+ )

.model nch_ss_16 nmos (
+ level = 54
+ pketa = 8.7750313e-15
+ pkt1 = -9.3484796e-16
+ pkt2 = 1.5926682e-15
+ ngate = 8e+20
+ lku0we = 2.5e-11
+ ngcon = 1
+ wpclm = -1.03603352e-6
+ epsrox = 3.9
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ wpdiblc2 = 7.4301235e-10
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ rdsmod = 0
+ bigbacc = 0.002588
+ rbdb = 50
+ pua1 = -1.9060214e-23
+ prwb = 0
+ prwg = 0
+ pub1 = 5.2875851e-32
+ puc1 = 1.47310838e-23
+ igbmod = 1
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ rdsw = 100
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ kvth0we = 0.00018
+ pbswgd = 0.95
+ pbswgs = 0.95
+ lintnoi = -1.5e-8
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ igcmod = 1
+ wkvth0we = 2e-12
+ rshg = 15.6
+ trnqsmod = 0
+ tvoff = 0.002919136
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ paigsd = 4.3875156e-23
+ ku0we = -0.0007
+ permod = 1
+ beta0 = 13
+ rgatemod = 0
+ leta0 = 1.5743207e-8
+ tnom = 25
+ letab = 3.0329695e-8
+ tnjtsswg = 1
+ toxe = 2.47e-9
+ toxm = 2.43e-9
+ nfactor = 1
+ ppclm = 5.7373356e-14
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ voffcv = -0.16942
+ wpemod = 1
+ a0 = 3.2177147
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 155039.51
+ cf = 7.5795e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.027015951000000003
+ k3 = -1.8419
+ em = 1000000.0
+ ll = 0
+ lw = 0
+ ags = 2.5974722
+ u0 = 0.0038051123
+ w0 = 0
+ ua = -2.19661343e-9
+ ub = 1.4860819409999996e-18
+ uc = 2.2595638e-10
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ wags = 1.2263301999999999e-6
+ xl = 5.6700000000000005e-9
+ ww = 0
+ xw = 3.4e-9
+ cjd = 0.00145199
+ cit = -0.0016245269000000001
+ cjs = 0.00145199
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dmcgt = 0
+ dlc = 3.26497e-9
+ wcit = 3.3404264e-9
+ tcjsw = 0.000357
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ nigbacc = 10
+ voff = -0.04075972859999999
+ acde = 0.4
+ la0 = -1.8141853e-7
+ vsat = 96253.58170000001
+ wint = 0
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.0028489849000000005
+ vth0 = 0.34597836060000003
+ kt1 = -0.20813859
+ lk2 = -3.6017846e-9
+ kt2 = -0.11042259
+ llc = 0
+ lln = 1
+ lu0 = 4.0177003000000003e-10
+ wkt1 = 2.0651446e-8
+ wkt2 = -4.9869936e-8
+ mjd = 0.26
+ bigsd = 0.00125
+ lua = 3.1699464000000005e-17
+ mjs = 0.26
+ lub = -1.5342368999999952e-27
+ luc = -8.94744e-18
+ lud = 0
+ wmax = 9.0026e-6
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ aigc = 0.011397597
+ wmin = 9.025999999999999e-7
+ njs = 1.02
+ pa0 = -1.9996651e-13
+ nsd = 1e+20
+ nigbinv = 10
+ pbd = 0.52
+ pat = 1.3158901000000001e-9
+ pbs = 0.52
+ pk2 = 3.3250012e-16
+ tpbswg = 0.0009
+ pu0 = -1.22411747e-16
+ prt = 0
+ pua = 2.7971342e-23
+ pub = -4.5926045000000006e-32
+ puc = -7.6781524e-24
+ pud = 0
+ wvoff = 8.333983999999995e-9
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 4.3071269e-10
+ ub1 = -9.826436099999999e-20
+ uc1 = 5.294111900000001e-10
+ wua1 = 4.7742754e-16
+ tpb = 0.0014
+ wub1 = -1.3888553900000001e-24
+ wuc1 = -3.71148e-16
+ wvsat = 0.04358437799999999
+ wa0 = 3.9431957e-6
+ wvth0 = -2.2369996999999977e-8
+ ute = -1
+ wat = -0.050249687
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -7.7369724e-9
+ bigc = 0.001442
+ wlc = 0
+ wln = 1
+ wu0 = 9.245876399999999e-10
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -5.5320853e-16
+ wub = 6.903720200000001e-25
+ wuc = 1.2647685e-16
+ wud = 0
+ wwlc = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ waigc = -9.3979847e-11
+ ptvoff = -3.4317401e-17
+ waigsd = 3.0706789e-12
+ fnoimod = 1
+ cdsc = 0
+ eigbinv = 1.1
+ cgbo = 0
+ cgdl = 3.0874977e-12
+ cgdo = 4.5622265999999996e-11
+ xtid = 3
+ lketa = -2.4929909e-8
+ xtis = 3
+ ijthsfwd = 0.01
+ diomod = 1
+ cgsl = 3.0874977e-12
+ cgso = 4.5622265999999996e-11
+ xpart = 1
+ wtvfbsdoff = 0
+ cigc = 0.000625
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 3.0174000000000004e-10
+ pku0we = -1.5e-18
+ cjswgs = 3.0174000000000004e-10
+ egidl = 0.29734
+ ltvfbsdoff = 0
+ ijthsrev = 0.01
+ mjswgd = 0.85
+ mjswgs = 0.85
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ cigbacc = 0.32875
+ pvfbsdoff = 0
+ tcjswg = 0.001
+ tnoimod = 0
+ k2we = 5e-5
+ dsub = 0.75
+ dtox = 2.7e-10
+ ptvfbsdoff = 0
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ cigbinv = 0.006
+ pvoff = -3.3017380000000365e-17
+ cdscb = 0
+ cdscd = 0
+ eta0 = -0.003716791
+ etab = -0.88927493
+ pvsat = -2.7040040500000002e-9
+ wk2we = 5e-12
+ pvth0 = 7.767441600000001e-16
+ drout = 0.56
+ version = 4.5
+ fprout = 300
+ paigc = 6.2522098e-18
+ tempmod = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ voffl = 0
+ weta0 = 2.2378028e-8
+ pkvth0we = -1.3e-19
+ wetab = 3.831648e-8
+ aigbacc = 0.02
+ wtvoff = 9.4004181e-10
+ lpclm = -7.043921000000001e-8
+ cgidl = 0.22
+ vfbsdoff = 0.02
+ capmod = 2
+ aigbinv = 0.0163
+ wku0we = 2e-11
+ mobmod = 0
+ pbswd = 0.8
+ pbsws = 0.8
+ paramchk = 1
+ pdits = 0
+ cigsd = 0.069865
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ poxedge = 1
+ ijthdfwd = 0.01
+ laigsd = -2.6649547e-17
+ pk2we = -1e-19
+ keta = 0.46877367
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ binunit = 2
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ tnoia = 0
+ lcit = 3.0456022999999997e-10
+ ijthdrev = 0.01
+ kt1l = 0
+ peta0 = -2.6027237e-15
+ petab = -2.4777955e-15
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ wketa = -1.7908228e-7
+ tpbsw = 0.0019
+ lint = 0
+ cjswd = 8.774000000000001e-11
+ cjsws = 8.774000000000001e-11
+ lkt1 = -3.805047e-9
+ lkt2 = 1.4303548e-9
+ mjswd = 0.11
+ lmax = 4.333e-8
+ mjsws = 0.11
+ agidl = 9.41e-8
+ lmin = 3.6e-8
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ minv = -0.3
+ lua1 = 9.2872684e-18
+ lub1 = -3.4169731800000003e-26
+ luc1 = -1.796249619e-17
+ ndep = 1e+18
+ lwlc = 0
+ lkvth0we = -2e-12
+ moin = 5.1
+ toxref = 3e-9
+ nigc = 3.083
+ scref = 1e-6
+ pigcd = 2.621
+ aigsd = 0.01077288
+ acnqsmod = 0
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ lvoff = -7.160218279999998e-9
+ tvfbsdoff = 0.022
+ njtsswg = 9
+ rbodymod = 0
+ lvsat = 0.001676600613
+ lvth0 = 2.7767160299999994e-9
+ ntox = -0.31099999999999994
+ ltvoff = -1.0782211e-10
+ pcit = -1.6585171e-16
+ pclm = 2.21669238
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ delta = 0.007595625
+ laigc = -6.9149623e-12
+ ckappad = 0.6
+ ckappas = 0.6
+ rnoia = 0
+ rnoib = 0
+ pdiblc1 = 0
+ pdiblc2 = 0.0068331981
+ phin = 0.15
+ pdiblcb = -0.3
+ )

.model nch_ss_17 nmos (
+ level = 54
+ cgbo = 0
+ cgdl = 3.0874977e-12
+ cgdo = 4.5622265999999996e-11
+ xtid = 3
+ pbswgd = 0.95
+ xtis = 3
+ pbswgs = 0.95
+ ijthdfwd = 0.01
+ cgsl = 3.0874977e-12
+ cgso = 4.5622265999999996e-11
+ aigbinv = 0.0163
+ cigc = 0.000625
+ voffl = 0
+ igcmod = 1
+ weta0 = -1.09928e-7
+ wetab = 2.7482e-8
+ ijthdrev = 0.01
+ cgidl = 0.22
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ poxedge = 1
+ k2we = 5e-5
+ pbswd = 0.8
+ pbsws = 0.8
+ dsub = 0.75
+ permod = 1
+ dtox = 2.7e-10
+ binunit = 2
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ pdits = 0
+ eta0 = 0.42133333
+ cigsd = 0.069865
+ etab = -0.29033333
+ lkvth0we = -2e-12
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ voffcv = -0.16942
+ wpemod = 1
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ acnqsmod = 0
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ tnoia = 0
+ rbodymod = 0
+ peta0 = 0
+ wketa = -3.7974654e-8
+ tpbsw = 0.0019
+ cjswd = 8.774000000000001e-11
+ tpbswg = 0.0009
+ cjsws = 8.774000000000001e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ wtvfbsdoff = 0
+ a0 = 2.2098167
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 72000
+ cf = 7.5795e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.018686228
+ k3 = -1.8419
+ em = 1000000.0
+ wpdiblc2 = -6.449088e-9
+ ll = 0
+ lw = 0
+ u0 = 0.0159465
+ w0 = 0
+ ua = -1.7855187e-9
+ ub = 2.0636167e-18
+ uc = 7.8391667e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 5.6700000000000005e-9
+ ptvoff = 0
+ ww = 0
+ xw = 3.4e-9
+ njtsswg = 9
+ ltvfbsdoff = 0
+ waigsd = 3.0876027e-12
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ diomod = 1
+ scref = 1e-6
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.025656394
+ pigcd = 2.621
+ pdiblcb = -0.3
+ pditsd = 0
+ pditsl = 0
+ aigsd = 0.010772862
+ cjswgd = 3.0174000000000004e-10
+ pku0we = -1.5e-18
+ cjswgs = 3.0174000000000004e-10
+ keta = 0.015093331
+ tvfbsdoff = 0.022
+ lvoff = 0
+ wkvth0we = 2e-12
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lvsat = 0.0003
+ lcit = 4e-12
+ lvth0 = 0
+ ptvfbsdoff = 0
+ kt1l = 0
+ mjswgd = 0.85
+ mjswgs = 0.85
+ trnqsmod = 0
+ delta = 0.007595625
+ bigbacc = 0.002588
+ tcjswg = 0.001
+ rnoia = 0
+ rnoib = 0
+ lint = 6.5375218e-9
+ kvth0we = 0.00018
+ lkt1 = 0
+ lmax = 2.001e-5
+ lmin = 8.99743e-6
+ ngate = 8e+20
+ lintnoi = -1.5e-8
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ ngcon = 1
+ bigbinv = 0.004953
+ wpclm = 5.7423639e-7
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ rgatemod = 0
+ minv = -0.3
+ lub1 = 0
+ gbmin = 1e-12
+ tnjtsswg = 1
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ ndep = 1e+18
+ lwlc = 0
+ moin = 5.1
+ fprout = 300
+ nigc = 3.083
+ xrcrg1 = 12
+ xrcrg2 = 1
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ wtvoff = 9.3503662e-10
+ ntox = -0.31099999999999994
+ pcit = 0
+ pclm = 0.629885
+ tvoff = 5.0359625e-5
+ capmod = 2
+ nfactor = 1
+ wku0we = 2e-11
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ phin = 0.15
+ mobmod = 0
+ pkt1 = 0
+ ku0we = -0.0007
+ beta0 = 13
+ leta0 = 0
+ nigbacc = 10
+ rbdb = 50
+ prwb = 0
+ prwg = 0
+ pub1 = 0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ ags = 0.72720097
+ dlcig = 2.5e-9
+ rdsw = 100
+ bgidl = 2320000000.0
+ cjd = 0.00145199
+ cit = 6.2896875e-5
+ cjs = 0.00145199
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 9.8024918e-9
+ ijthsfwd = 0.01
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ nigbinv = 10
+ la0 = 0
+ jsd = 6.11e-7
+ dmcgt = 0
+ jss = 6.11e-7
+ lat = 0.0004
+ kt1 = -0.28314411
+ kt2 = -0.074391698
+ tcjsw = 0.000357
+ llc = 0
+ lln = 1
+ lu0 = -6e-12
+ mjd = 0.26
+ mjs = 0.26
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 0
+ ijthsrev = 0.01
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 6e-11
+ pbs = 0.52
+ rshg = 15.6
+ pu0 = 0
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ prt = 0
+ pud = 0
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = -6.8749055e-10
+ ub1 = 1.0341951e-18
+ uc1 = 4.5339833e-11
+ fnoimod = 1
+ bigsd = 0.00125
+ tpb = 0.0014
+ wa0 = 7.159061e-7
+ eigbinv = 1.1
+ ute = -2.01925
+ wat = 0
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 3.760485e-9
+ wlc = 0
+ wln = 1
+ wu0 = -1.03669e-10
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -7.132277e-17
+ wub = 7.28273e-26
+ wuc = -1.167985e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ wvoff = 1.0181215e-9
+ wvsat = -0.0045771271
+ wvth0 = -6.1727395e-9
+ tnom = 25
+ toxe = 2.47e-9
+ waigc = 5.0140497e-11
+ toxm = 2.43e-9
+ toxref = 3e-9
+ cigbacc = 0.32875
+ xpart = 1
+ tnoimod = 0
+ wags = 1.2493247e-7
+ egidl = 0.29734
+ pkvth0we = -1.3e-19
+ wcit = 4.4907306e-10
+ cigbinv = 0.006
+ voff = -0.11158375
+ ltvoff = 0
+ acde = 0.4
+ vsat = 106133.02
+ vfbsdoff = 0.02
+ wint = 0
+ pvfbsdoff = 0
+ vth0 = 0.37572953000000003
+ wkt1 = 3.5275480999999994e-8
+ wkt2 = 1.5939759e-8
+ wmax = 9.025999999999999e-7
+ aigc = 0.011740211
+ wmin = 5.426e-7
+ version = 4.5
+ tempmod = 0
+ lku0we = 2.5e-11
+ epsrox = 3.9
+ paramchk = 1
+ wua1 = 1.0731531e-15
+ wub1 = -9.2968455e-25
+ wuc1 = -1.4414309e-17
+ aigbacc = 0.02
+ rdsmod = 0
+ bigc = 0.001442
+ pvoff = -7e-17
+ wute = 5.565105e-7
+ wwlc = 0
+ igbmod = 1
+ cdscb = 0
+ cdscd = 0
+ pvsat = 0
+ wk2we = 5e-12
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ pvth0 = 2.3e-16
+ cdsc = 0
+ drout = 0.56
+ )

.model nch_ss_18 nmos (
+ level = 54
+ kt1l = 0
+ nigbacc = 10
+ tvoff = -0.0002433276
+ paigsd = 1.3573222e-22
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ lint = 6.5375218e-9
+ lkt1 = 8.6246405e-8
+ lkt2 = 5.1456509e-9
+ lmax = 8.99743e-6
+ lmin = 8.974099999999999e-7
+ permod = 1
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ nigbinv = 10
+ ags = 0.68161289
+ ku0we = -0.0007
+ ppdiblc2 = 1.9760389e-14
+ beta0 = 13
+ cjd = 0.00145199
+ leta0 = 0
+ cit = -0.00011782923
+ cjs = 0.00145199
+ minv = -0.3
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ lua1 = 1.38467e-15
+ lub1 = -1.4892591e-24
+ luc1 = 1.0686128e-16
+ dlc = 9.8024918e-9
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ ndep = 1e+18
+ lute = 1.0068051e-6
+ lwlc = 0
+ moin = 5.1
+ dlcig = 2.5e-9
+ voffcv = -0.16942
+ wpemod = 1
+ bgidl = 2320000000.0
+ la0 = -1.1479603e-6
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ nigc = 3.083
+ lat = 0.085745067
+ kt1 = -0.2927377
+ lk2 = -1.3507419e-8
+ kt2 = -0.074964073
+ llc = 0
+ lln = 1
+ lu0 = -2.0064396000000002e-9
+ fnoimod = 1
+ mjd = 0.26
+ lua = -1.5028094e-16
+ mjs = 0.26
+ lub = -1.4426347e-25
+ luc = -5.2935673e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = -5.1713984e-13
+ eigbinv = 1.1
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 6e-11
+ pbs = 0.52
+ pk2 = -1.6553107e-15
+ pu0 = 1.3573224e-17
+ prt = 0
+ noff = 2.7195
+ pua = -3.5916841e-23
+ pub = 6.5823852e-32
+ puc = 3.1761344e-23
+ pud = 0
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ pkvth0we = -1.3e-19
+ dmcgt = 0
+ rsh = 17.5
+ tcjsw = 0.000357
+ tcj = 0.00076
+ ua1 = -8.4151391e-10
+ ub1 = 1.1998524e-18
+ uc1 = 3.3453151e-11
+ tpb = 0.0014
+ wa0 = 7.7343e-7
+ pags = -1.4569295e-13
+ ute = -2.1312417
+ wtvfbsdoff = 0
+ wat = 0
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 3.944613e-9
+ wlc = 0
+ wln = 1
+ ntox = -0.31099999999999994
+ wu0 = -1.0517881e-10
+ pcit = -6.2947523e-16
+ xgl = -1.09e-8
+ pclm = 0.629885
+ xgw = 0
+ wua = -6.7327571e-17
+ wub = 6.5505403e-26
+ wuc = -1.5212814e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ vfbsdoff = 0.02
+ tpbswg = 0.0009
+ bigsd = 0.00125
+ ltvfbsdoff = 0
+ phin = 0.15
+ cigbacc = 0.32875
+ wvoff = 8.2208115e-10
+ pkt1 = -6.952314e-14
+ pkt2 = -1.5079533e-14
+ paramchk = 1
+ tnoimod = 0
+ wvsat = -0.0045771271
+ wvth0 = -6.4760901e-9
+ ptvoff = -2.0299898e-15
+ waigsd = 3.0875876e-12
+ waigc = 5.030718e-11
+ rbdb = 50
+ pua1 = -1.044071e-21
+ prwb = 0
+ prwg = 0
+ pub1 = 9.8799081e-31
+ cigbinv = 0.006
+ puc1 = -4.3746501e-23
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ pute = -5.4971558e-13
+ diomod = 1
+ rdsw = 100
+ ptvfbsdoff = 0
+ lketa = -1.3350472e-7
+ ijthdfwd = 0.01
+ pditsd = 0
+ xpart = 1
+ pditsl = 0
+ cjswgd = 3.0174000000000004e-10
+ pku0we = -1.5e-18
+ cjswgs = 3.0174000000000004e-10
+ version = 4.5
+ tempmod = 0
+ egidl = 0.29734
+ mjswgd = 0.85
+ mjswgs = 0.85
+ ijthdrev = 0.01
+ aigbacc = 0.02
+ a0 = 2.3375097
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ rshg = 15.6
+ at = 62506.667
+ cf = 7.5795e-11
+ tcjswg = 0.001
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.020188722
+ k3 = -1.8419
+ em = 1000000.0
+ pvfbsdoff = 0
+ ll = 0
+ lw = 0
+ u0 = 0.016169018
+ lpdiblc2 = -2.2119558e-8
+ w0 = 0
+ ua = -1.7688022e-9
+ ub = 2.0796638e-18
+ uc = 8.4279951e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 5.6700000000000005e-9
+ ww = 0
+ xw = 3.4e-9
+ aigbinv = 0.0163
+ tnom = 25
+ pvoff = 1.6924031e-15
+ toxe = 2.47e-9
+ toxm = 2.43e-9
+ cdscb = 0
+ cdscd = 0
+ fprout = 300
+ pvsat = 0
+ lkvth0we = -2e-12
+ wk2we = 5e-12
+ pvth0 = 2.9571226999999997e-15
+ drout = 0.56
+ xrcrg1 = 12
+ xrcrg2 = 1
+ paigc = -1.4984839e-18
+ voffl = 0
+ poxedge = 1
+ acnqsmod = 0
+ wtvoff = 1.1608419e-9
+ wags = 1.4113859e-7
+ weta0 = -1.09928e-7
+ wetab = 2.7482e-8
+ wcit = 5.1909255e-10
+ binunit = 2
+ rbodymod = 0
+ voff = -0.1094379
+ acde = 0.4
+ capmod = 2
+ cgidl = 0.22
+ vsat = 106133.02
+ wint = 0
+ wku0we = 2e-11
+ vth0 = 0.36994059
+ wkt1 = 4.3008867e-8
+ wkt2 = 1.7617127e-8
+ wmax = 9.025999999999999e-7
+ mobmod = 0
+ aigc = 0.011757817
+ wmin = 5.426e-7
+ pbswd = 0.8
+ pbsws = 0.8
+ wua1 = 1.1892901e-15
+ wub1 = -1.0395834e-24
+ wuc1 = -9.5481798e-18
+ wpdiblc2 = -8.647129e-9
+ bigc = 0.001442
+ wute = 6.1765795e-7
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ wwlc = 0
+ pdits = 0
+ cigsd = 0.069865
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ laigsd = -2.4859383e-16
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.0874977e-12
+ cgdo = 4.5622265999999996e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.0874977e-12
+ cgso = 4.5622265999999996e-11
+ cigc = 0.000625
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ wkvth0we = 2e-12
+ tnoia = 0
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ trnqsmod = 0
+ peta0 = 0
+ njtsswg = 9
+ wketa = -4.7550208e-8
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ tpbsw = 0.0019
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ cjswd = 8.774000000000001e-11
+ cjsws = 8.774000000000001e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.028116857
+ k2we = 5e-5
+ pdiblcb = -0.3
+ dsub = 0.75
+ dtox = 2.7e-10
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ rgatemod = 0
+ tnjtsswg = 1
+ toxref = 3e-9
+ eta0 = 0.42133333
+ etab = -0.29033333
+ bigbacc = 0.002588
+ scref = 1e-6
+ pigcd = 2.621
+ aigsd = 0.010772862
+ kvth0we = 0.00018
+ tvfbsdoff = 0.022
+ lvoff = -1.9291251e-8
+ lintnoi = -1.5e-8
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ ltvoff = 2.6402481e-9
+ lvsat = 0.0003
+ lvth0 = 5.2042566e-8
+ delta = 0.007595625
+ laigc = -1.5827875e-10
+ rnoia = 0
+ rnoib = 0
+ lku0we = 2.5e-11
+ pketa = 8.6084224e-14
+ epsrox = 3.9
+ ngate = 8e+20
+ ngcon = 1
+ wvfbsdoff = 0
+ wpclm = 5.7423639e-7
+ lvfbsdoff = 0
+ rdsmod = 0
+ gbmin = 1e-12
+ igbmod = 1
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ pbswgd = 0.95
+ pbswgs = 0.95
+ nfactor = 1
+ ijthsfwd = 0.01
+ igcmod = 1
+ keta = 0.029943688
+ lags = 4.0983681e-7
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 1.6287277e-9
+ ijthsrev = 0.01
+ )

.model nch_ss_19 nmos (
+ level = 54
+ rgatemod = 0
+ tnom = 25
+ tnjtsswg = 1
+ toxe = 2.47e-9
+ toxm = 2.43e-9
+ pdits = 0
+ cigsd = 0.069865
+ voffcv = -0.16942
+ wpemod = 1
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ njtsswg = 9
+ wtvfbsdoff = 0
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ ltvfbsdoff = 0
+ ckappad = 0.6
+ ckappas = 0.6
+ wags = -7.73542e-7
+ pdiblc1 = 0
+ pdiblc2 = -0.019237439
+ pdiblcb = -0.3
+ wcit = -4.5548514e-10
+ tnoia = 0
+ voff = -0.12566406
+ acde = 0.4
+ peta0 = 0
+ vsat = 106133.02
+ wketa = 9.2259042e-8
+ wint = 0
+ tpbswg = 0.0009
+ vth0 = 0.42814179
+ tpbsw = 0.0019
+ wkt1 = -6.8753249e-8
+ wkt2 = 3.7202325e-9
+ wmax = 9.025999999999999e-7
+ bigbacc = 0.002588
+ cjswd = 8.774000000000001e-11
+ aigc = 0.01160027
+ cjsws = 8.774000000000001e-11
+ wmin = 5.426e-7
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ ptvfbsdoff = 0
+ kvth0we = 0.00018
+ ptvoff = 9.96032e-16
+ wua1 = 1.1798319e-17
+ wub1 = 1.8760115e-25
+ wuc1 = -8.2926019e-17
+ lintnoi = -1.5e-8
+ waigsd = 3.0878745e-12
+ bigbinv = 0.004953
+ bigc = 0.001442
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ wwlc = 0
+ diomod = 1
+ cdsc = 0
+ cgbo = 0
+ pditsd = 0
+ pditsl = 0
+ cgdl = 3.0874977e-12
+ cgdo = 4.5622265999999996e-11
+ xtid = 3
+ xtis = 3
+ cjswgd = 3.0174000000000004e-10
+ ijthsfwd = 0.01
+ scref = 1e-6
+ pku0we = -1.5e-18
+ cjswgs = 3.0174000000000004e-10
+ cgsl = 3.0874977e-12
+ cgso = 4.5622265999999996e-11
+ cigc = 0.000625
+ pigcd = 2.621
+ tvfbsdoff = 0.022
+ aigsd = 0.010772861
+ lvoff = -4.8499703e-9
+ mjswgd = 0.85
+ mjswgs = 0.85
+ lvsat = 0.0003
+ lvth0 = 2.434924e-10
+ ijthsrev = 0.01
+ tcjswg = 0.001
+ delta = 0.007595625
+ laigc = -1.8062176e-11
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ rnoia = 0
+ rnoib = 0
+ nfactor = 1
+ pketa = -3.8346008e-14
+ ngate = 8e+20
+ k2we = 5e-5
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ ngcon = 1
+ dsub = 0.75
+ wpclm = 5.7423639e-7
+ dtox = 2.7e-10
+ ppdiblc2 = -1.3176269e-14
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ fprout = 300
+ eta0 = 0.42133333
+ etab = -0.29033333
+ xrcrg1 = 12
+ xrcrg2 = 1
+ nigbacc = 10
+ a0 = 1.6362276
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 209176.65
+ cf = 7.5795e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.016938797999999998
+ k3 = -1.8419
+ em = 1000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.015647274
+ w0 = 0
+ ua = -1.7708735e-9
+ ub = 1.8600147e-18
+ uc = 2.580063e-11
+ ud = 0
+ wtvoff = -2.2391826e-9
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 5.6700000000000005e-9
+ ww = 0
+ xw = 3.4e-9
+ pkvth0we = -1.3e-19
+ nigbinv = 10
+ capmod = 2
+ wku0we = 2e-11
+ tvoff = 0.004406442
+ vfbsdoff = 0.02
+ mobmod = 0
+ ags = 2.547561
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ cjd = 0.00145199
+ cit = 0.0020125208
+ cjs = 0.00145199
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 9.8024918e-9
+ k3b = 1.9326
+ fnoimod = 1
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ eigbinv = 1.1
+ paramchk = 1
+ ku0we = -0.0007
+ beta0 = 13
+ la0 = -5.2381924e-7
+ leta0 = 0
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.04479122
+ kt1 = -0.12585017
+ lk2 = -1.0614987e-8
+ kt2 = -0.061139846
+ llc = 0
+ lln = 1
+ lu0 = -1.5420873e-9
+ mjd = 0.26
+ lua = -1.4843753e-16
+ mjs = 0.26
+ lub = 5.1224193e-26
+ luc = -8.8907704e-19
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 9.5948774e-14
+ nsd = 1e+20
+ pbd = 0.52
+ pat = -4.9144129999999995e-9
+ pbs = 0.52
+ laigsd = 2.1900591e-16
+ pk2 = -1.0578878e-15
+ pu0 = 1.1957724e-17
+ dlcig = 2.5e-9
+ prt = 0
+ pua = 5.0063903e-23
+ pub = -8.0709098e-32
+ puc = -9.2074471e-24
+ pud = 0
+ bgidl = 2320000000.0
+ ijthdfwd = 0.01
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 7.2552224e-10
+ ub1 = -4.8701436e-19
+ uc1 = 1.8003493e-10
+ tpb = 0.0014
+ wa0 = 8.4566389e-8
+ ute = -1
+ wat = 0.0055892281
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 3.2733514e-9
+ keta = -0.17327473
+ cigbacc = 0.32875
+ wlc = 0
+ wln = 1
+ wu0 = -1.0336364000000001e-10
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -1.6393515e-16
+ wub = 2.3014917e-25
+ wuc = 3.0819536e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ dmcgt = 0
+ tcjsw = 0.000357
+ lags = -1.250857e-6
+ tnoimod = 0
+ jswd = 1.28e-13
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ jsws = 1.28e-13
+ lcit = -2.672838e-10
+ ijthdrev = 0.01
+ kt1l = 0
+ cigbinv = 0.006
+ lpdiblc2 = 2.0025765e-8
+ bigsd = 0.00125
+ lint = 6.5375218e-9
+ lkt1 = -6.2283496e-8
+ lkt2 = -7.1579117e-9
+ lmax = 8.974099999999999e-7
+ lmin = 4.4741e-7
+ wvoff = 5.2999378e-9
+ lpe0 = 9.2e-8
+ version = 4.5
+ lpeb = 2.5e-7
+ tempmod = 0
+ wvsat = -0.0045771271
+ wvth0 = -4.9199227000000006e-9
+ minv = -0.3
+ lua1 = -9.9922063e-18
+ lub1 = 1.2052288e-26
+ luc1 = -2.3596511e-17
+ toxref = 3e-9
+ waigc = 6.3350032e-11
+ ndep = 1e+18
+ aigbacc = 0.02
+ lwlc = 0
+ lkvth0we = -2e-12
+ moin = 5.1
+ lketa = 4.735968e-8
+ nigc = 3.083
+ xpart = 1
+ acnqsmod = 0
+ aigbinv = 0.0163
+ egidl = 0.29734
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ ltvoff = -1.4980468e-9
+ rbodymod = 0
+ pags = 6.6837277e-13
+ ntox = -0.31099999999999994
+ pvfbsdoff = 0
+ pcit = 2.3789891e-16
+ pclm = 0.629885
+ phin = 0.15
+ lku0we = 2.5e-11
+ epsrox = 3.9
+ pkt1 = 2.9945144e-14
+ pkt2 = -2.7112972e-15
+ poxedge = 1
+ rdsmod = 0
+ igbmod = 1
+ wpdiblc2 = 2.8360352e-8
+ pvoff = -2.2928893999999998e-15
+ binunit = 2
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ rbdb = 50
+ pua1 = 3.8966634e-24
+ prwb = 0
+ prwg = 0
+ pub1 = -1.0420346e-31
+ cdscb = 0
+ cdscd = 0
+ puc1 = 2.1559776e-23
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ pvsat = 0
+ rbsb = 50
+ pvag = 1.2
+ pbswgd = 0.95
+ pbswgs = 0.95
+ wk2we = 5e-12
+ pvth0 = 1.5721336999999999e-15
+ drout = 0.56
+ rdsw = 100
+ igcmod = 1
+ paigc = -1.3106622e-17
+ voffl = 0
+ weta0 = -1.09928e-7
+ wetab = 2.7482e-8
+ wkvth0we = 2e-12
+ trnqsmod = 0
+ cgidl = 0.22
+ rshg = 15.6
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ paigsd = -1.1957726e-22
+ permod = 1
+ pbswd = 0.8
+ pbsws = 0.8
+ )

.model nch_ss_20 nmos (
+ level = 54
+ rgatemod = 0
+ tnom = 25
+ tnjtsswg = 1
+ toxe = 2.47e-9
+ toxm = 2.43e-9
+ pdits = 0
+ cigsd = 0.069865
+ voffcv = -0.16942
+ wpemod = 1
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ njtsswg = 9
+ wtvfbsdoff = 0
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ ltvfbsdoff = 0
+ ckappad = 0.6
+ ckappas = 0.6
+ wags = 2.5246629999999998e-6
+ pdiblc1 = 0
+ pdiblc2 = 0.041730695
+ pdiblcb = -0.3
+ wcit = 1.5646633e-10
+ tnoia = 0
+ voff = -0.11119538
+ acde = 0.4
+ peta0 = 0
+ vsat = 99029.765
+ wketa = 8.4379468e-9
+ wint = 0
+ tpbswg = 0.0009
+ vth0 = 0.43649989
+ tpbsw = 0.0019
+ wkt1 = 1.1516763e-8
+ wkt2 = -6.4493333e-9
+ wmax = 9.025999999999999e-7
+ bigbacc = 0.002588
+ cjswd = 8.774000000000001e-11
+ aigc = 0.011620363
+ cjsws = 8.774000000000001e-11
+ wmin = 5.426e-7
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ ptvfbsdoff = 0
+ kvth0we = 0.00018
+ ptvoff = -1.0913215e-16
+ wua1 = 2.6150731e-17
+ wub1 = -7.4432483e-26
+ wuc1 = -3.5091334e-17
+ lintnoi = -1.5e-8
+ waigsd = 3.0877293e-12
+ bigbinv = 0.004953
+ bigc = 0.001442
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ wwlc = 0
+ diomod = 1
+ cdsc = 0
+ cgbo = 0
+ pditsd = 0
+ pditsl = 0
+ cgdl = 3.0874977e-12
+ cgdo = 4.5622265999999996e-11
+ xtid = 3
+ xtis = 3
+ cjswgd = 3.0174000000000004e-10
+ ijthsfwd = 0.01
+ scref = 1e-6
+ pku0we = -1.5e-18
+ cjswgs = 3.0174000000000004e-10
+ cgsl = 3.0874977e-12
+ cgso = 4.5622265999999996e-11
+ cigc = 0.000625
+ pigcd = 2.621
+ tvfbsdoff = 0.022
+ aigsd = 0.010772861
+ lvoff = -1.121619e-8
+ mjswgd = 0.85
+ mjswgs = 0.85
+ lvsat = 0.0034254309
+ lvth0 = -3.434068e-9
+ ijthsrev = 0.01
+ tcjswg = 0.001
+ delta = 0.007595625
+ laigc = -2.6902885e-11
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ rnoia = 0
+ rnoib = 0
+ nfactor = 1
+ pketa = -1.4647263e-15
+ ngate = 8e+20
+ k2we = 5e-5
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ ngcon = 1
+ dsub = 0.75
+ wpclm = 5.7423639e-7
+ dtox = 2.7e-10
+ ppdiblc2 = 1.3236303e-15
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ fprout = 300
+ eta0 = 0.42133333
+ etab = -0.29033333
+ xrcrg1 = 12
+ xrcrg2 = 1
+ nigbacc = 10
+ a0 = -0.63009793
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 152816.98
+ cf = 7.5795e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.01590817
+ k3 = -1.8419
+ em = 1000000.0
+ ll = -1.18e-13
+ lw = 0
+ u0 = 0.013570664999999999
+ w0 = 0
+ ua = -2.0345741e-9
+ ub = 2.0265059e-18
+ uc = 2.0750138e-11
+ ud = 0
+ wtvoff = 2.7255415e-10
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 5.6700000000000005e-9
+ ww = 0
+ xw = 3.4e-9
+ pkvth0we = -1.3e-19
+ nigbinv = 10
+ capmod = 2
+ wku0we = 2e-11
+ tvoff = 0.001369836
+ vfbsdoff = 0.02
+ mobmod = 0
+ ags = -5.4134702
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ cjd = 0.00145199
+ cit = 0.0010906361
+ cjs = 0.00145199
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 1.30529375e-8
+ k3b = 1.9326
+ fnoimod = 1
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ eigbinv = 1.1
+ paramchk = 1
+ ku0we = -0.0007
+ beta0 = 13
+ la0 = 4.73364e-7
+ leta0 = 0
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.019992964
+ kt1 = -0.257877
+ lk2 = -1.0161511e-8
+ kt2 = -0.061294719
+ llc = -1.18e-13
+ lln = 0.7
+ lu0 = -6.2837936e-10
+ mjd = 0.26
+ lua = -3.2409276e-17
+ mjs = 0.26
+ lub = -2.2031936e-26
+ luc = 1.3331392e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = -5.6835585e-13
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 5.5480901e-9
+ pbs = 0.52
+ laigsd = 6.148791e-17
+ pk2 = 5.7885716e-16
+ pu0 = 5.5708054e-18
+ dlcig = 2.5e-9
+ prt = 0
+ pua = 1.3198419e-23
+ pub = -1.7542132e-32
+ puc = -4.6237685e-24
+ pud = 0
+ bgidl = 2320000000.0
+ ijthdfwd = 0.01
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 7.2295613e-10
+ ub1 = -3.1143135e-19
+ uc1 = 1.5561971e-10
+ tpb = 0.0014
+ wa0 = 1.5943496e-6
+ ute = -1
+ wat = -0.018189188
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -4.4652352e-10
+ keta = -0.031454297
+ cigbacc = 0.32875
+ wlc = 0
+ wln = 1
+ wu0 = -8.884792000000001e-11
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -8.0149958e-17
+ wub = 8.6587882e-26
+ wuc = 2.0402085e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ dmcgt = 0
+ tcjsw = 0.000357
+ lags = 2.2519967e-6
+ tnoimod = 0
+ jswd = 1.28e-13
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ jsws = 1.28e-13
+ lcit = 1.3834545000000002e-10
+ ijthdrev = 0.01
+ kt1l = 0
+ cigbinv = 0.006
+ lpdiblc2 = -6.8002141e-9
+ bigsd = 0.00125
+ lint = 9.7879675e-9
+ lkt1 = -4.1916909e-9
+ lkt2 = -7.0897675e-9
+ lmax = 4.4741e-7
+ lmin = 2.1410000000000002e-7
+ wvoff = -5.5871857e-9
+ lpe0 = 9.2e-8
+ version = 4.5
+ lpeb = 2.5e-7
+ tempmod = 0
+ wvsat = 0.0018584193
+ wvth0 = -3.8953081e-9
+ minv = -0.3
+ lua1 = -8.8631172e-18
+ lub1 = -6.5204234e-26
+ luc1 = -1.2853813e-17
+ toxref = 3e-9
+ waigc = 3.2137522e-11
+ ndep = 1e+18
+ aigbacc = 0.02
+ lwlc = 0
+ lkvth0we = -2e-12
+ moin = 5.1
+ lketa = -1.5041313e-8
+ nigc = 3.083
+ xpart = 1
+ acnqsmod = 0
+ aigbinv = 0.0163
+ egidl = 0.29734
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ ltvoff = -1.6194017e-10
+ rbodymod = 0
+ pags = -7.8283743e-13
+ ntox = -0.31099999999999994
+ pvfbsdoff = 0
+ pcit = -3.1359735e-17
+ pclm = 0.629885
+ phin = 0.15
+ lku0we = 2.5e-11
+ epsrox = 3.9
+ pkt1 = -5.3736613e-15
+ pkt2 = 1.7633117e-15
+ poxedge = 1
+ rdsmod = 0
+ igbmod = 1
+ wpdiblc2 = -4.5939646e-9
+ pvoff = 2.497445e-15
+ binunit = 2
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ rbdb = 50
+ pua1 = -2.4183981e-24
+ prwb = 0
+ prwg = 0
+ pub1 = 1.1091342e-32
+ cdscb = 0
+ cdscd = 0
+ puc1 = 5.125141e-25
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ pvsat = -2.8316404e-9
+ rbsb = 50
+ pvag = 1.2
+ pbswgd = 0.95
+ pbswgs = 0.95
+ wk2we = 5e-12
+ pvth0 = 1.12130324e-15
+ drout = 0.56
+ rdsw = 100
+ igcmod = 1
+ paigc = 6.2688273e-19
+ voffl = 0
+ weta0 = -1.09928e-7
+ wetab = 2.7482e-8
+ wkvth0we = 2e-12
+ trnqsmod = 0
+ cgidl = 0.22
+ rshg = 15.6
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ paigsd = -5.5708045e-23
+ permod = 1
+ pbswd = 0.8
+ pbsws = 0.8
+ )

.model nch_ss_21 nmos (
+ level = 54
+ acnqsmod = 0
+ dmcgt = 0
+ version = 4.5
+ tcjsw = 0.000357
+ ptvfbsdoff = 0
+ tempmod = 0
+ rbodymod = 0
+ tpbswg = 0.0009
+ aigbacc = 0.02
+ bigsd = 0.00125
+ wvoff = 4.2089489999999885e-10
+ ptvoff = 6.7086074e-18
+ wvsat = -0.0116031636
+ waigsd = 3.0872445e-12
+ aigbinv = 0.0163
+ wvth0 = 1.0890214590000001e-8
+ wpdiblc2 = 3.4958017e-9
+ waigc = 1.7847398e-12
+ diomod = 1
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 3.0174000000000004e-10
+ pku0we = -1.5e-18
+ cjswgs = 3.0174000000000004e-10
+ lketa = -3.6124213e-8
+ xpart = 1
+ keta = 0.068466797
+ egidl = 0.29734
+ mjswgd = 0.85
+ mjswgs = 0.85
+ wkvth0we = 2e-12
+ poxedge = 1
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ tcjswg = 0.001
+ lcit = 6.5521194e-11
+ pvfbsdoff = 0
+ kt1l = 0
+ trnqsmod = 0
+ binunit = 2
+ lint = 9.7879675e-9
+ lkt1 = 7.1588252e-10
+ lkt2 = 9.4878496e-10
+ lmax = 2.1410000000000002e-7
+ lmin = 8.833e-8
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ rgatemod = 0
+ minv = -0.3
+ lua1 = 1.428412e-17
+ pvoff = 1.2297136100000002e-15
+ lub1 = -6.3260104e-26
+ luc1 = -5.9196014e-18
+ tnjtsswg = 1
+ fprout = 300
+ ndep = 1e+18
+ cdscb = 0
+ cdscd = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ pvsat = 8.752865999999776e-12
+ lwlc = 0
+ wk2we = 5e-12
+ pvth0 = -1.9984174400000003e-15
+ moin = 5.1
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ drout = 0.56
+ nigc = 3.083
+ paigc = 7.0313197e-18
+ wtvoff = -2.7645419e-10
+ voffl = 0
+ noff = 2.7195
+ weta0 = -1.09928e-7
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ wetab = 2.7482e-8
+ lpclm = 5.9671804e-8
+ capmod = 2
+ wku0we = 2e-11
+ ntox = -0.31099999999999994
+ cgidl = 0.22
+ pcit = -3.3161007e-17
+ pclm = 0.34708024
+ mobmod = 0
+ njtsswg = 9
+ phin = 0.15
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ pkt1 = -1.1050175e-15
+ pkt2 = -1.739649e-15
+ pbswd = 0.8
+ pbsws = 0.8
+ a0 = 1.2892878
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 51380.779
+ cf = 7.5795e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = -0.031282087
+ k3 = -1.8419
+ em = 1000000.0
+ ckappad = 0.6
+ ckappas = 0.6
+ ll = -1.18e-13
+ lw = 0
+ u0 = 0.011699764
+ w0 = 0
+ ua = -2.2703742e-9
+ ub = 2.053795462e-18
+ uc = 5.2246809e-11
+ ud = 0
+ pdiblc1 = 0
+ pdiblc2 = 0.010471563
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 5.6700000000000005e-9
+ ww = 0
+ xw = 3.4e-9
+ pdiblcb = -0.3
+ rbdb = 50
+ pua1 = -9.0422848e-24
+ prwb = 0
+ pdits = 0
+ laigsd = -6.8373623e-17
+ prwg = 0
+ pub1 = 1.3277736e-32
+ puc1 = 4.9546192e-24
+ cigsd = 0.069865
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ rdsw = 100
+ ijthsfwd = 0.01
+ bigbacc = 0.002588
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ kvth0we = 0.00018
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ tnoia = 0
+ ijthsrev = 0.01
+ lintnoi = -1.5e-8
+ bigbinv = 0.004953
+ peta0 = 0
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ rshg = 15.6
+ wketa = -5.2502872e-8
+ tpbsw = 0.0019
+ cjswd = 8.774000000000001e-11
+ cjsws = 8.774000000000001e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ ppdiblc2 = -3.8331042e-16
+ toxref = 3e-9
+ tnom = 25
+ toxe = 2.47e-9
+ toxm = 2.43e-9
+ scref = 1e-6
+ tvfbsdoff = 0.022
+ pigcd = 2.621
+ aigsd = 0.010772862
+ nfactor = 1
+ ltvoff = 9.6416574e-11
+ wags = -1.185467e-6
+ lvoff = -8.878213999999996e-10
+ pkvth0we = -1.3e-19
+ wcit = 1.6500316e-10
+ lvsat = 6.182528999999987e-5
+ lvth0 = -6.196310299999999e-9
+ voff = -0.16014500000000004
+ acde = 0.4
+ delta = 0.007595625
+ laigc = -1.4310771e-11
+ vfbsdoff = 0.02
+ vsat = 114971.1026
+ wint = 0
+ vth0 = 0.449591107
+ rnoia = 0
+ rnoib = 0
+ lku0we = 2.5e-11
+ wkt1 = -8.7137768e-9
+ wkt2 = 1.0152376e-8
+ nigbacc = 10
+ wmax = 9.025999999999999e-7
+ epsrox = 3.9
+ aigc = 0.011560684
+ wmin = 5.426e-7
+ wvfbsdoff = 0
+ pketa = 1.139354e-14
+ lvfbsdoff = 0
+ ngate = 8e+20
+ rdsmod = 0
+ ngcon = 1
+ paramchk = 1
+ wpclm = 8.9560432e-7
+ igbmod = 1
+ wua1 = 5.7543559e-17
+ wub1 = -8.4794537e-26
+ wuc1 = -5.6143964e-17
+ gbmin = 1e-12
+ nigbinv = 10
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ bigc = 0.001442
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ wwlc = 0
+ pbswgd = 0.95
+ pbswgs = 0.95
+ cdsc = 0
+ igcmod = 1
+ cgbo = 0
+ cgdl = 3.0874977e-12
+ cgdo = 4.5622265999999996e-11
+ xtid = 3
+ ijthdfwd = 0.01
+ xtis = 3
+ cgsl = 3.0874977e-12
+ cgso = 4.5622265999999996e-11
+ cigc = 0.000625
+ fnoimod = 1
+ eigbinv = 1.1
+ ags = 5.2595
+ ijthdrev = 0.01
+ cjd = 0.00145199
+ cit = 0.0014357747
+ cjs = 0.00145199
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 1.30529375e-8
+ paigsd = 4.6587859e-23
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ tvoff = 0.00014539643
+ lpdiblc2 = -2.045371e-10
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ permod = 1
+ la0 = 6.8373618e-8
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = 0.0014100743
+ kt1 = -0.28113564
+ lk2 = -2.0436616e-10
+ kt2 = -0.099392124
+ llc = -1.18e-13
+ lln = 0.7
+ wtvfbsdoff = 0
+ lu0 = -2.3361917e-10
+ mjd = 0.26
+ lua = 1.7344554e-17
+ mjs = 0.26
+ lub = -2.7790142600000004e-26
+ luc = -5.3126584e-18
+ lud = 0
+ k2we = 5e-5
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = -4.6587862e-14
+ nsd = 1e+20
+ dsub = 0.75
+ pbd = 0.52
+ pat = -1.7332973e-9
+ pbs = 0.52
+ pk2 = -1.7344476e-15
+ cigbacc = 0.32875
+ dtox = 2.7e-10
+ ku0we = -0.0007
+ pu0 = 3.028211e-18
+ beta0 = 13
+ prt = 0
+ pua = 1.2335294e-23
+ pub = -1.88032504e-32
+ puc = -1.1996375e-24
+ pud = 0
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ leta0 = 0
+ ltvfbsdoff = 0
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 6.1325358e-10
+ ub1 = -3.2064524e-19
+ uc1 = 1.2275615e-10
+ tnoimod = 0
+ tpb = 0.0014
+ ppclm = -6.7808634e-14
+ wa0 = -8.7848444e-7
+ voffcv = -0.16942
+ wpemod = 1
+ ute = -1
+ wat = 0.016319757
+ eta0 = 0.42133333
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 1.0517006e-8
+ lkvth0we = -2e-12
+ etab = -0.29033333
+ wlc = 0
+ wln = 1
+ wu0 = -7.6797711e-11
+ xgl = -1.09e-8
+ xgw = 0
+ dlcig = 2.5e-9
+ wua = -7.6059319e-17
+ wub = 9.256491399999999e-26
+ wuc = 4.1739756e-18
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ bgidl = 2320000000.0
+ cigbinv = 0.006
+ )

.model nch_ss_22 nmos (
+ level = 54
+ phin = 0.15
+ cjswd = 8.774000000000001e-11
+ cjsws = 8.774000000000001e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ pkt1 = -2.447551e-15
+ pkt2 = 8.0276583e-16
+ ptvoff = -9.1490879e-17
+ nfactor = 1
+ paramchk = 1
+ waigsd = 3.0879615e-12
+ diomod = 1
+ rbdb = 50
+ pua1 = -1.6477593e-25
+ prwb = 0
+ prwg = 0
+ pub1 = 1.4533022e-32
+ puc1 = 1.5607499999999994e-24
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ pditsd = 0
+ pditsl = 0
+ rbsb = 50
+ pvag = 1.2
+ cjswgd = 3.0174000000000004e-10
+ pku0we = -1.5e-18
+ cjswgs = 3.0174000000000004e-10
+ rdsw = 100
+ ijthdfwd = 0.01
+ scref = 1e-6
+ tvfbsdoff = 0.022
+ nigbacc = 10
+ pigcd = 2.621
+ aigsd = 0.010772861
+ mjswgd = 0.85
+ mjswgs = 0.85
+ lvoff = -4.968304999999992e-10
+ tcjswg = 0.001
+ lvsat = 0.0020364239840000003
+ ijthdrev = 0.01
+ lvth0 = 2.877403999999998e-10
+ nigbinv = 10
+ delta = 0.007595625
+ rshg = 15.6
+ laigc = -8.7106488e-12
+ lpdiblc2 = -4.1841324e-15
+ rnoia = 0
+ rnoib = 0
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ pketa = -2.7052976e-14
+ ngate = 8e+20
+ ngcon = 1
+ wpclm = 4.0103412e-7
+ fnoimod = 1
+ fprout = 300
+ eigbinv = 1.1
+ gbmin = 1e-12
+ tnom = 25
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ xrcrg1 = 12
+ xrcrg2 = 1
+ toxe = 2.47e-9
+ toxm = 2.43e-9
+ lkvth0we = -2e-12
+ wtvoff = 7.682212e-10
+ ags = 5.2595
+ cjd = 0.00145199
+ cit = 0.00012466993000000007
+ cjs = 0.00145199
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ acnqsmod = 0
+ dlc = 3.26497e-9
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ wags = -1.185467e-6
+ capmod = 2
+ wcit = -2.7211382e-10
+ cigbacc = 0.32875
+ rbodymod = 0
+ wku0we = 2e-11
+ la0 = -1.9182963e-7
+ voff = -0.164304478
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.00129425008
+ acde = 0.4
+ kt1 = -0.33033037
+ lk2 = -1.3785596e-9
+ kt2 = -0.066210327
+ mobmod = 0
+ llc = 0
+ lln = 1
+ lu0 = -3.5042418999999997e-11
+ tnoimod = 0
+ mjd = 0.26
+ tvoff = 0.00053139469
+ lua = 2.7860169e-17
+ mjs = 0.26
+ lub = -2.7395085e-26
+ luc = 1.41139916e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ vsat = 93964.74900000001
+ njs = 1.02
+ pa0 = 2.0809981e-13
+ wint = 0
+ vth0 = 0.38061184800000003
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 2.13894442e-9
+ pbs = 0.52
+ pk2 = 9.5324632e-16
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ wkt1 = 5.5684939e-9
+ wkt2 = -1.689459e-8
+ pu0 = -2.33571417e-17
+ wmax = 9.025999999999999e-7
+ prt = 0
+ pua = -6.3654423e-24
+ pub = 7.034010899999999e-33
+ puc = -7.127418999999999e-24
+ pud = 0
+ cigbinv = 0.006
+ aigc = 0.011501109
+ wmin = 5.426e-7
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 8.1588744e-10
+ ub1 = -6.9089562e-19
+ uc1 = 5.5536722999999985e-11
+ tpb = 0.0014
+ wa0 = -3.5879278e-6
+ ute = -1
+ wat = -0.024874303599999998
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -1.8075483e-8
+ ku0we = -0.0007
+ wlc = 0
+ wln = 1
+ wu0 = 2.03897552e-10
+ xgl = -1.09e-8
+ xgw = 0
+ beta0 = 13
+ wua = 1.2288469e-16
+ wub = -1.8229956900000002e-25
+ wua1 = -3.6898024e-17
+ wuc = 6.7235478e-17
+ wud = 0
+ wub1 = -9.8148649e-26
+ wuc1 = -2.0038907999999998e-17
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ leta0 = -1.0826782e-8
+ wpdiblc2 = -5.8202891e-10
+ letab = -2.2164189e-8
+ version = 4.5
+ bigc = 0.001442
+ laigsd = 3.8113519e-17
+ tempmod = 0
+ wwlc = 0
+ ppclm = -2.1319035e-14
+ dlcig = 2.5e-9
+ cdsc = 0
+ bgidl = 2320000000.0
+ cgbo = 0
+ cgdl = 3.0874977e-12
+ cgdo = 4.5622265999999996e-11
+ xtid = 3
+ aigbacc = 0.02
+ xtis = 3
+ cgsl = 3.0874977e-12
+ cgso = 4.5622265999999996e-11
+ cigc = 0.000625
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ dmcgt = 0
+ tcjsw = 0.000357
+ wkvth0we = 2e-12
+ aigbinv = 0.0163
+ a0 = 4.0574074
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 80150.18699999999
+ cf = 7.5795e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = -0.018790666999999997
+ k3 = -1.8419
+ em = 1000000.0
+ ll = 0
+ lw = 0
+ trnqsmod = 0
+ u0 = 0.009587245
+ w0 = 0
+ ua = -2.3822425e-9
+ ub = 2.049592666e-18
+ uc = -1.5441968e-10
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 5.6700000000000005e-9
+ ww = 0
+ xw = 3.4e-9
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ bigsd = 0.00125
+ wvoff = 3.044252900000001e-8
+ k2we = 5e-5
+ dsub = 0.75
+ dtox = 2.7e-10
+ wvsat = -0.020780859999999998
+ toxref = 3e-9
+ wvth0 = -3.2732843e-8
+ rgatemod = 0
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ tnjtsswg = 1
+ poxedge = 1
+ waigc = 1.9067031e-10
+ eta0 = 0.53651186
+ etab = -0.054544089
+ binunit = 2
+ lketa = 6.7720908e-8
+ xpart = 1
+ ltvoff = 6.0132739e-11
+ egidl = 0.29734
+ pvfbsdoff = 0
+ lku0we = 2.5e-11
+ epsrox = 3.9
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ rdsmod = 0
+ igbmod = 1
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ pvoff = -1.5923199999999998e-15
+ pbswgd = 0.95
+ pbswgs = 0.95
+ cdscb = 0
+ cdscd = 0
+ pvsat = 8.714606e-10
+ wk2we = 5e-12
+ igcmod = 1
+ pvth0 = 2.1021500000000004e-15
+ drout = 0.56
+ paigc = -1.0723924e-17
+ ijthsfwd = 0.01
+ njtsswg = 9
+ voffl = 0
+ keta = -1.0362685
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ weta0 = -2.7932191e-7
+ wetab = 6.5877739e-8
+ wtvfbsdoff = 0
+ lpclm = -1.3225653e-8
+ ckappad = 0.6
+ ckappas = 0.6
+ jswd = 1.28e-13
+ pdiblc1 = 0
+ jsws = 1.28e-13
+ pdiblc2 = 0.0082956805
+ lcit = 1.8876511000000002e-10
+ paigsd = -2.0809977e-23
+ pdiblcb = -0.3
+ ijthsrev = 0.01
+ kt1l = 0
+ cgidl = 0.22
+ ltvfbsdoff = 0
+ permod = 1
+ lint = 0
+ lkt1 = 5.3401869e-9
+ lkt2 = -2.1703039e-9
+ lmax = 8.833e-8
+ lmin = 5.233e-8
+ pbswd = 0.8
+ pbsws = 0.8
+ bigbacc = 0.002588
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ ppdiblc2 = 5.6582339e-21
+ minv = -0.3
+ kvth0we = 0.00018
+ lua1 = -4.7634626e-18
+ lub1 = -2.8456569e-26
+ luc1 = 3.9907281000000113e-19
+ voffcv = -0.16942
+ wpemod = 1
+ pdits = 0
+ ndep = 1e+18
+ lintnoi = -1.5e-8
+ cigsd = 0.069865
+ ptvfbsdoff = 0
+ lwlc = 0
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ moin = 5.1
+ vtsswgs = 4.2
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ nigc = 3.083
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ pkvth0we = -1.3e-19
+ tnoia = 0
+ tpbswg = 0.0009
+ peta0 = 1.5923028e-14
+ ntox = -0.31099999999999994
+ pcit = 7.928002500000001e-18
+ petab = -3.6091995e-15
+ pclm = 1.1225851
+ vfbsdoff = 0.02
+ wketa = 3.5650261e-7
+ tpbsw = 0.0019
+ )

.model nch_ss_23 nmos (
+ level = 54
+ pditsl = 0
+ cjswgd = 3.0174000000000004e-10
+ pku0we = -1.5e-18
+ cjswgs = 3.0174000000000004e-10
+ cdsc = 0
+ lketa = -2.0578185e-8
+ cgbo = 0
+ cgdl = 3.0874977e-12
+ cgdo = 4.5622265999999996e-11
+ ijthsfwd = 0.01
+ xtid = 3
+ xtis = 3
+ xpart = 1
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ cgsl = 3.0874977e-12
+ cgso = 4.5622265999999996e-11
+ cigc = 0.000625
+ mjswgd = 0.85
+ mjswgs = 0.85
+ egidl = 0.29734
+ tcjswg = 0.001
+ pvfbsdoff = 0
+ ijthsrev = 0.01
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ njtsswg = 9
+ k2we = 5e-5
+ dsub = 0.75
+ dtox = 2.7e-10
+ fprout = 300
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ xrcrg1 = 12
+ xrcrg2 = 1
+ pvoff = -3.995098540000001e-15
+ ckappad = 0.6
+ ckappas = 0.6
+ cdscb = 0
+ pdiblc1 = 0
+ pdiblc2 = 0.0082956083
+ cdscd = 0
+ pdiblcb = -0.3
+ pvsat = 3.857754111e-9
+ eta0 = 0.49180426
+ etab = -1.1686036
+ wk2we = 5e-12
+ pvth0 = 4.973404900000001e-15
+ drout = 0.56
+ wtvoff = -4.625476e-9
+ paigc = -1.7630641e-18
+ voffl = 0
+ weta0 = 1.6706711e-7
+ capmod = 2
+ bigbacc = 0.002588
+ wetab = -6.7375536e-8
+ pkvth0we = -1.3e-19
+ lpclm = -4.9784452e-8
+ wku0we = 2e-11
+ mobmod = 0
+ kvth0we = 0.00018
+ cgidl = 0.22
+ vfbsdoff = 0.02
+ lintnoi = -1.5e-8
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ pbswd = 0.8
+ pbsws = 0.8
+ paramchk = 1
+ laigsd = -3.1577826e-17
+ pdits = 0
+ cigsd = 0.069865
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ ijthdfwd = 0.01
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ keta = 0.48612964
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ nfactor = 1
+ tnoia = 0
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ ijthdrev = 0.01
+ lcit = 3.4212035e-10
+ peta0 = -9.9675358e-15
+ kt1l = 0
+ petab = 4.1194905e-15
+ wketa = -1.8474011e-7
+ tpbsw = 0.0019
+ lint = 0
+ cjswd = 8.774000000000001e-11
+ cjsws = 8.774000000000001e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ lkt1 = -1.4874128e-8
+ lkt2 = -1.4213753e-9
+ lmax = 5.233e-8
+ lmin = 4.333e-8
+ nigbacc = 10
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ toxref = 3e-9
+ minv = -0.3
+ lua1 = 7.7308837e-17
+ lub1 = -1.78071462e-25
+ luc1 = -1.2025833999999998e-17
+ ndep = 1e+18
+ lkvth0we = -2e-12
+ nigbinv = 10
+ lwlc = 0
+ moin = 5.1
+ a0 = 11.080765
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 31524.241299999994
+ cf = 7.5795e-11
+ ef = 1.0
+ k1 = 0.274
+ tvfbsdoff = 0.022
+ k2 = 0.015147898
+ k3 = -1.8419
+ em = 1000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.00027638826
+ scref = 1e-6
+ nigc = 3.083
+ w0 = 0
+ ua = -5.2066121e-9
+ ub = 5.20056154e-18
+ uc = 2.7090556e-10
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 5.6700000000000005e-9
+ ww = 0
+ xw = 3.4e-9
+ pigcd = 2.621
+ aigsd = 0.010772862
+ ltvoff = -1.4697355e-10
+ acnqsmod = 0
+ lvoff = 1.6118058999999991e-9
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ fnoimod = 1
+ lvsat = -0.0058544363700000004
+ rbodymod = 0
+ lvth0 = -3.5936672999999988e-9
+ eigbinv = 1.1
+ ntox = -0.31099999999999994
+ delta = 0.007595625
+ pcit = 6.5486977e-17
+ lku0we = 2.5e-11
+ pclm = 1.7529092
+ laigc = -1.8175152e-11
+ epsrox = 3.9
+ rnoia = 0
+ rnoib = 0
+ wvfbsdoff = 0
+ phin = 0.15
+ lvfbsdoff = 0
+ rdsmod = 0
+ pketa = 4.339103e-15
+ igbmod = 1
+ ngate = 8e+20
+ pkt1 = 1.1940455e-14
+ pkt2 = 3.1759909e-15
+ ngcon = 1
+ wpclm = -7.2697212e-7
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ wpdiblc2 = -5.8193135e-10
+ pbswgd = 0.95
+ gbmin = 1e-12
+ pbswgs = 0.95
+ cigbacc = 0.32875
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ ags = 5.2595
+ rbdb = 50
+ pua1 = -6.2039198e-23
+ prwb = 0
+ prwg = 0
+ pub1 = 1.25797289e-31
+ puc1 = 1.5186895599999997e-23
+ igcmod = 1
+ wtvfbsdoff = 0
+ cjd = 0.00145199
+ cit = -0.0025193893
+ cjs = 0.00145199
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ dlc = 3.26497e-9
+ k3b = 1.9326
+ tnoimod = 0
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ rdsw = 100
+ ltvfbsdoff = 0
+ cigbinv = 0.006
+ la0 = -5.9918439e-7
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = 0.0015260548200000004
+ kt1 = 0.018192305
+ lk2 = -3.3469964e-9
+ kt2 = -0.079122889
+ llc = 0
+ lln = 1
+ lu0 = 5.0498706e-10
+ mjd = 0.26
+ lua = 1.9167361e-16
+ mjs = 0.26
+ lub = -2.101512744e-25
+ luc = -1.0554871600000002e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 1.4611928e-13
+ wkvth0we = 2e-12
+ nsd = 1e+20
+ pbd = 0.52
+ pat = -1.3855335799999999e-9
+ pbs = 0.52
+ pk2 = 2.1253177e-15
+ paigsd = 1.0451534e-29
+ pu0 = -2.7232224e-17
+ prt = 0
+ pua = -7.1470289e-23
+ pub = 9.665873609999999e-32
+ puc = 4.556057900000002e-24
+ pud = 0
+ version = 4.5
+ rsh = 17.5
+ trnqsmod = 0
+ tcj = 0.00076
+ ua1 = -5.9915221e-10
+ ub1 = 1.88867097e-18
+ uc1 = 2.697591899999999e-10
+ rshg = 15.6
+ tempmod = 0
+ tvoff = 0.0041021928
+ tpb = 0.0014
+ wa0 = -2.5192978e-6
+ permod = 1
+ ute = -1
+ wat = 0.035892558
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -3.8283609e-8
+ xjbvd = 1
+ xjbvs = 1
+ wlc = 0
+ wln = 1
+ lk2we = -1.5e-12
+ wu0 = 2.7070790000000004e-10
+ xgl = -1.09e-8
+ xgw = 0
+ wua = 1.2453821e-15
+ wub = -1.72755342e-24
+ wuc = -1.3420376999999993e-16
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ ptvfbsdoff = 0
+ aigbacc = 0.02
+ ku0we = -0.0007
+ beta0 = 13
+ rgatemod = 0
+ leta0 = -8.2337409e-9
+ letab = 4.245126e-8
+ voffcv = -0.16942
+ wpemod = 1
+ tnom = 25
+ tnjtsswg = 1
+ toxe = 2.47e-9
+ toxm = 2.43e-9
+ aigbinv = 0.0163
+ ppclm = 4.4105328e-14
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ wags = -1.185467e-6
+ dmcgt = 0
+ tcjsw = 0.000357
+ wcit = -1.26451726e-9
+ tpbswg = 0.0009
+ voff = -0.20066027000000003
+ acde = 0.4
+ poxedge = 1
+ vsat = 230014.02399999995
+ wint = 0
+ vth0 = 0.44753267
+ bigsd = 0.00125
+ binunit = 2
+ wkt1 = -2.4250058e-7
+ wkt2 = -5.7812263e-8
+ wmax = 9.025999999999999e-7
+ aigc = 0.01166429
+ wmin = 5.426e-7
+ ptvoff = 2.2134356e-16
+ wvoff = 7.186973409999998e-8
+ waigsd = 3.0876027e-12
+ wvsat = -0.07226864247
+ wua1 = 1.0299024e-15
+ wub1 = -2.01649781e-24
+ wuc1 = -2.54972289e-16
+ wvth0 = -8.223723199999997e-8
+ diomod = 1
+ bigc = 0.001442
+ waigc = 3.6172725e-11
+ wwlc = 0
+ pditsd = 0
+ )

.model nch_ss_24 nmos (
+ level = 54
+ lvsat = -0.0033603521999999992
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lvth0 = 5.278952700000001e-9
+ lcit = 2.3309058e-10
+ trnqsmod = 0
+ kt1l = 0
+ cigbacc = 0.32875
+ delta = 0.007595625
+ laigc = -7.4258513e-12
+ rnoia = 0
+ rnoib = 0
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ tnoimod = 0
+ lint = 0
+ lkt1 = 1.0114149e-9
+ lkt2 = 6.4873536e-9
+ lmax = 4.333e-8
+ pketa = 3.05233408e-14
+ ags = 5.2595
+ ngate = 8e+20
+ lmin = 3.6e-8
+ cigbinv = 0.006
+ ngcon = 1
+ lpe0 = 9.2e-8
+ cjd = 0.00145199
+ cit = -0.0002942959999999999
+ fprout = 300
+ cjs = 0.00145199
+ clc = 1e-7
+ wpclm = 9.524622100000001e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ lpeb = 2.5e-7
+ dlc = 3.26497e-9
+ k3b = 1.9326
+ xrcrg1 = 12
+ xrcrg2 = 1
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ rgatemod = 0
+ gbmin = 1e-12
+ minv = -0.3
+ tnjtsswg = 1
+ lua1 = -6.7547343e-17
+ lub1 = 1.43021154e-25
+ luc1 = 6.782260000000001e-18
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ ndep = 1e+18
+ la0 = -5.581062559999999e-7
+ version = 4.5
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.00127504779
+ wtvoff = -5.6534448e-10
+ lwlc = 0
+ kt1 = -0.30600245
+ lk2 = -3.4047834e-9
+ kt2 = -0.24052552
+ llc = 0
+ moin = 5.1
+ lln = 1
+ lu0 = 7.0945495e-10
+ tempmod = 0
+ mjd = 0.26
+ lua = 1.9963428e-16
+ mjs = 0.26
+ lub = -1.86515944e-25
+ luc = -1.3855022100000003e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 1.41312605e-13
+ nigc = 3.083
+ nsd = 1e+20
+ pbd = 0.52
+ pat = -1.1010081000000005e-10
+ pbs = 0.52
+ pk2 = 1.540171e-16
+ pu0 = -4.0117431000000003e-16
+ prt = 0
+ pua = -1.24177601e-22
+ pub = 1.2166737845000001e-31
+ puc = -3.231882900000001e-24
+ pud = 0
+ aigbacc = 0.02
+ capmod = 2
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 2.3570964e-9
+ ub1 = -4.6642377000000004e-18
+ uc1 = -1.1408099999999994e-10
+ tpb = 0.0014
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ wku0we = 2e-11
+ wa0 = -2.4212027299999997e-6
+ ute = -1
+ wat = 0.009863318999999999
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 1.947015e-9
+ wlc = 0
+ wln = 1
+ wu0 = 7.902177499999999e-9
+ xgl = -1.09e-8
+ mobmod = 0
+ xgw = 0
+ wua = 2.32104147e-15
+ wub = -2.2379339299999998e-24
+ wuc = 2.4733810000000014e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ ntox = -0.31099999999999994
+ pcit = -1.0110125699999999e-16
+ pclm = 0.021884800000000038
+ tvoff = 0.0045807103
+ aigbinv = 0.0163
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ phin = 0.15
+ pkt1 = -5.2985624e-15
+ pkt2 = -2.9889728e-15
+ ku0we = -0.0007
+ beta0 = 13
+ laigsd = 2.1777751e-17
+ leta0 = 6.023777099999999e-9
+ letab = 3.2196399e-8
+ ppclm = -3.8186956000000005e-14
+ rbdb = 50
+ pua1 = 5.0551945e-23
+ prwb = 0
+ prwg = 0
+ pub1 = -1.0765901599999999e-31
+ puc1 = -7.6876879e-24
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ poxedge = 1
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ rdsw = 100
+ ijthsfwd = 0.01
+ binunit = 2
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ dmcgt = 0
+ tcjsw = 0.000357
+ ijthsrev = 0.01
+ rshg = 15.6
+ bigsd = 0.00125
+ wvoff = -4.371822099999998e-8
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ toxref = 3e-9
+ wvsat = -0.03148762100000001
+ wvth0 = 4.9674833e-8
+ tnom = 25
+ waigc = -1.3685053e-10
+ toxe = 2.47e-9
+ toxm = 2.43e-9
+ lketa = -4.89346675e-8
+ xpart = 1
+ ltvoff = -1.7042091e-10
+ egidl = 0.29734
+ njtsswg = 9
+ wags = -1.185467e-6
+ pkvth0we = -1.3e-19
+ pvfbsdoff = 0
+ wcit = 2.1352386e-9
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ voff = 0.016693055000000012
+ lku0we = 2.5e-11
+ acde = 0.4
+ ckappad = 0.6
+ epsrox = 3.9
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.0082956083
+ vfbsdoff = 0.02
+ pdiblcb = -0.3
+ vsat = 179114.496
+ wint = 0
+ vth0 = 0.266458765
+ wkt1 = 1.0931611e-7
+ wkt2 = 6.8003321e-8
+ rdsmod = 0
+ wtvfbsdoff = 0
+ wmax = 9.025999999999999e-7
+ aigc = 0.011444916
+ wmin = 5.426e-7
+ igbmod = 1
+ a0 = 10.24243689
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 88689.602
+ cf = 7.5795e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.016327223000000002
+ k3 = -1.8419
+ em = 1000000.0
+ ll = 0
+ lw = 0
+ u0 = -0.0038964158
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ paramchk = 1
+ w0 = 0
+ ua = -5.369074800000001e-9
+ ub = 4.718207719999999e-18
+ uc = 3.3825556e-10
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 5.6700000000000005e-9
+ ww = 0
+ xw = 3.4e-9
+ ltvfbsdoff = 0
+ pbswgd = 0.95
+ pbswgs = 0.95
+ wua1 = -1.2678761e-15
+ wub1 = 2.74791671e-24
+ wuc1 = 2.1185608000000002e-16
+ bigbacc = 0.002588
+ pvoff = 1.6687133299999993e-15
+ bigc = 0.001442
+ igcmod = 1
+ wwlc = 0
+ cdscb = 0
+ cdscd = 0
+ kvth0we = 0.00018
+ pvsat = 1.85948003e-9
+ wk2we = 5e-12
+ pvth0 = -1.4902817e-15
+ drout = 0.56
+ cdsc = 0
+ lintnoi = -1.5e-8
+ paigc = 6.7150752e-18
+ cgbo = 0
+ ijthdfwd = 0.01
+ cgdl = 3.0874977e-12
+ cgdo = 4.5622265999999996e-11
+ xtid = 3
+ xtis = 3
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ cgsl = 3.0874977e-12
+ cgso = 4.5622265999999996e-11
+ voffl = 0
+ cigc = 0.000625
+ ptvfbsdoff = 0
+ weta0 = -1.6294544599999998e-7
+ wetab = 1.0177792e-7
+ paigsd = 4.9710031e-30
+ lpclm = 3.5035747999999996e-8
+ ijthdrev = 0.01
+ cgidl = 0.22
+ permod = 1
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ pbswd = 0.8
+ pbsws = 0.8
+ k2we = 5e-5
+ dsub = 0.75
+ dtox = 2.7e-10
+ voffcv = -0.16942
+ wpemod = 1
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ nfactor = 1
+ pdits = 0
+ cigsd = 0.069865
+ eta0 = 0.20083450200000003
+ lkvth0we = -2e-12
+ etab = -0.95932067
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ acnqsmod = 0
+ nigbacc = 10
+ tpbswg = 0.0009
+ tnoia = 0
+ rbodymod = 0
+ peta0 = 6.20307972e-15
+ petab = -4.1690291e-15
+ wketa = -7.1911233e-7
+ tpbsw = 0.0019
+ nigbinv = 10
+ cjswd = 8.774000000000001e-11
+ cjsws = 8.774000000000001e-11
+ ptvoff = 2.2397114e-17
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ waigsd = 3.0876027e-12
+ diomod = 1
+ wpdiblc2 = -5.8193135e-10
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 3.0174000000000004e-10
+ pku0we = -1.5e-18
+ fnoimod = 1
+ cjswgs = 3.0174000000000004e-10
+ eigbinv = 1.1
+ tvfbsdoff = 0.022
+ scref = 1e-6
+ pigcd = 2.621
+ mjswgd = 0.85
+ aigsd = 0.010772861
+ mjswgs = 0.85
+ keta = 1.06483334
+ tcjswg = 0.001
+ lvoff = -9.038509000000001e-9
+ wkvth0we = 2e-12
+ )

.model nch_ss_25 nmos (
+ level = 54
+ fprout = 300
+ xrcrg1 = 12
+ xrcrg2 = 1
+ pvoff = -7e-17
+ tnom = 25
+ cdscb = 0
+ cdscd = 0
+ toxe = 2.47e-9
+ toxm = 2.43e-9
+ wtvoff = 0
+ pvsat = 0
+ lkvth0we = -2e-12
+ wk2we = 5e-12
+ pvth0 = 2.3e-16
+ drout = 0.56
+ voffl = 0
+ capmod = 2
+ acnqsmod = 0
+ wku0we = 2e-11
+ weta0 = -1.1162667e-8
+ wags = -5.5469040000000005e-8
+ wetab = 2.2325333e-8
+ mobmod = 0
+ wcit = 2.963688e-10
+ rbodymod = 0
+ nfactor = 1
+ voff = -0.13478422
+ acde = 0.4
+ cgidl = 0.22
+ vsat = 102889.02
+ wint = 0
+ vth0 = 0.39220512
+ wkt1 = 1.102940613e-9
+ wkt2 = -5.3296152e-9
+ wmax = 5.426e-7
+ aigc = 0.011779434
+ wmin = 2.726e-7
+ pbswd = 0.8
+ pbsws = 0.8
+ wua1 = -1.874362e-16
+ nigbacc = 10
+ wub1 = 1.1464267e-25
+ wuc1 = -2.7527136e-17
+ wpdiblc2 = 4.9914968e-9
+ bigc = 0.001442
+ pdits = 0
+ wwlc = 0
+ cigsd = 0.069865
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.0874977e-12
+ cgdo = 4.5622265999999996e-11
+ xtid = 3
+ nigbinv = 10
+ xtis = 3
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ cgsl = 3.0874977e-12
+ cgso = 4.5622265999999996e-11
+ cigc = 0.000625
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ wkvth0we = 2e-12
+ tnoia = 0
+ trnqsmod = 0
+ peta0 = 0
+ fnoimod = 1
+ wketa = 1.6322115e-8
+ eigbinv = 1.1
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ tpbsw = 0.0019
+ dmdg = 0
+ cjswd = 8.774000000000001e-11
+ cjsws = 8.774000000000001e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ toxref = 3e-9
+ k2we = 5e-5
+ dsub = 0.75
+ dtox = 2.7e-10
+ rgatemod = 0
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ tnjtsswg = 1
+ tvfbsdoff = 0.022
+ eta0 = 0.24044444
+ etab = -0.28088889
+ cigbacc = 0.32875
+ ltvoff = 0
+ scref = 1e-6
+ pigcd = 2.621
+ tnoimod = 0
+ aigsd = 0.010772818
+ wtvfbsdoff = 0
+ lvoff = 0
+ cigbinv = 0.006
+ lvsat = 0.0003
+ lku0we = 2.5e-11
+ lvth0 = 0
+ ltvfbsdoff = 0
+ epsrox = 3.9
+ delta = 0.007595625
+ ags = 1.05760667
+ wvfbsdoff = 0
+ cjd = 0.00145199
+ cit = 0.000342575
+ version = 4.5
+ cjs = 0.00145199
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ lvfbsdoff = 0
+ rnoia = 0
+ rnoib = 0
+ rdsmod = 0
+ dlc = 9.8024918e-9
+ k3b = 1.9326
+ tempmod = 0
+ igbmod = 1
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ ngate = 8e+20
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ ngcon = 1
+ la0 = 0
+ wpclm = 9.3989653e-8
+ pbswgd = 0.95
+ jsd = 6.11e-7
+ pbswgs = 0.95
+ jss = 6.11e-7
+ lat = 0.0004
+ aigbacc = 0.02
+ kt1 = -0.22055704
+ kt2 = -0.0354368
+ llc = 0
+ lln = 1
+ lu0 = -6e-12
+ mjd = 0.26
+ mjs = 0.26
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ gbmin = 1e-12
+ njs = 1.02
+ pa0 = 0
+ igcmod = 1
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 6e-11
+ jswgd = 1.28e-13
+ ptvfbsdoff = 0
+ pbs = 0.52
+ jswgs = 1.28e-13
+ pu0 = 0
+ prt = 0
+ pud = 0
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 1.6212811e-9
+ ub1 = -8.7849211e-19
+ uc1 = 6.9356e-11
+ tpb = 0.0014
+ aigbinv = 0.0163
+ wa0 = -1.17208e-8
+ ijthsfwd = 0.01
+ ute = -1
+ wat = 0.071441067
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 1.8596306e-9
+ wlc = 0
+ wln = 1
+ wu0 = -1.2637067000000002e-9
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -1.3097991e-16
+ wub = 9.54408e-26
+ wuc = -2.4557867e-18
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ keta = -0.084351302
+ a0 = 3.5424667
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = -58844.444
+ cf = 7.5795e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.022167646
+ k3 = -1.8419
+ em = 1000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.018071111
+ jswd = 1.28e-13
+ w0 = 0
+ jsws = 1.28e-13
+ ijthsrev = 0.01
+ ua = -1.6762565e-9
+ ub = 2.0222e-18
+ uc = 6.1497778e-11
+ ud = 0
+ lcit = 4e-12
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 5.6700000000000005e-9
+ ww = 0
+ xw = 3.4e-9
+ permod = 1
+ kt1l = 0
+ tvoff = 0.0017628809
+ xjbvd = 1
+ xjbvs = 1
+ poxedge = 1
+ lk2we = -1.5e-12
+ lint = 6.5375218e-9
+ lkt1 = 0
+ lmax = 2.001e-5
+ binunit = 2
+ lmin = 8.99743e-6
+ lpe0 = 9.2e-8
+ voffcv = -0.16942
+ wpemod = 1
+ lpeb = 2.5e-7
+ ku0we = -0.0007
+ beta0 = 13
+ leta0 = 0
+ minv = -0.3
+ lub1 = 0
+ ndep = 1e+18
+ lwlc = 0
+ dlcig = 2.5e-9
+ moin = 5.1
+ bgidl = 2320000000.0
+ nigc = 3.083
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ noff = 2.7195
+ dmcgt = 0
+ noia = 3.11e+42
+ noib = 1.22e+22
+ pkvth0we = -1.3e-19
+ noic = 45200000.0
+ tpbswg = 0.0009
+ tcjsw = 0.000357
+ ntox = -0.31099999999999994
+ pcit = 0
+ pclm = 1.5094578
+ vfbsdoff = 0.02
+ bigsd = 0.00125
+ ptvoff = 0
+ phin = 0.15
+ waigsd = 3.1112026e-12
+ wvoff = 1.3685577e-8
+ pkt1 = 0
+ paramchk = 1
+ diomod = 1
+ wvsat = -0.0028059037
+ wvth0 = -1.5168414e-8
+ njtsswg = 9
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 3.0174000000000004e-10
+ pku0we = -1.5e-18
+ cjswgs = 3.0174000000000004e-10
+ waigc = 2.8724444e-11
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ rbdb = 50
+ prwb = 0
+ prwg = 0
+ pub1 = 0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.0047029422
+ rdsw = 100
+ pdiblcb = -0.3
+ ijthdfwd = 0.01
+ mjswgd = 0.85
+ xpart = 1
+ mjswgs = 0.85
+ tcjswg = 0.001
+ egidl = 0.29734
+ pvfbsdoff = 0
+ bigbacc = 0.002588
+ ijthdrev = 0.01
+ rshg = 15.6
+ kvth0we = 0.00018
+ lintnoi = -1.5e-8
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ )

.model nch_ss_26 nmos (
+ level = 54
+ poxedge = 1
+ capmod = 2
+ wku0we = 2e-11
+ binunit = 2
+ mobmod = 0
+ pkvth0we = -1.3e-19
+ tvoff = 0.0019388906
+ vfbsdoff = 0.02
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ laigsd = -2.019482e-16
+ paramchk = 1
+ ku0we = -0.0007
+ beta0 = 13
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ leta0 = 0
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ ijthdfwd = 0.01
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ keta = -0.091670067
+ dmcgt = 0
+ tcjsw = 0.000357
+ lags = -1.7808411e-7
+ njtsswg = 9
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ ijthdrev = 0.01
+ lcit = 6.7178289e-10
+ kt1l = 0
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ lpdiblc2 = 2.6261368e-8
+ bigsd = 0.00125
+ ckappad = 0.6
+ ckappas = 0.6
+ lint = 6.5375218e-9
+ pdiblc1 = 0
+ pdiblc2 = 0.0017817666
+ toxref = 3e-9
+ pdiblcb = -0.3
+ lkt1 = 9.0572759e-9
+ lkt2 = -2.1662043e-8
+ lmax = 8.99743e-6
+ wvoff = 1.395365e-8
+ lmin = 8.974099999999999e-7
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ wvsat = -0.0028059037
+ wvth0 = -1.5516317e-8
+ minv = -0.3
+ wtvfbsdoff = 0
+ lua1 = -8.9279603e-16
+ lub1 = 6.8544226e-25
+ luc1 = -5.9256432e-18
+ waigc = 2.989874e-11
+ bigbacc = 0.002588
+ ndep = 1e+18
+ lkvth0we = -2e-12
+ lwlc = 0
+ moin = 5.1
+ ltvoff = -1.582327e-9
+ ltvfbsdoff = 0
+ lketa = 6.5795695e-8
+ kvth0we = 0.00018
+ nigc = 3.083
+ xpart = 1
+ lintnoi = -1.5e-8
+ acnqsmod = 0
+ pvfbsdoff = 0
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ egidl = 0.29734
+ vtsswgs = 4.2
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ lku0we = 2.5e-11
+ rbodymod = 0
+ epsrox = 3.9
+ pags = 1.7531187e-13
+ ntox = -0.31099999999999994
+ pcit = -1.0698337e-16
+ pclm = 1.5094578
+ rdsmod = 0
+ ptvfbsdoff = 0
+ igbmod = 1
+ phin = 0.15
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ pbswgd = 0.95
+ pkt1 = -2.7377875e-14
+ pkt2 = -4.4253241e-16
+ pbswgs = 0.95
+ igcmod = 1
+ wpdiblc2 = 5.7318301e-9
+ pvoff = -2.4799793e-15
+ cdscb = 0
+ cdscd = 0
+ rbdb = 50
+ pua1 = 1.9942546e-22
+ prwb = 0
+ prwg = 0
+ pub1 = -1.9939615e-31
+ puc1 = 1.7835157e-23
+ nfactor = 1
+ pvsat = 0
+ rbpb = 50
+ rbpd = 50
+ wk2we = 5e-12
+ rbps = 50
+ pvth0 = 3.3576501999999996e-15
+ rbsb = 50
+ pvag = 1.2
+ drout = 0.56
+ rdsw = 100
+ paigc = -1.0556924e-17
+ voffl = 0
+ paigsd = 1.1026372e-22
+ weta0 = -1.1162667e-8
+ wetab = 2.2325333e-8
+ wkvth0we = 2e-12
+ nigbacc = 10
+ permod = 1
+ trnqsmod = 0
+ cgidl = 0.22
+ rshg = 15.6
+ nigbinv = 10
+ pbswd = 0.8
+ pbsws = 0.8
+ voffcv = -0.16942
+ wpemod = 1
+ rgatemod = 0
+ tnjtsswg = 1
+ tnom = 25
+ pdits = 0
+ toxe = 2.47e-9
+ toxm = 2.43e-9
+ a0 = 3.8452644
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ cigsd = 0.069865
+ b1 = 0
+ at = -81312.781
+ cf = 7.5795e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.023723392000000003
+ k3 = -1.8419
+ em = 1000000.0
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ ll = 0
+ lw = 0
+ u0 = 0.01832456
+ w0 = 0
+ fnoimod = 1
+ ua = -1.6436128e-9
+ ub = 2.0158412e-18
+ uc = 5.8736458e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 5.6700000000000005e-9
+ ww = 0
+ xw = 3.4e-9
+ eigbinv = 1.1
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ tpbswg = 0.0009
+ wags = -7.4969804e-8
+ wcit = 3.0826906e-10
+ tnoia = 0
+ voff = -0.13348839
+ peta0 = 0
+ acde = 0.4
+ wketa = 1.8850903e-8
+ vsat = 102889.02
+ ptvoff = 2.7553621e-16
+ wint = 0
+ tpbsw = 0.0019
+ vth0 = 0.38649778
+ cigbacc = 0.32875
+ waigsd = 3.1111904e-12
+ wkt1 = 4.1483105e-9
+ wkt2 = -5.2803902e-9
+ cjswd = 8.774000000000001e-11
+ cjsws = 8.774000000000001e-11
+ wmax = 5.426e-7
+ mjswd = 0.11
+ aigc = 0.011795195
+ mjsws = 0.11
+ wmin = 2.726e-7
+ agidl = 9.41e-8
+ diomod = 1
+ tnoimod = 0
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 3.0174000000000004e-10
+ pku0we = -1.5e-18
+ wua1 = -2.0961923e-16
+ wub1 = 1.3682244e-25
+ cjswgs = 3.0174000000000004e-10
+ wuc1 = -2.9511024e-17
+ cigbinv = 0.006
+ bigc = 0.001442
+ wwlc = 0
+ tvfbsdoff = 0.022
+ cdsc = 0
+ mjswgd = 0.85
+ mjswgs = 0.85
+ scref = 1e-6
+ version = 4.5
+ ijthsfwd = 0.01
+ cgbo = 0
+ cgdl = 3.0874977e-12
+ cgdo = 4.5622265999999996e-11
+ xtid = 3
+ xtis = 3
+ pigcd = 2.621
+ cgsl = 3.0874977e-12
+ tcjswg = 0.001
+ cgso = 4.5622265999999996e-11
+ tempmod = 0
+ aigsd = 0.010772818
+ cigc = 0.000625
+ ags = 1.0774158
+ lvoff = -1.1649525e-8
+ cjd = 0.00145199
+ cit = 0.00026829437
+ cjs = 0.00145199
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ aigbacc = 0.02
+ dlc = 9.8024918e-9
+ lvsat = 0.0003
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ lvth0 = 5.1308999e-8
+ ijthsrev = 0.01
+ delta = 0.007595625
+ laigc = -1.416882e-10
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ la0 = -2.722152e-6
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ rnoia = 0
+ rnoib = 0
+ dmdg = 0
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = 0.20239035000000002
+ kt1 = -0.22156452
+ lk2 = -1.3986155e-8
+ kt2 = -0.033027229
+ llc = 0
+ lln = 1
+ lu0 = -2.2845026e-9
+ mjd = 0.26
+ aigbinv = 0.0163
+ lua = -2.9346741e-16
+ mjs = 0.26
+ lub = 5.7165214e-26
+ luc = 2.4824263e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 3.4236885e-13
+ fprout = 300
+ nsd = 1e+20
+ pbd = 0.52
+ pat = -6.3628324e-8
+ pbs = 0.52
+ pketa = -2.2733801e-14
+ pk2 = -1.3939214e-15
+ ngate = 8e+20
+ pu0 = 1.6539558e-16
+ xrcrg1 = 12
+ xrcrg2 = 1
+ k2we = 5e-5
+ prt = 0
+ pua = 4.226297e-23
+ pub = -4.4156209e-32
+ puc = -1.0695581e-23
+ pud = 0
+ ngcon = 1
+ wpclm = 9.3989653e-8
+ dsub = 0.75
+ rsh = 17.5
+ tcj = 0.00076
+ dtox = 2.7e-10
+ ua1 = 1.720591e-9
+ ub1 = -9.5473708e-19
+ uc1 = 7.0015137e-11
+ ppdiblc2 = -6.6555967e-15
+ tpb = 0.0014
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ wa0 = -4.9804098e-8
+ gbmin = 1e-12
+ ute = -1
+ wat = 0.078525419
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 2.0146831e-9
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ wtvoff = -3.0649189e-11
+ wlc = 0
+ wln = 1
+ wu0 = -1.2821044000000001e-9
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -1.3568102e-16
+ wub = 1.003525e-25
+ wuc = -1.2660669e-18
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ eta0 = 0.24044444
+ etab = -0.28088889
+ )

.model nch_ss_27 nmos (
+ level = 54
+ ntox = -0.31099999999999994
+ pcit = -1.1605802e-16
+ pclm = 1.5094578
+ fnoimod = 1
+ phin = 0.15
+ eigbinv = 1.1
+ pbswd = 0.8
+ pbsws = 0.8
+ pkt1 = 4.8128443e-15
+ pkt2 = 2.2738921e-15
+ pdits = 0
+ rbdb = 50
+ pua1 = -2.6369043e-23
+ prwb = 0
+ prwg = 0
+ pub1 = 4.8759292e-32
+ cigsd = 0.069865
+ puc1 = 6.8677984e-24
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ dvt0w = 0
+ pvag = 1.2
+ dvt1w = 0
+ dvt2w = 0
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ rdsw = 100
+ ijthsfwd = 0.01
+ cigbacc = 0.32875
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ tnoimod = 0
+ tnoia = 0
+ ijthsrev = 0.01
+ cigbinv = 0.006
+ peta0 = 0
+ rshg = 15.6
+ wketa = -2.2122195e-8
+ wtvfbsdoff = 0
+ tpbsw = 0.0019
+ toxref = 3e-9
+ cjswd = 8.774000000000001e-11
+ cjsws = 8.774000000000001e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ version = 4.5
+ ltvfbsdoff = 0
+ tempmod = 0
+ ppdiblc2 = 1.7501102e-15
+ tnom = 25
+ aigbacc = 0.02
+ tvfbsdoff = 0.022
+ toxe = 2.47e-9
+ toxm = 2.43e-9
+ ltvoff = 1.3913801e-9
+ ags = 0.40766657
+ scref = 1e-6
+ cjd = 0.00145199
+ cit = 0.00059502911
+ cjs = 0.00145199
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 9.8024918e-9
+ pigcd = 2.621
+ k3b = 1.9326
+ aigsd = 0.010772818
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ ptvfbsdoff = 0
+ aigbinv = 0.0163
+ lvoff = -5.0132203e-10
+ wags = 3.9484036e-7
+ lku0we = 2.5e-11
+ pkvth0we = -1.3e-19
+ la0 = 3.6355951e-7
+ epsrox = 3.9
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.052338453
+ kt1 = -0.19312528
+ lk2 = -1.4722356e-8
+ kt2 = -0.039065148
+ wcit = 3.184653e-10
+ lvsat = 0.0003
+ llc = 0
+ lln = 1
+ lu0 = -1.7576993e-9
+ mjd = 0.26
+ lvth0 = -8.2158156e-9
+ lua = -1.1159069e-16
+ mjs = 0.26
+ lub = -2.3732546e-26
+ luc = -2.9405776e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ voff = -0.14601446
+ njs = 1.02
+ pa0 = -3.8856002e-13
+ nsd = 1e+20
+ delta = 0.007595625
+ acde = 0.4
+ pbd = 0.52
+ wvfbsdoff = 0
+ pat = -7.9362363e-10
+ pbs = 0.52
+ rdsmod = 0
+ pk2 = 1.1847359e-15
+ lvfbsdoff = 0
+ laigc = -3.3762752e-11
+ pu0 = 1.2968191e-16
+ vfbsdoff = 0.02
+ igbmod = 1
+ prt = 0
+ pua = 2.9945529e-23
+ pub = -3.9782718e-32
+ puc = 6.3626704e-24
+ pud = 0
+ vsat = 102889.02
+ wint = 0
+ rnoia = 0
+ rnoib = 0
+ vth0 = 0.45337959
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 6.6639379e-10
+ ub1 = 1.1665789e-19
+ uc1 = 5.9635906e-11
+ wkt1 = -3.2021037e-8
+ wkt2 = -8.3325526e-9
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ tpb = 0.0014
+ wmax = 5.426e-7
+ wa0 = 7.714643e-7
+ aigc = 0.01167393
+ wmin = 2.726e-7
+ ute = -1
+ wat = 0.0079246317
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -8.8268726e-10
+ pbswgd = 0.95
+ pketa = 1.3732256e-14
+ poxedge = 1
+ pbswgs = 0.95
+ ngate = 8e+20
+ wlc = 0
+ wln = 1
+ wu0 = -1.2419767e-9
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -1.218412e-16
+ wub = 9.5438468e-26
+ wuc = -2.0432641e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ ngcon = 1
+ paramchk = 1
+ wpclm = 9.3989653e-8
+ igcmod = 1
+ binunit = 2
+ wua1 = 4.4082452e-17
+ wub1 = -1.420039e-25
+ wuc1 = -1.718815e-17
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ bigc = 0.001442
+ wwlc = 0
+ cdsc = 0
+ ijthdfwd = 0.01
+ cgbo = 0
+ cgdl = 3.0874977e-12
+ cgdo = 4.5622265999999996e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.0874977e-12
+ cgso = 4.5622265999999996e-11
+ cigc = 0.000625
+ permod = 1
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ ijthdrev = 0.01
+ tvoff = -0.0014023534
+ lpdiblc2 = -7.3119259e-9
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ voffcv = -0.16942
+ wpemod = 1
+ k2we = 5e-5
+ ku0we = -0.0007
+ dsub = 0.75
+ dtox = 2.7e-10
+ beta0 = 13
+ leta0 = 0
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ njtsswg = 9
+ lkvth0we = -2e-12
+ eta0 = 0.24044444
+ etab = -0.28088889
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.039504569
+ pdiblcb = -0.3
+ tpbswg = 0.0009
+ acnqsmod = 0
+ dmcgt = 0
+ tcjsw = 0.000357
+ rbodymod = 0
+ ptvoff = -5.8159511e-16
+ bigbacc = 0.002588
+ waigsd = 3.1113143e-12
+ bigsd = 0.00125
+ a0 = 0.37817284
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 204899.36
+ cf = 7.5795e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.024550589999999997
+ k3 = -1.8419
+ em = 1000000.0
+ kvth0we = 0.00018
+ diomod = 1
+ ll = 0
+ lw = 0
+ u0 = 0.017732646
+ w0 = 0
+ wvoff = 1.6411259e-8
+ ua = -1.8479686e-9
+ ub = 2.1067376e-18
+ uc = 1.1966909e-10
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 5.6700000000000005e-9
+ ww = 0
+ xw = 3.4e-9
+ lintnoi = -1.5e-8
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 3.0174000000000004e-10
+ pku0we = -1.5e-18
+ cjswgs = 3.0174000000000004e-10
+ bigbinv = 0.004953
+ wvsat = -0.0028059037
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ wvth0 = -1.8699761e-8
+ wpdiblc2 = -3.7127843e-9
+ waigc = 2.313153e-11
+ mjswgd = 0.85
+ mjswgs = 0.85
+ lketa = -4.8021757e-8
+ tcjswg = 0.001
+ xpart = 1
+ pvfbsdoff = 0
+ keta = 0.03621471
+ egidl = 0.29734
+ wkvth0we = 2e-12
+ lags = 4.1799271e-7
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 3.8098897e-10
+ trnqsmod = 0
+ kt1l = 0
+ nfactor = 1
+ lint = 6.5375218e-9
+ fprout = 300
+ lkt1 = -1.6253643e-8
+ lkt2 = -1.6288295e-8
+ xrcrg1 = 12
+ xrcrg2 = 1
+ lmax = 8.974099999999999e-7
+ lmin = 4.4741e-7
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ rgatemod = 0
+ wtvoff = 9.3241971e-10
+ pvoff = -4.6672513e-15
+ minv = -0.3
+ tnjtsswg = 1
+ lua1 = 4.5439491e-17
+ lub1 = -2.6809927e-25
+ luc1 = 3.3118724e-18
+ cdscb = 0
+ cdscd = 0
+ nigbacc = 10
+ ndep = 1e+18
+ pvsat = 0
+ wk2we = 5e-12
+ pvth0 = 6.1909158e-15
+ lwlc = 0
+ drout = 0.56
+ moin = 5.1
+ capmod = 2
+ paigc = -4.5341069e-18
+ nigc = 3.083
+ voffl = 0
+ wku0we = 2e-11
+ nigbinv = 10
+ mobmod = 0
+ weta0 = -1.1162667e-8
+ wetab = 2.2325333e-8
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ pags = -2.4281917e-13
+ cgidl = 0.22
+ )

.model nch_ss_28 nmos (
+ level = 54
+ wuc1 = -1.3268706e-17
+ bigc = 0.001442
+ ppclm = -7.9196439e-14
+ wwlc = 0
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ cdsc = 0
+ bigbacc = 0.002588
+ cgbo = 0
+ cgdl = 3.0874977e-12
+ cgdo = 4.5622265999999996e-11
+ xtid = 3
+ xtis = 3
+ wtvfbsdoff = 0
+ cgsl = 3.0874977e-12
+ cgso = 4.5622265999999996e-11
+ cigc = 0.000625
+ kvth0we = 0.00018
+ dmcgt = 0
+ tcjsw = 0.000357
+ wkvth0we = 2e-12
+ lintnoi = -1.5e-8
+ ltvfbsdoff = 0
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ trnqsmod = 0
+ toxref = 3e-9
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ bigsd = 0.00125
+ wvoff = 5.1767953e-9
+ k2we = 5e-5
+ dsub = 0.75
+ wvsat = -0.0054199005
+ dtox = 2.7e-10
+ ptvfbsdoff = 0
+ wvth0 = -1.0869543e-9
+ rgatemod = 0
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ tnjtsswg = 1
+ waigc = -1.6608588e-12
+ ltvoff = -7.6859018e-11
+ eta0 = 0.24044444
+ etab = -0.28088889
+ lketa = -5.7215427e-9
+ nfactor = 1
+ xpart = 1
+ pvfbsdoff = 0
+ lku0we = 2.5e-11
+ egidl = 0.29734
+ epsrox = 3.9
+ rdsmod = 0
+ igbmod = 1
+ nigbacc = 10
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ pbswgd = 0.95
+ pbswgs = 0.95
+ igcmod = 1
+ nigbinv = 10
+ pvoff = 2.7591262e-16
+ cdscb = 0
+ cdscd = 0
+ pvsat = 1.1501586e-9
+ wk2we = 5e-12
+ pvth0 = -1.5587192000000002e-15
+ drout = 0.56
+ paigc = 6.374544e-18
+ ijthsfwd = 0.01
+ paigsd = 2.2627557e-23
+ voffl = 0
+ fnoimod = 1
+ eigbinv = 1.1
+ keta = -0.05992214
+ weta0 = -1.1162667e-8
+ wetab = 2.2325333e-8
+ permod = 1
+ lpclm = 1.4504842e-7
+ lags = 5.906061e-7
+ jswd = 1.28e-13
+ ijthsrev = 0.01
+ jsws = 1.28e-13
+ lcit = 9.7365571e-11
+ cgidl = 0.22
+ kt1l = 0
+ lint = 9.7879675e-9
+ voffcv = -0.16942
+ wpemod = 1
+ lkt1 = 8.8603069e-9
+ lkt2 = -2.5638367e-9
+ lmax = 4.4741e-7
+ cigbacc = 0.32875
+ pbswd = 0.8
+ pbsws = 0.8
+ lmin = 2.1410000000000002e-7
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ ppdiblc2 = -5.242001e-17
+ tnoimod = 0
+ minv = -0.3
+ lua1 = -4.6794128e-17
+ lub1 = -3.2889654e-26
+ luc1 = -2.1335001e-17
+ pdits = 0
+ ndep = 1e+18
+ cigsd = 0.069865
+ cigbinv = 0.006
+ dvt0w = 0
+ lwlc = 0
+ dvt1w = 0
+ dvt2w = 0
+ moin = 5.1
+ nigc = 3.083
+ tpbswg = 0.0009
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ version = 4.5
+ tempmod = 0
+ pkvth0we = -1.3e-19
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ tnoia = 0
+ pags = 1.2428184e-13
+ peta0 = 0
+ ptvoff = -1.5558646e-16
+ aigbacc = 0.02
+ ntox = -0.31099999999999994
+ pcit = -8.9847229e-18
+ pclm = 1.1798023
+ waigsd = 3.1112628e-12
+ wketa = 2.3981389e-8
+ vfbsdoff = 0.02
+ tpbsw = 0.0019
+ cjswd = 8.774000000000001e-11
+ cjsws = 8.774000000000001e-11
+ diomod = 1
+ mjswd = 0.11
+ phin = 0.15
+ mjsws = 0.11
+ agidl = 9.41e-8
+ pditsd = 0
+ pditsl = 0
+ aigbinv = 0.0163
+ pkt1 = -1.2500052e-14
+ pkt2 = -7.0784646e-16
+ cjswgd = 3.0174000000000004e-10
+ pku0we = -1.5e-18
+ cjswgs = 3.0174000000000004e-10
+ paramchk = 1
+ ags = 0.015363416000000005
+ cjd = 0.00145199
+ tvfbsdoff = 0.022
+ cit = 0.0012396277
+ cjs = 0.00145199
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 1.30529375e-8
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ rbdb = 50
+ pua1 = 1.8291934e-23
+ prwb = 0
+ prwg = 0
+ pub1 = -6.5524188e-33
+ puc1 = 5.143243e-24
+ mjswgd = 0.85
+ mjswgs = 0.85
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ tcjswg = 0.001
+ rdsw = 100
+ scref = 1e-6
+ ijthdfwd = 0.01
+ la0 = -6.0902319e-7
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.014636938
+ kt1 = -0.25020244
+ lk2 = -1.0681005e-8
+ kt2 = -0.070257098
+ pigcd = 2.621
+ llc = -1.18e-13
+ lln = 0.7
+ aigsd = 0.010772818
+ lu0 = -7.1183626e-10
+ mjd = 0.26
+ lua = -1.8564943e-17
+ mjs = 0.26
+ lub = -5.2748233e-26
+ luc = -4.2757753e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 2.2627554e-14
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 2.6237001000000004e-9
+ poxedge = 1
+ pbs = 0.52
+ pk2 = 8.6250113e-16
+ lvoff = -7.1474494e-9
+ a0 = 2.5885881
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ pu0 = 5.1138272e-17
+ at = 119214.09
+ cf = 7.5795e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.015365692
+ k3 = -1.8419
+ em = 1000000.0
+ prt = 0
+ pua = 5.6394132e-24
+ pub = -7.710339e-34
+ puc = -1.5613012e-24
+ pud = 0
+ ll = -1.18e-13
+ lw = 0
+ u0 = 0.015355684
+ w0 = 0
+ ua = -2.0593908e-9
+ ub = 2.1726824e-18
+ uc = 6.2555449e-11
+ ud = 0
+ wl = 0
+ rsh = 17.5
+ wr = 1
+ xj = 8.6e-8
+ xl = 5.6700000000000005e-9
+ ww = 0
+ xw = 3.4e-9
+ tcj = 0.00076
+ ua1 = 8.7601565e-10
+ lvsat = -0.0038672412000000005
+ ub1 = -4.1790941e-19
+ uc1 = 1.1565153e-10
+ binunit = 2
+ lvth0 = 1.474398e-9
+ ijthdrev = 0.01
+ tpb = 0.0014
+ wvfbsdoff = 0
+ wa0 = -1.6305293e-7
+ lvfbsdoff = 0
+ ute = -1
+ wat = 0.00015798693
+ delta = 0.007595625
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -1.5033038e-10
+ laigc = -3.7429738e-11
+ wlc = 0
+ wln = 1
+ rshg = 15.6
+ wu0 = -1.0634684000000002e-9
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -6.6600022e-17
+ wub = 6.7755498e-27
+ wuc = -2.4236148e-18
+ wud = 0
+ lpdiblc2 = -4.2799755e-9
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ rnoia = 0
+ rnoib = 0
+ fprout = 300
+ xrcrg1 = 12
+ xrcrg2 = 1
+ pketa = -6.5533207e-15
+ ngate = 8e+20
+ ngcon = 1
+ wpclm = 2.7398156e-7
+ wtvoff = -3.5781771e-11
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ tnom = 25
+ jswgs = 1.28e-13
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ toxe = 2.47e-9
+ toxm = 2.43e-9
+ lkvth0we = -2e-12
+ capmod = 2
+ wku0we = 2e-11
+ mobmod = 0
+ acnqsmod = 0
+ wags = -4.3948013e-7
+ wcit = 7.5116891e-11
+ rbodymod = 0
+ voff = -0.13090963
+ acde = 0.4
+ tvoff = 0.0019345538
+ njtsswg = 9
+ vsat = 112360.02
+ wint = 0
+ xjbvd = 1
+ xjbvs = 1
+ vth0 = 0.43135638000000004
+ lk2we = -1.5e-12
+ wkt1 = 7.3264548e-9
+ wkt2 = -1.5558741e-9
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ wmax = 5.426e-7
+ laigsd = -8.1983894e-17
+ aigc = 0.011682264
+ wmin = 2.726e-7
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.032613772
+ pdiblcb = -0.3
+ ku0we = -0.0007
+ beta0 = 13
+ leta0 = 0
+ wua1 = -5.7419768e-17
+ wpdiblc2 = 3.8387521e-10
+ wub1 = -1.6295463e-26
+ )

.model nch_ss_29 nmos (
+ level = 54
+ keta = 0.0092481698
+ aigbinv = 0.0163
+ tnoia = 0
+ ijthdrev = 0.01
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = -9.537106e-12
+ peta0 = 0
+ ptvfbsdoff = 0
+ kt1l = 0
+ wketa = -2.0169501e-8
+ toxref = 3e-9
+ lpdiblc2 = -9.0824285e-10
+ tpbsw = 0.0019
+ ags = 2.8144443999999997
+ cjswd = 8.774000000000001e-11
+ cjsws = 8.774000000000001e-11
+ lint = 9.7879675e-9
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ cjd = 0.00145199
+ cit = 0.0017462755
+ cjs = 0.00145199
+ clc = 1e-7
+ cle = 0.6
+ lkt1 = -2.5262126e-9
+ bvd = 8.7
+ lkt2 = -3.9513595e-9
+ bvs = 8.7
+ lmax = 2.1410000000000002e-7
+ dlc = 1.30529375e-8
+ lmin = 8.833e-8
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ poxedge = 1
+ tvfbsdoff = 0.022
+ la0 = -2.075695e-7
+ minv = -0.3
+ jsd = 6.11e-7
+ ltvoff = 5.8839234e-11
+ jss = 6.11e-7
+ lat = -0.0011937311
+ lua1 = -5.8912951e-18
+ lub1 = -2.9377439e-26
+ luc1 = 1.0640856e-17
+ kt1 = -0.1962379
+ lk2 = -3.2022951e-9
+ kt2 = -0.063681161
+ llc = -1.18e-13
+ binunit = 2
+ lln = 0.7
+ lu0 = -2.6151767e-10
+ mjd = 0.26
+ lua = 5.2959027e-17
+ mjs = 0.26
+ lub = -7.97606935e-26
+ luc = -8.8267893e-18
+ lud = 0
+ lwc = 0
+ ndep = 1e+18
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ lkvth0we = -2e-12
+ njs = 1.02
+ pa0 = 1.0407708e-13
+ nsd = 1e+20
+ lwlc = 0
+ pbd = 0.52
+ pat = -3.1161951e-10
+ pbs = 0.52
+ pk2 = -9.7578421e-17
+ moin = 5.1
+ pu0 = 1.8260797e-17
+ prt = 0
+ pua = -7.1102082e-24
+ pub = 9.57267e-33
+ puc = 7.19078e-25
+ pud = 0
+ scref = 1e-6
+ nigc = 3.083
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 6.8216336e-10
+ pigcd = 2.621
+ ub1 = -4.3455498e-19
+ uc1 = -3.5892821e-11
+ aigsd = 0.010772818
+ tpb = 0.0014
+ lku0we = 2.5e-11
+ wa0 = -5.4906963e-7
+ acnqsmod = 0
+ ute = -1
+ wat = 0.014069454
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 4.3998097e-9
+ epsrox = 3.9
+ lvoff = 2.33236653e-9
+ wlc = 0
+ wln = 1
+ wu0 = -9.076509899999999e-10
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -6.1752756e-18
+ wub = -4.2246744000000004e-26
+ wuc = -1.3231099e-17
+ wud = 0
+ wwc = 0
+ noff = 2.7195
+ wwl = 0
+ wwn = 1
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ lvsat = -0.00015734827000000009
+ rbodymod = 0
+ rdsmod = 0
+ wvfbsdoff = 0
+ lvth0 = -1.2194990599999998e-8
+ lvfbsdoff = 0
+ igbmod = 1
+ delta = 0.007595625
+ laigc = 2.6175146e-12
+ ntox = -0.31099999999999994
+ pcit = 7.8208248e-18
+ jtsswgd = 2.3e-7
+ pclm = 2.3689724
+ jtsswgs = 2.3e-7
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ rnoia = 0
+ rnoib = 0
+ pbswgd = 0.95
+ pbswgs = 0.95
+ phin = 0.15
+ pketa = 2.762517e-15
+ ngate = 8e+20
+ igcmod = 1
+ ngcon = 1
+ pkt1 = 6.6516645e-16
+ pkt2 = 9.3582987e-16
+ wpclm = -2.0834879e-7
+ wpdiblc2 = 1.3111248e-10
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ rbdb = 50
+ pua1 = 1.9734917e-24
+ prwb = 0
+ prwg = 0
+ pub1 = -5.2222001e-33
+ puc1 = -4.0873907e-24
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ njtsswg = 9
+ paigsd = -9.4615512e-24
+ rdsw = 100
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ permod = 1
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.016633997
+ pdiblcb = -0.3
+ wkvth0we = 2e-12
+ trnqsmod = 0
+ tvoff = 0.0012914341
+ rshg = 15.6
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ voffcv = -0.16942
+ wpemod = 1
+ bigbacc = 0.002588
+ ku0we = -0.0007
+ kvth0we = 0.00018
+ beta0 = 13
+ leta0 = 0
+ rgatemod = 0
+ lintnoi = -1.5e-8
+ tnjtsswg = 1
+ tnom = 25
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ ppclm = 2.2575265e-14
+ vtsswgs = 4.2
+ toxe = 2.47e-9
+ toxm = 2.43e-9
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ tpbswg = 0.0009
+ dmcgt = 0
+ wags = 1.4953333e-7
+ tcjsw = 0.000357
+ wcit = -4.5302538e-12
+ ptvoff = 2.7225835e-17
+ voff = -0.175837897
+ waigsd = 3.1114149e-12
+ acde = 0.4
+ vsat = 94777.65030000001
+ wint = 0
+ bigsd = 0.00125
+ vth0 = 0.49614045399999995
+ diomod = 1
+ wkt1 = -5.5067946e-8
+ wkt2 = -9.3458092e-9
+ wmax = 5.426e-7
+ aigc = 0.011492467
+ wmin = 2.726e-7
+ nfactor = 1
+ pditsd = 0
+ pditsl = 0
+ wvoff = 8.989216699999998e-9
+ cjswgd = 3.0174000000000004e-10
+ pku0we = -1.5e-18
+ cjswgs = 3.0174000000000004e-10
+ wvsat = -0.0005775380999999999
+ wvth0 = -1.4525727999999998e-8
+ wua1 = 1.991882e-17
+ wub1 = -2.2599817e-26
+ wuc1 = 3.0478373e-17
+ waigc = 3.9031408e-11
+ bigc = 0.001442
+ mjswgd = 0.85
+ mjswgs = 0.85
+ wwlc = 0
+ tcjswg = 0.001
+ nigbacc = 10
+ lketa = -2.0316478e-8
+ cdsc = 0
+ ijthsfwd = 0.01
+ cgbo = 0
+ xpart = 1
+ cgdl = 3.0874977e-12
+ cgdo = 4.5622265999999996e-11
+ pvfbsdoff = 0
+ xtid = 3
+ xtis = 3
+ cgsl = 3.0874977e-12
+ cgso = 4.5622265999999996e-11
+ cigc = 0.000625
+ egidl = 0.29734
+ nigbinv = 10
+ ijthsrev = 0.01
+ fprout = 300
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ fnoimod = 1
+ k2we = 5e-5
+ wtvoff = -9.0219076e-10
+ eigbinv = 1.1
+ dsub = 0.75
+ dtox = 2.7e-10
+ ppdiblc2 = 9.1292629e-19
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ pvoff = -5.285090499999998e-16
+ a0 = 0.68596391
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 55502.213
+ cf = 7.5795e-11
+ cdscb = 0
+ cdscd = 0
+ ef = 1.0
+ k1 = 0.274
+ k2 = -0.02007843
+ k3 = -1.8419
+ em = 1000000.0
+ ll = -1.18e-13
+ lw = 0
+ u0 = 0.013221473
+ pvsat = 1.2842156000000008e-10
+ w0 = 0
+ ua = -2.398367e-9
+ ub = 2.300703286e-18
+ uc = 8.4124236e-11
+ ud = 0
+ wk2we = 5e-12
+ capmod = 2
+ wl = 0
+ wr = 1
+ pvth0 = 1.276862e-15
+ xj = 8.6e-8
+ xl = 5.6700000000000005e-9
+ ww = 0
+ eta0 = 0.24044444
+ xw = 3.4e-9
+ drout = 0.56
+ etab = -0.28088889
+ wku0we = 2e-11
+ paigc = -2.2115244e-18
+ mobmod = 0
+ voffl = 0
+ cigbacc = 0.32875
+ weta0 = -1.1162667e-8
+ wetab = 2.2325333e-8
+ pkvth0we = -1.3e-19
+ lpclm = -1.0586647e-7
+ tnoimod = 0
+ cgidl = 0.22
+ vfbsdoff = 0.02
+ cigbinv = 0.006
+ laigsd = 3.4280989e-17
+ pbswd = 0.8
+ pbsws = 0.8
+ paramchk = 1
+ version = 4.5
+ wtvfbsdoff = 0
+ tempmod = 0
+ pdits = 0
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ cigsd = 0.069865
+ ltvfbsdoff = 0
+ dvt0w = 0
+ aigbacc = 0.02
+ dvt1w = 0
+ dvt2w = 0
+ ijthdfwd = 0.01
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ )

.model nch_ss_30 nmos (
+ level = 54
+ keta = -0.29566775
+ aigbinv = 0.0163
+ tnoia = 0
+ ijthdrev = 0.01
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 2.6988428000000004e-10
+ peta0 = -9.3037135e-16
+ ptvfbsdoff = 0
+ petab = -1.2138265e-15
+ kt1l = 0
+ wketa = -4.7865407e-8
+ toxref = 3e-9
+ lpdiblc2 = 8.2379047e-15
+ tpbsw = 0.0019
+ ags = 2.8144443999999997
+ cjswd = 8.774000000000001e-11
+ cjsws = 8.774000000000001e-11
+ lint = 0
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ cjd = 0.00145199
+ cit = -0.0012262896700000001
+ cjs = 0.00145199
+ clc = 1e-7
+ cle = 0.6
+ lkt1 = -8.4950836e-9
+ bvd = 8.7
+ lkt2 = 3.8424987e-10
+ bvs = 8.7
+ lmax = 8.833e-8
+ dlc = 3.26497e-9
+ lmin = 5.233e-8
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ poxedge = 1
+ tvfbsdoff = 0.022
+ la0 = 3.9829889e-7
+ minv = -0.3
+ jsd = 6.11e-7
+ ltvoff = -2.7237524e-10
+ jss = 6.11e-7
+ lat = 0.00568560498
+ lua1 = -1.2736334e-17
+ lub1 = 1.6085594e-26
+ luc1 = -2.4540957899999996e-18
+ kt1 = -0.13273927
+ lk2 = 1.0502722e-9
+ kt2 = -0.10980467
+ llc = 0
+ binunit = 2
+ lln = 1
+ lu0 = -2.1075966000000001e-10
+ mjd = 0.26
+ lua = -7.6887484e-18
+ mjs = 0.26
+ lub = 6.3606825e-27
+ luc = -3.2720592999999998e-18
+ lud = 0
+ lwc = 0
+ ndep = 1e+18
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ lkvth0we = -2e-12
+ njs = 1.02
+ pa0 = -1.1411036e-13
+ nsd = 1e+20
+ lwlc = 0
+ pbd = 0.52
+ pat = -1.6720563e-9
+ pbs = 0.52
+ pk2 = -3.7289588e-16
+ moin = 5.1
+ pu0 = 7.2584501e-17
+ prt = 0
+ pua = 1.3044266e-23
+ pub = -1.13966382e-32
+ puc = 2.3653651e-24
+ pud = 0
+ scref = 1e-6
+ nigc = 3.083
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 7.5498293e-10
+ pigcd = 2.621
+ ub1 = -9.1820427e-19
+ uc1 = 1.03415541e-10
+ aigsd = 0.010772818
+ tpb = 0.0014
+ lku0we = 2.5e-11
+ wa0 = 1.7720733e-6
+ acnqsmod = 0
+ ute = -1
+ wat = 0.028542186400000003
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 7.3287188e-9
+ epsrox = 3.9
+ lvoff = -3.2511799e-9
+ wlc = 0
+ wln = 1
+ wu0 = -1.4855627e-9
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -2.2058458e-16
+ wub = 1.80830997e-25
+ wuc = -3.0744792e-17
+ wud = 0
+ wwc = 0
+ noff = 2.7195
+ wwl = 0
+ wwn = 1
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ lvsat = 0.0056945043
+ rbodymod = 0
+ rdsmod = 0
+ wvfbsdoff = 0
+ lvth0 = 3.589724300000001e-9
+ lvfbsdoff = 0
+ igbmod = 1
+ delta = 0.007595625
+ laigc = -3.0244582e-11
+ ntox = -0.31099999999999994
+ pcit = -3.6362976e-17
+ jtsswgd = 2.3e-7
+ pclm = 1.7776553
+ jtsswgs = 2.3e-7
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ rnoia = 0
+ rnoib = 0
+ pbswgd = 0.95
+ pbswgs = 0.95
+ phin = 0.15
+ pketa = 5.3659323e-15
+ ngate = 8e+20
+ igcmod = 1
+ ngcon = 1
+ pkt1 = 5.1065068e-15
+ pkt2 = -5.9202052e-16
+ wpclm = 4.3365813e-8
+ wpdiblc2 = 1.4083642e-10
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ rbdb = 50
+ pua1 = 4.1884121e-24
+ prwb = 0
+ prwg = 0
+ pub1 = -9.7869988e-33
+ puc1 = 3.1185952000000005e-24
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ njtsswg = 9
+ rdsw = 100
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ permod = 1
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.0069717513
+ pdiblcb = -0.3
+ wkvth0we = 2e-12
+ trnqsmod = 0
+ tvoff = 0.0048149924
+ rshg = 15.6
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ voffcv = -0.16942
+ wpemod = 1
+ bigbacc = 0.002588
+ ku0we = -0.0007
+ kvth0we = 0.00018
+ beta0 = 13
+ leta0 = 2.0040249e-8
+ rgatemod = 0
+ letab = -2.6551319e-8
+ lintnoi = -1.5e-8
+ tnjtsswg = 1
+ tnom = 25
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ ppclm = -1.085908e-15
+ vtsswgs = 4.2
+ toxe = 2.47e-9
+ toxm = 2.43e-9
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ tpbswg = 0.0009
+ dmcgt = 0
+ wags = 1.4953333e-7
+ tcjsw = 0.000357
+ wcit = 4.6550956e-10
+ ptvoff = 9.0058483e-17
+ voff = -0.116438471
+ waigsd = 3.1113143e-12
+ acde = 0.4
+ vsat = 32523.893000000004
+ wint = 0
+ bigsd = 0.00125
+ vth0 = 0.328217953
+ diomod = 1
+ wkt1 = -1.0231625000000001e-7
+ wkt2 = 6.9079183e-9
+ wmax = 5.426e-7
+ aigc = 0.011842064
+ wmin = 2.726e-7
+ nfactor = 1
+ pditsd = 0
+ pditsl = 0
+ wvoff = 4.307686799999997e-9
+ cjswgd = 3.0174000000000004e-10
+ pku0we = -1.5e-18
+ cjswgs = 3.0174000000000004e-10
+ wvsat = 0.0127657745
+ wvth0 = -4.1257771e-9
+ wua1 = -3.6441631e-18
+ wub1 = 2.5961869999999995e-26
+ wuc1 = -4.618107e-17
+ waigc = 4.5087747e-12
+ bigc = 0.001442
+ mjswgd = 0.85
+ mjswgs = 0.85
+ wwlc = 0
+ tcjswg = 0.001
+ nigbacc = 10
+ lketa = 8.345618e-9
+ cdsc = 0
+ ijthsfwd = 0.01
+ cgbo = 0
+ xpart = 1
+ cgdl = 3.0874977e-12
+ cgdo = 4.5622265999999996e-11
+ pvfbsdoff = 0
+ xtid = 3
+ xtis = 3
+ cgsl = 3.0874977e-12
+ cgso = 4.5622265999999996e-11
+ cigc = 0.000625
+ egidl = 0.29734
+ nigbinv = 10
+ ijthsrev = 0.01
+ fprout = 300
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ fnoimod = 1
+ k2we = 5e-5
+ wtvoff = -1.5706231e-9
+ eigbinv = 1.1
+ dsub = 0.75
+ dtox = 2.7e-10
+ ppdiblc2 = -1.1241984e-21
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ pvoff = -8.844511799999994e-17
+ a0 = -5.7594444
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = -17682.2125
+ cf = 7.5795e-11
+ cdscb = 0
+ cdscd = 0
+ ef = 1.0
+ k1 = 0.274
+ k2 = -0.065318509
+ k3 = -1.8419
+ em = 1000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.012681494
+ pvsat = -1.1258518e-9
+ w0 = 0
+ ua = -1.7531779e-9
+ ub = 1.3845184050000002e-18
+ uc = 2.5031363e-11
+ ud = 0
+ wk2we = 5e-12
+ capmod = 2
+ wl = 0
+ wr = 1
+ pvth0 = 2.9926666000000004e-16
+ xj = 8.6e-8
+ xl = 5.6700000000000005e-9
+ ww = 0
+ eta0 = 0.027250304
+ xw = 3.4e-9
+ drout = 0.56
+ etab = 0.001571952
+ wku0we = 2e-11
+ paigc = 1.0336032e-18
+ mobmod = 0
+ voffl = 0
+ cigbacc = 0.32875
+ weta0 = -1.2650991e-9
+ wetab = 3.5238381e-8
+ pkvth0we = -1.3e-19
+ lpclm = -5.0282662e-8
+ tnoimod = 0
+ cgidl = 0.22
+ vfbsdoff = 0.02
+ cigbinv = 0.006
+ pbswd = 0.8
+ pbsws = 0.8
+ paramchk = 1
+ version = 4.5
+ wtvfbsdoff = 0
+ tempmod = 0
+ pdits = 0
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ cigsd = 0.069865
+ ltvfbsdoff = 0
+ dvt0w = 0
+ aigbacc = 0.02
+ dvt1w = 0
+ dvt2w = 0
+ ijthdfwd = 0.01
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ )

.model nch_ss_31 nmos (
+ level = 54
+ nigbacc = 10
+ wvoff = 2.6164685300000083e-9
+ wvsat = 0.004955544200000002
+ wvth0 = -2.7687313000000006e-8
+ ltvoff = 2.6647905e-10
+ waigc = 1.8753243e-11
+ tnom = 25
+ nigbinv = 10
+ toxe = 2.47e-9
+ toxm = 2.43e-9
+ lketa = -2.3617222e-8
+ pvfbsdoff = 0
+ xpart = 1
+ lku0we = 2.5e-11
+ epsrox = 3.9
+ egidl = 0.29734
+ fnoimod = 1
+ pkvth0we = -1.3e-19
+ wags = 1.4953333e-7
+ rdsmod = 0
+ eigbinv = 1.1
+ wcit = 5.6353234e-10
+ igbmod = 1
+ voff = -0.07382279000000001
+ acde = 0.4
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ vfbsdoff = 0.02
+ vsat = 88577.58000000002
+ pbswgd = 0.95
+ pbswgs = 0.95
+ wint = 0
+ vth0 = 0.34762439000000006
+ wkt1 = -1.5494349e-8
+ wkt2 = -2.0876247e-8
+ wmax = 5.426e-7
+ igcmod = 1
+ aigc = 0.011696193
+ wmin = 2.726e-7
+ paramchk = 1
+ cigbacc = 0.32875
+ wua1 = -1.1132499e-16
+ wub1 = 7.746798000000004e-26
+ wuc1 = 2.2143851000000003e-16
+ pvoff = 9.645440000000495e-18
+ bigc = 0.001442
+ cdscb = 0
+ cdscd = 0
+ tnoimod = 0
+ wwlc = 0
+ pvsat = -6.72859e-10
+ wk2we = 5e-12
+ pvth0 = 1.6658357999999994e-15
+ drout = 0.56
+ paigsd = 1.7624612e-23
+ cdsc = 0
+ paigc = 2.0742404e-19
+ cigbinv = 0.006
+ ijthdfwd = 0.01
+ cgbo = 0
+ cgdl = 3.0874977e-12
+ cgdo = 4.5622265999999996e-11
+ xtid = 3
+ xtis = 3
+ voffl = 0
+ cgsl = 3.0874977e-12
+ cgso = 4.5622265999999996e-11
+ cigc = 0.000625
+ permod = 1
+ weta0 = -1.2005104e-7
+ wetab = 5.6750807e-8
+ lpclm = 5.458214e-8
+ version = 4.5
+ tempmod = 0
+ ijthdrev = 0.01
+ cgidl = 0.22
+ voffcv = -0.16942
+ wpemod = 1
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ aigbacc = 0.02
+ pbswd = 0.8
+ pbsws = 0.8
+ k2we = 5e-5
+ dsub = 0.75
+ dtox = 2.7e-10
+ aigbinv = 0.0163
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ pdits = 0
+ cigsd = 0.069865
+ lkvth0we = -2e-12
+ eta0 = 1.0176617
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ etab = -1.3959412
+ tpbswg = 0.0009
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ acnqsmod = 0
+ tnoia = 0
+ ptvoff = -4.401556e-18
+ poxedge = 1
+ rbodymod = 0
+ ags = 2.8144443999999997
+ waigsd = 3.1110104e-12
+ peta0 = 5.9592132e-15
+ cjd = 0.00145199
+ cit = -0.0058674639
+ cjs = 0.00145199
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ petab = -2.4615472e-15
+ dlc = 3.26497e-9
+ binunit = 2
+ wketa = -5.877032e-8
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ diomod = 1
+ tpbsw = 0.0019
+ cjswd = 8.774000000000001e-11
+ cjsws = 8.774000000000001e-11
+ mjswd = 0.11
+ pditsd = 0
+ pditsl = 0
+ mjsws = 0.11
+ agidl = 9.41e-8
+ cjswgd = 3.0174000000000004e-10
+ pku0we = -1.5e-18
+ cjswgs = 3.0174000000000004e-10
+ la0 = -1.4097724e-8
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.0003194376999999999
+ kt1 = -0.39757001
+ lk2 = 7.4338958e-10
+ kt2 = -0.14677127
+ llc = 0
+ lln = 1
+ lu0 = 5.7832928e-10
+ mjd = 0.26
+ lua = 6.4763643e-17
+ mjs = 0.26
+ lub = -2.3096342000000002e-26
+ luc = -1.0931136000000001e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = -1.7333804e-13
+ nsd = 1e+20
+ pbd = 0.52
+ pat = -3.7789471e-10
+ tvfbsdoff = 0.022
+ pbs = 0.52
+ pk2 = -1.0803308e-16
+ wpdiblc2 = 1.4081704e-10
+ pu0 = -6.727698299999999e-17
+ prt = 0
+ pua = -2.1774501e-24
+ pub = -5.473259300000002e-33
+ puc = 4.761497700000001e-24
+ pud = 0
+ mjswgd = 0.85
+ mjswgs = 0.85
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 1.4910078e-9
+ ub1 = -1.94643208e-18
+ uc1 = -6.027858599999999e-10
+ tpb = 0.0014
+ tcjswg = 0.001
+ wa0 = 2.7932403e-6
+ ute = -1
+ wat = 0.006229054600000004
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 2.7621189e-9
+ wlc = 0
+ wln = 1
+ wu0 = 9.258426e-10
+ jtsswgd = 2.3e-7
+ xgl = -1.09e-8
+ jtsswgs = 2.3e-7
+ xgw = 0
+ wua = 4.1858808e-17
+ wub = 7.870378029999999e-26
+ wuc = -7.2057435e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ scref = 1e-6
+ pigcd = 2.621
+ aigsd = 0.010772819
+ keta = 0.2554158
+ lvoff = -5.722889800000002e-9
+ wkvth0we = 2e-12
+ wvfbsdoff = 0
+ lvsat = 0.0024434015700000003
+ lvfbsdoff = 0
+ lvth0 = 2.4641506e-9
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 5.390715899999999e-10
+ trnqsmod = 0
+ delta = 0.007595625
+ laigc = -2.1784105e-11
+ kt1l = 0
+ fprout = 300
+ xrcrg1 = 12
+ xrcrg2 = 1
+ rnoia = 0
+ rnoib = 0
+ lint = 0
+ njtsswg = 9
+ lkt1 = 6.8650994e-9
+ lkt2 = 2.528313e-9
+ pketa = 5.998417e-15
+ ngate = 8e+20
+ lmax = 5.233e-8
+ lmin = 4.333e-8
+ wtvoff = 5.799816e-11
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ ngcon = 1
+ wpclm = 2.4669208e-7
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ ckappad = 0.6
+ ckappas = 0.6
+ rgatemod = 0
+ gbmin = 1e-12
+ pdiblc1 = 0
+ pdiblc2 = 0.0069718933
+ pdiblcb = -0.3
+ tnjtsswg = 1
+ minv = -0.3
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ lua1 = -5.5425775e-17
+ lub1 = 7.572278e-26
+ luc1 = 3.8505613e-17
+ capmod = 2
+ ndep = 1e+18
+ wku0we = 2e-11
+ lwlc = 0
+ moin = 5.1
+ mobmod = 0
+ nigc = 3.083
+ bigbacc = 0.002588
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ kvth0we = 0.00018
+ wtvfbsdoff = 0
+ lintnoi = -1.5e-8
+ bigbinv = 0.004953
+ tvoff = -0.0044755986
+ ntox = -0.31099999999999994
+ vtsswgd = 4.2
+ pcit = -4.2048497e-17
+ vtsswgs = 4.2
+ pclm = -0.030358553
+ laigsd = -6.385731e-17
+ xjbvd = 1
+ a0 = 1.350842
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ xjbvs = 1
+ lk2we = -1.5e-12
+ at = 85853.00300000001
+ cf = 7.5795e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = -0.060027428
+ k3 = -1.8419
+ em = 1000000.0
+ ltvfbsdoff = 0
+ ll = 0
+ lw = 0
+ u0 = -0.0009234929531000001
+ w0 = 0
+ ua = -3.002357e-9
+ ub = 1.89239813e-18
+ uc = 1.5708441000000004e-10
+ ud = 0
+ phin = 0.15
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 5.6700000000000005e-9
+ ww = 0
+ xw = 3.4e-9
+ pkt1 = 7.083666e-17
+ pkt2 = 1.019461e-15
+ ku0we = -0.0007
+ beta0 = 13
+ leta0 = -3.7403611e-8
+ letab = 5.4504443e-8
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ ppclm = -1.2878832e-14
+ rbdb = 50
+ pua1 = 1.04339e-23
+ prwb = 0
+ prwg = 0
+ pub1 = -1.27743519e-32
+ puc1 = -1.24033186e-23
+ rbpb = 50
+ rbpd = 50
+ dlcig = 2.5e-9
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ bgidl = 2320000000.0
+ ptvfbsdoff = 0
+ rdsw = 100
+ ijthsfwd = 0.01
+ nfactor = 1
+ dmcgt = 0
+ tcjsw = 0.000357
+ ijthsrev = 0.01
+ toxref = 3e-9
+ rshg = 15.6
+ bigsd = 0.00125
+ )

.model nch_ss_32 nmos (
+ level = 54
+ eta0 = -0.25440451
+ etab = -0.81370191
+ scref = 1e-6
+ lku0we = 2.5e-11
+ pigcd = 2.621
+ epsrox = 3.9
+ aigsd = 0.010772817
+ njtsswg = 9
+ lvoff = -7.2316898e-9
+ rdsmod = 0
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ igbmod = 1
+ lvsat = -0.0021690246
+ ckappad = 0.6
+ ckappas = 0.6
+ lvth0 = -6.79131000000006e-11
+ pdiblc1 = 0
+ pdiblc2 = 0.0069718933
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ pdiblcb = -0.3
+ delta = 0.007595625
+ laigc = 9.707156e-12
+ pbswgd = 0.95
+ pbswgs = 0.95
+ rnoia = 0
+ rnoib = 0
+ igcmod = 1
+ pketa = -6.053668000000001e-15
+ ngate = 8e+20
+ ngcon = 1
+ wpclm = 1.6305740000000013e-7
+ bigbacc = 0.002588
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ kvth0we = 0.00018
+ paigsd = -1.2154906e-23
+ lintnoi = -1.5e-8
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ ijthsfwd = 0.01
+ permod = 1
+ keta = -0.59506219
+ ijthsrev = 0.01
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = -4.4084e-11
+ tvoff = 0.0034020192
+ kt1l = 0
+ voffcv = -0.16942
+ wpemod = 1
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ lint = 0
+ lkt1 = -1.8529946e-8
+ lkt2 = 1.0897551e-9
+ lmax = 4.333e-8
+ lmin = 3.6e-8
+ ku0we = -0.0007
+ nfactor = 1
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ beta0 = 13
+ leta0 = 2.4927632200000002e-8
+ letab = 2.5974719e-8
+ minv = -0.3
+ lua1 = 7.6118385e-17
+ lub1 = -1.5665095e-25
+ luc1 = -2.1832442999999997e-17
+ ppclm = -8.780734400000002e-15
+ ndep = 1e+18
+ dlcig = 2.5e-9
+ lwlc = 0
+ tpbswg = 0.0009
+ bgidl = 2320000000.0
+ moin = 5.1
+ nigc = 3.083
+ nigbacc = 10
+ dmcgt = 0
+ pkvth0we = -1.3e-19
+ noff = 2.7195
+ tcjsw = 0.000357
+ ptvoff = -5.392468e-18
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ waigsd = 3.1116181e-12
+ nigbinv = 10
+ diomod = 1
+ ntox = -0.31099999999999994
+ pcit = 5.0236409e-17
+ vfbsdoff = 0.02
+ pclm = 1.46768105
+ bigsd = 0.00125
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 3.0174000000000004e-10
+ pku0we = -1.5e-18
+ cjswgs = 3.0174000000000004e-10
+ phin = 0.15
+ wvoff = -1.1108948e-8
+ paramchk = 1
+ pkt1 = 5.3710205e-15
+ pkt2 = -4.1883975e-17
+ wvsat = -0.03344995599999999
+ wvth0 = -2.2856158999999997e-8
+ fnoimod = 1
+ mjswgd = 0.85
+ mjswgs = 0.85
+ eigbinv = 1.1
+ waigc = 7.6854687e-11
+ tcjswg = 0.001
+ rbdb = 50
+ pua1 = -2.7889543e-23
+ prwb = 0
+ prwg = 0
+ pub1 = 5.5961859e-32
+ puc1 = 7.935933e-24
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ pvfbsdoff = 0
+ lketa = 1.80561909e-8
+ ijthdfwd = 0.01
+ rdsw = 100
+ xpart = 1
+ egidl = 0.29734
+ cigbacc = 0.32875
+ ijthdrev = 0.01
+ fprout = 300
+ rshg = 15.6
+ xrcrg1 = 12
+ xrcrg2 = 1
+ tnoimod = 0
+ cigbinv = 0.006
+ wtvoff = 7.822084e-11
+ pvoff = 6.821929600000002e-16
+ version = 4.5
+ capmod = 2
+ tnom = 25
+ cdscb = 0
+ cdscd = 0
+ tempmod = 0
+ toxe = 2.47e-9
+ toxm = 2.43e-9
+ pvsat = 1.20901182e-9
+ wku0we = 2e-11
+ lkvth0we = -2e-12
+ wk2we = 5e-12
+ pvth0 = 1.42910679e-15
+ drout = 0.56
+ mobmod = 0
+ wtvfbsdoff = 0
+ paigc = -2.6395467e-18
+ aigbacc = 0.02
+ voffl = 0
+ acnqsmod = 0
+ ltvfbsdoff = 0
+ weta0 = 8.5615058e-8
+ wetab = 2.2270081e-8
+ wags = 1.4953333e-7
+ lpclm = -1.8821805999999992e-8
+ wcit = -1.3198261000000002e-9
+ rbodymod = 0
+ aigbinv = 0.0163
+ voff = -0.04303087299999998
+ cgidl = 0.22
+ acde = 0.4
+ laigsd = 4.4039511e-17
+ vsat = 182708.442
+ wint = 0
+ vth0 = 0.399299171
+ wkt1 = -1.2366136999999998e-7
+ wkt2 = 7.8385579e-10
+ wmax = 5.426e-7
+ aigc = 0.011053515
+ wmin = 2.726e-7
+ pbswd = 0.8
+ pbsws = 0.8
+ ptvfbsdoff = 0
+ wpdiblc2 = 1.4081704e-10
+ wua1 = 6.7078609e-16
+ wub1 = -1.3253118999999999e-24
+ wuc1 = -1.9364911e-16
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ poxedge = 1
+ bigc = 0.001442
+ pdits = 0
+ wwlc = 0
+ cigsd = 0.069865
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ binunit = 2
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.0874977e-12
+ cgdo = 4.5622265999999996e-11
+ xtid = 3
+ xtis = 3
+ ags = 2.8144443999999997
+ cgsl = 3.0874977e-12
+ pk2we = -1e-19
+ cgso = 4.5622265999999996e-11
+ cigc = 0.000625
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ a0 = 10.55945905
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 51568.057
+ cf = 7.5795e-11
+ cjd = 0.00145199
+ cit = 0.0060336591999999994
+ cjs = 0.00145199
+ clc = 1e-7
+ ef = 1.0
+ k1 = 0.274
+ cle = 0.6
+ k2 = 0.041127322
+ k3 = -1.8419
+ em = 1000000.0
+ bvd = 8.7
+ bvs = 8.7
+ ll = 0
+ lw = 0
+ dlc = 3.26497e-9
+ u0 = 0.0085132265
+ w0 = 0
+ k3b = 1.9326
+ ua = -1.7148580999999998e-9
+ ub = 1.250859149999999e-18
+ uc = 5.4381728e-10
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 5.6700000000000005e-9
+ dwb = 0
+ ww = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ xw = 3.4e-9
+ wkvth0we = 2e-12
+ tnoia = 0
+ toxref = 3e-9
+ peta0 = -4.1184253e-15
+ la0 = -4.65319969e-7
+ trnqsmod = 0
+ petab = -7.719916e-16
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = 0.0013605251200000002
+ kt1 = 0.12069622
+ lk2 = -4.2131932e-9
+ kt2 = -0.11741295
+ wketa = 1.87190595e-7
+ llc = 0
+ lln = 1
+ lu0 = 1.1593053e-10
+ mjd = 0.26
+ lua = 1.6761980000000137e-18
+ mjs = 0.26
+ lub = 8.339062399999967e-27
+ luc = -2.98810456e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ tpbsw = 0.0019
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 9.065128000000001e-14
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ nsd = 1e+20
+ pbd = 0.52
+ pat = -1.54912428e-9
+ pbs = 0.52
+ pk2 = 5.9540883e-16
+ cjswd = 8.774000000000001e-11
+ cjsws = 8.774000000000001e-11
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ pu0 = -7.710994e-17
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ prt = 0
+ pua = -1.6092489999999997e-23
+ pub = 1.5276544400000003e-32
+ puc = 5.518326299999999e-24
+ pud = 0
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = -1.1935669e-9
+ ub1 = 2.7958892300000004e-18
+ uc1 = 6.286009700000002e-10
+ tpb = 0.0014
+ k2we = 5e-5
+ wa0 = -2.59429679e-6
+ tvfbsdoff = 0.022
+ ute = -1
+ wat = 0.0301316685
+ dsub = 0.75
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -1.1593839e-8
+ ltvoff = -1.1952424e-10
+ dtox = 2.7e-10
+ wlc = 0
+ wln = 1
+ rgatemod = 0
+ wu0 = 1.1265157e-9
+ xgl = -1.09e-8
+ xgw = 0
+ wua = 3.2583921000000013e-16
+ wub = -3.447615700000002e-25
+ wuc = -8.750290400000002e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ tnjtsswg = 1
+ )

.model nch_ss_33 nmos (
+ level = 54
+ rbodymod = 0
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ version = 4.5
+ pbswgd = 0.95
+ pbswgs = 0.95
+ ntox = -0.31099999999999994
+ pcit = 0
+ pclm = 1.8851852
+ tempmod = 0
+ igcmod = 1
+ phin = 0.15
+ aigbacc = 0.02
+ pkt1 = 0
+ wpdiblc2 = -2.9834e-10
+ pvoff = -7e-17
+ cdscb = 0
+ cdscd = 0
+ pvsat = 0
+ aigbinv = 0.0163
+ rbdb = 50
+ prwb = 0
+ prwg = 0
+ pub1 = 0
+ wk2we = 5e-12
+ pvth0 = 2.3e-16
+ drout = 0.56
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ rdsw = 100
+ permod = 1
+ voffl = 0
+ weta0 = 0
+ wkvth0we = 2e-12
+ cgidl = 0.22
+ trnqsmod = 0
+ voffcv = -0.16942
+ wpemod = 1
+ poxedge = 1
+ rshg = 15.6
+ binunit = 2
+ pbswd = 0.8
+ pbsws = 0.8
+ rgatemod = 0
+ tnjtsswg = 1
+ tnom = 25
+ pdits = 0
+ ags = 0.75882593
+ cigsd = 0.069865
+ toxe = 2.47e-9
+ toxm = 2.43e-9
+ tpbswg = 0.0009
+ cjd = 0.00145199
+ dvt0w = 0
+ cit = 0.002342713
+ dvt1w = 0
+ cjs = 0.00145199
+ clc = 1e-7
+ cle = 0.6
+ dvt2w = 0
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 9.8024918e-9
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ jtsswgd = 2.3e-7
+ pk2we = -1e-19
+ jtsswgs = 2.3e-7
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ la0 = 0
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = 0.0004
+ kt1 = -0.21767878
+ kt2 = -0.055117852
+ ptvoff = 0
+ llc = 0
+ lln = 1
+ lu0 = -6e-12
+ wags = 2.6994444e-8
+ mjd = 0.26
+ mjs = 0.26
+ lub = 0
+ lud = 0
+ lwc = 0
+ waigsd = 3.1789128e-12
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 0
+ tnoia = 0
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 6e-11
+ wcit = -2.5566928e-10
+ pbs = 0.52
+ pu0 = 0
+ prt = 0
+ pub = 0
+ pud = 0
+ peta0 = 0
+ diomod = 1
+ voff = -0.095952978
+ acde = 0.4
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 9.5347726e-10
+ wketa = -1.1490089e-9
+ ub1 = -5.3850981e-19
+ uc1 = -6.0041111e-11
+ tpb = 0.0014
+ tpbsw = 0.0019
+ pditsd = 0
+ pditsl = 0
+ vsat = 84306.193
+ wa0 = 0
+ cjswgd = 3.0174000000000004e-10
+ pku0we = -1.5e-18
+ cjswgs = 3.0174000000000004e-10
+ wint = 0
+ ute = -1
+ wat = 0
+ vth0 = 0.34069411000000005
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 3.0219344e-9
+ cjswd = 8.774000000000001e-11
+ cjsws = 8.774000000000001e-11
+ wlc = 0
+ wln = 1
+ wu0 = 4.3306667e-11
+ wkt1 = 3.0854175e-10
+ wkt2 = 1.0235511e-10
+ xgl = -1.09e-8
+ mjswd = 0.11
+ xgw = 0
+ mjsws = 0.11
+ wua = -1.6467997e-17
+ wub = 3.619626e-26
+ wuc = -1.4955111e-18
+ wud = 0
+ agidl = 9.41e-8
+ wmax = 2.726e-7
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ aigc = 0.01181895
+ wmin = 1.08e-7
+ tvfbsdoff = 0.022
+ njtsswg = 9
+ mjswgd = 0.85
+ mjswgs = 0.85
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ wua1 = -3.1223388e-18
+ wub1 = 2.0807554e-26
+ wuc1 = 8.1864667e-18
+ tcjswg = 0.001
+ bigc = 0.001442
+ ckappad = 0.6
+ ckappas = 0.6
+ wwlc = 0
+ pdiblc1 = 0
+ pdiblc2 = 0.023869018
+ pdiblcb = -0.3
+ scref = 1e-6
+ cdsc = 0
+ ijthsfwd = 0.01
+ cgbo = 0
+ cgdl = 3.0874977e-12
+ cgdo = 4.5622265999999996e-11
+ xtid = 3
+ xtis = 3
+ pigcd = 2.621
+ aigsd = 0.010772573
+ cgsl = 3.0874977e-12
+ cgso = 4.5622265999999996e-11
+ cigc = 0.000625
+ lvoff = 0
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ bigbacc = 0.002588
+ lvsat = 0.0003
+ lvth0 = 0
+ fprout = 300
+ ijthsrev = 0.01
+ delta = 0.007595625
+ xrcrg1 = 12
+ xrcrg2 = 1
+ kvth0we = 0.00018
+ rnoia = 0
+ rnoib = 0
+ lintnoi = -1.5e-8
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ wtvoff = 2.5061202e-10
+ ngate = 8e+20
+ wtvfbsdoff = 0
+ ngcon = 1
+ wpclm = -9.7111111e-9
+ k2we = 5e-5
+ dsub = 0.75
+ dtox = 2.7e-10
+ gbmin = 1e-12
+ capmod = 2
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ ltvfbsdoff = 0
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ wku0we = 2e-11
+ mobmod = 0
+ eta0 = 0.2
+ etab = -0.2
+ pkvth0we = -1.3e-19
+ nfactor = 1
+ ptvfbsdoff = 0
+ tvoff = 0.00085486634
+ vfbsdoff = 0.02
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ paramchk = 1
+ nigbacc = 10
+ ku0we = -0.0007
+ beta0 = 13
+ leta0 = 0
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ dlcig = 2.5e-9
+ nigbinv = 10
+ bgidl = 2320000000.0
+ ijthdfwd = 0.01
+ keta = -0.021050128
+ dmcgt = 0
+ tcjsw = 0.000357
+ toxref = 3e-9
+ ijthdrev = 0.01
+ fnoimod = 1
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 4e-12
+ eigbinv = 1.1
+ kt1l = 0
+ bigsd = 0.00125
+ lint = 6.5375218e-9
+ lkt1 = 0
+ wvoff = 2.9681533e-9
+ lmax = 2.001e-5
+ lmin = 8.99743e-6
+ ltvoff = 0
+ lpe0 = 9.2e-8
+ wvsat = 0.002322956
+ lpeb = 2.5e-7
+ wvth0 = -9.513738999999998e-10
+ a0 = 3.5
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 200000
+ cf = 7.5795e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.017956400999999997
+ k3 = -1.8419
+ em = 1000000.0
+ minv = -0.3
+ waigc = 1.7818122e-11
+ ll = 0
+ lw = 0
+ u0 = 0.013335556
+ w0 = 0
+ lub1 = 0
+ ua = -2.0911548e-9
+ ub = 2.2368542e-18
+ uc = 5.8018519e-11
+ ud = 0
+ cigbacc = 0.32875
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 5.6700000000000005e-9
+ ww = 0
+ xw = 3.4e-9
+ ndep = 1e+18
+ lkvth0we = -2e-12
+ pvfbsdoff = 0
+ lwlc = 0
+ moin = 5.1
+ lku0we = 2.5e-11
+ tnoimod = 0
+ epsrox = 3.9
+ xpart = 1
+ nigc = 3.083
+ cigbinv = 0.006
+ acnqsmod = 0
+ rdsmod = 0
+ egidl = 0.29734
+ igbmod = 1
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ )

.model nch_ss_34 nmos (
+ level = 54
+ paramchk = 1
+ wpclm = -9.7111111e-9
+ gbmin = 1e-12
+ wua1 = -1.7574281e-19
+ wub1 = 1.7597088e-26
+ wuc1 = 8.3134424e-18
+ jswgd = 1.28e-13
+ nfactor = 1
+ jswgs = 1.28e-13
+ paigsd = -3.8370159e-23
+ bigc = 0.001442
+ wwlc = 0
+ permod = 1
+ cdsc = 0
+ ijthdfwd = 0.01
+ cgbo = 0
+ cgdl = 3.0874977e-12
+ cgdo = 4.5622265999999996e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.0874977e-12
+ cgso = 4.5622265999999996e-11
+ cigc = 0.000625
+ nigbacc = 10
+ ijthdrev = 0.01
+ voffcv = -0.16942
+ wpemod = 1
+ tvoff = 0.00082419905
+ lpdiblc2 = -9.2950492e-9
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ nigbinv = 10
+ k2we = 5e-5
+ ku0we = -0.0007
+ beta0 = 13
+ dsub = 0.75
+ leta0 = 0
+ dtox = 2.7e-10
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ tpbswg = 0.0009
+ fnoimod = 1
+ lkvth0we = -2e-12
+ eigbinv = 1.1
+ dlcig = 2.5e-9
+ eta0 = 0.2
+ bgidl = 2320000000.0
+ etab = -0.2
+ acnqsmod = 0
+ ptvoff = -2.3727895e-16
+ waigsd = 3.1789171e-12
+ dmcgt = 0
+ tcjsw = 0.000357
+ rbodymod = 0
+ diomod = 1
+ cigbacc = 0.32875
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 3.0174000000000004e-10
+ pku0we = -1.5e-18
+ cjswgs = 3.0174000000000004e-10
+ bigsd = 0.00125
+ tnoimod = 0
+ wvoff = 3.141381e-9
+ mjswgd = 0.85
+ mjswgs = 0.85
+ cigbinv = 0.006
+ wvsat = 0.002322956
+ wvth0 = -1.1363659000000002e-9
+ wpdiblc2 = -6.4961636e-10
+ tcjswg = 0.001
+ waigc = 1.8291238e-11
+ pvfbsdoff = 0
+ version = 4.5
+ lketa = -2.7750915e-8
+ tempmod = 0
+ xpart = 1
+ egidl = 0.29734
+ aigbacc = 0.02
+ keta = -0.017963263
+ wkvth0we = 2e-12
+ wtvfbsdoff = 0
+ fprout = 300
+ lags = 4.3821463e-7
+ xrcrg1 = 12
+ xrcrg2 = 1
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = -5.265105499999999e-12
+ trnqsmod = 0
+ kt1l = 0
+ ltvfbsdoff = 0
+ aigbinv = 0.0163
+ wtvoff = 2.7700567e-10
+ lint = 6.5375218e-9
+ lkt1 = -8.8818468e-8
+ lkt2 = -1.6837724e-8
+ lmax = 8.99743e-6
+ lmin = 8.974099999999999e-7
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ capmod = 2
+ rgatemod = 0
+ pvoff = -1.6273171999999999e-15
+ tnjtsswg = 1
+ wku0we = 2e-11
+ minv = -0.3
+ lua1 = -7.4262143e-17
+ lub1 = -1.4158035e-25
+ luc1 = 6.2830403e-17
+ cdscb = 0
+ cdscd = 0
+ mobmod = 0
+ pvsat = 0
+ ndep = 1e+18
+ wk2we = 5e-12
+ pvth0 = 1.8930782e-15
+ ptvfbsdoff = 0
+ drout = 0.56
+ lwlc = 0
+ poxedge = 1
+ moin = 5.1
+ paigc = -4.2533129e-18
+ nigc = 3.083
+ voffl = 0
+ binunit = 2
+ weta0 = 0
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ laigsd = 3.3658034e-16
+ pags = 5.2134206e-15
+ cgidl = 0.22
+ ntox = -0.31099999999999994
+ pcit = 7.9881874e-17
+ pclm = 1.8851852
+ phin = 0.15
+ pbswd = 0.8
+ pbsws = 0.8
+ ags = 0.71008125
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ pkt1 = -3.6416964e-16
+ pkt2 = -1.7740443e-15
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ cjd = 0.00145199
+ cit = 0.0023437436
+ cjs = 0.00145199
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 9.8024918e-9
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ pdits = 0
+ cigsd = 0.069865
+ rbdb = 50
+ pua1 = -2.6489898e-23
+ prwb = 0
+ prwg = 0
+ pub1 = 2.886209e-32
+ puc1 = -1.1415122e-24
+ dvt0w = 0
+ la0 = -1.6207075e-6
+ dvt1w = 0
+ dvt2w = 0
+ rbpb = 50
+ rbpd = 50
+ jsd = 6.11e-7
+ rbps = 50
+ jss = 6.11e-7
+ lat = -0.042822769000000004
+ rbsb = 50
+ pvag = 1.2
+ kt1 = -0.20779908
+ lk2 = -1.5849432e-8
+ kt2 = -0.053244913
+ llc = 0
+ lln = 1
+ lu0 = -1.6852432e-9
+ mjd = 0.26
+ lua = -1.2813977e-16
+ mjs = 0.26
+ lub = -8.5009677e-26
+ luc = -2.2547224e-17
+ lud = 0
+ ijthsfwd = 0.01
+ lwc = 0
+ lwl = 0
+ rdsw = 100
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 3.8370159e-14
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 4.0504965e-9
+ pbs = 0.52
+ pk2 = -8.7965669e-16
+ pk2we = -1e-19
+ pu0 = -1.6281621e-30
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ prt = 0
+ pua = -3.3674591e-24
+ pub = -4.9159389e-33
+ puc = 2.3789498e-24
+ pud = 0
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 9.6173779e-10
+ ub1 = -5.2276116e-19
+ uc1 = -6.7030033e-11
+ njtsswg = 9
+ tpb = 0.0014
+ toxref = 3e-9
+ wa0 = -4.2680933e-9
+ tnoia = 0
+ ute = -1
+ wat = -0.0004438817
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 3.1197827e-9
+ wlc = 0
+ wln = 1
+ wu0 = 4.3306667e-11
+ ijthsrev = 0.01
+ xgl = -1.09e-8
+ xtsswgd = 0.18
+ xgw = 0
+ xtsswgs = 0.18
+ wua = -1.6093419e-17
+ wub = 3.6743083e-26
+ wuc = -1.7601329e-18
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ peta0 = 0
+ wketa = -1.4921751e-9
+ ckappad = 0.6
+ ckappas = 0.6
+ rshg = 15.6
+ pdiblc1 = 0
+ pdiblc2 = 0.02490295
+ tpbsw = 0.0019
+ pdiblcb = -0.3
+ cjswd = 8.774000000000001e-11
+ cjsws = 8.774000000000001e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ tvfbsdoff = 0.022
+ ltvoff = 2.7569894e-10
+ ppdiblc2 = 3.1579745e-15
+ bigbacc = 0.002588
+ tnom = 25
+ toxe = 2.47e-9
+ toxm = 2.43e-9
+ kvth0we = 0.00018
+ lku0we = 2.5e-11
+ epsrox = 3.9
+ scref = 1e-6
+ lintnoi = -1.5e-8
+ pigcd = 2.621
+ bigbinv = 0.004953
+ aigsd = 0.010772573
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ rdsmod = 0
+ wvfbsdoff = 0
+ igbmod = 1
+ lvoff = -1.4738881e-8
+ lvfbsdoff = 0
+ pkvth0we = -1.3e-19
+ wags = 2.6414531e-8
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ lvsat = 0.0003
+ wcit = -2.6455491e-10
+ lvth0 = 5.661542e-8
+ pbswgd = 0.95
+ pbswgs = 0.95
+ voff = -0.094313503
+ delta = 0.007595625
+ laigc = -1.6452737e-10
+ acde = 0.4
+ a0 = 3.6802789
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ vfbsdoff = 0.02
+ igcmod = 1
+ at = 204807.87
+ cf = 7.5795e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.019719408
+ k3 = -1.8419
+ em = 1000000.0
+ rnoia = 0
+ rnoib = 0
+ ll = 0
+ lw = 0
+ vsat = 84306.193
+ u0 = 0.013522346
+ w0 = 0
+ wint = 0
+ ua = -2.0769012e-9
+ ub = 2.2463102e-18
+ uc = 6.0526552e-11
+ ud = 0
+ vth0 = 0.33439651000000004
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 5.6700000000000005e-9
+ ww = 0
+ xw = 3.4e-9
+ wkt1 = 3.4905004999999996e-10
+ wkt2 = 2.996904e-10
+ wmax = 2.726e-7
+ aigc = 0.011837251
+ wmin = 1.08e-7
+ pketa = 3.0850638e-15
+ ngate = 8e+20
+ ngcon = 1
+ )

.model nch_ss_35 nmos (
+ level = 54
+ a0 = 2.7573663
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ voffl = 0
+ at = 225908.74
+ cf = 7.5795e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.012686581
+ k3 = -1.8419
+ em = 1000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.013112289999999999
+ w0 = 0
+ ua = -2.2251639e-9
+ ub = 2.3450974e-18
+ uc = 3.6825844e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 5.6700000000000005e-9
+ ww = 0
+ xw = 3.4e-9
+ weta0 = 0
+ keta = -0.063873893
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ voffcv = -0.16942
+ wpemod = 1
+ lags = -4.2829945e-7
+ ijthsrev = 0.01
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ cgidl = 0.22
+ lcit = -6.1490204e-10
+ kt1l = 0
+ ags = 1.6836926
+ cjd = 0.00145199
+ cit = 0.0030287289
+ cjs = 0.00145199
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 9.8024918e-9
+ k3b = 1.9326
+ lint = 6.5375218e-9
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ lkt1 = 4.9051427e-8
+ lkt2 = -1.4519819e-8
+ pbswd = 0.8
+ pbsws = 0.8
+ lmax = 8.974099999999999e-7
+ lmin = 4.4741e-7
+ lpe0 = 9.2e-8
+ la0 = -7.9931523e-7
+ lpeb = 2.5e-7
+ jsd = 6.11e-7
+ ppdiblc2 = -1.3141262e-15
+ jss = 6.11e-7
+ lat = -0.061602545
+ kt1 = -0.36270908
+ lk2 = -9.5902228e-9
+ kt2 = -0.0558493
+ llc = 0
+ lln = 1
+ lu0 = -1.3202934e-9
+ njtsswg = 9
+ mjd = 0.26
+ lua = 3.8140531e-18
+ mjs = 0.26
+ lub = -1.7293024e-25
+ luc = -1.4535934e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ tpbswg = 0.0009
+ njd = 1.02
+ minv = -0.3
+ njs = 1.02
+ pa0 = -6.7606598e-14
+ lua1 = -1.6437259e-16
+ lub1 = 2.2818043e-26
+ nsd = 1e+20
+ pdits = 0
+ luc1 = 5.6450349e-17
+ pbd = 0.52
+ pat = 1.7632657e-9
+ pbs = 0.52
+ pk2 = -2.3173279e-16
+ cigsd = 0.069865
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ pu0 = 8.9578742e-18
+ prt = 0
+ ndep = 1e+18
+ pua = -1.9061799e-24
+ pub = 1.3958464e-33
+ puc = -1.352132e-24
+ pud = 0
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ lwlc = 0
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 1.0629855e-9
+ ckappad = 0.6
+ ub1 = -7.0747845e-19
+ moin = 5.1
+ uc1 = -5.9861432e-11
+ ckappas = 0.6
+ tpb = 0.0014
+ pdiblc1 = 0
+ pdiblc2 = 0.01020022
+ pdiblcb = -0.3
+ wa0 = 1.1480691e-7
+ ute = -1
+ nigc = 3.083
+ wat = 0.0021260405
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 2.3917793e-9
+ wlc = 0
+ pk2we = -1e-19
+ ptvoff = -4.8469984e-16
+ wln = 1
+ wu0 = 3.3241639999999996e-11
+ xgl = -1.09e-8
+ dvtp0 = 4e-7
+ xgw = 0
+ dvtp1 = 0.01
+ wua = -1.7735306e-17
+ wub = 2.9651178e-26
+ wuc = 2.4320938e-18
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ waigsd = 3.178874e-12
+ pkvth0we = -1.3e-19
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ tnoia = 0
+ diomod = 1
+ bigbacc = 0.002588
+ peta0 = 0
+ pags = -9.2425378e-15
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 3.0174000000000004e-10
+ pku0we = -1.5e-18
+ cjswgs = 3.0174000000000004e-10
+ wketa = 5.5022601e-9
+ vfbsdoff = 0.02
+ ntox = -0.31099999999999994
+ pcit = 1.588079e-16
+ pclm = 1.8851852
+ tpbsw = 0.0019
+ kvth0we = 0.00018
+ cjswd = 8.774000000000001e-11
+ cjsws = 8.774000000000001e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ phin = 0.15
+ tvfbsdoff = 0.022
+ lintnoi = -1.5e-8
+ bigbinv = 0.004953
+ mjswgd = 0.85
+ mjswgs = 0.85
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ paramchk = 1
+ pkt1 = -1.3211355e-14
+ pkt2 = 1.7857928e-15
+ tcjswg = 0.001
+ wtvfbsdoff = 0
+ rbdb = 50
+ pua1 = 3.1539092e-23
+ prwb = 0
+ prwg = 0
+ pub1 = -3.1533886e-32
+ puc1 = -7.798421e-24
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ scref = 1e-6
+ ijthdfwd = 0.01
+ rdsw = 100
+ pigcd = 2.621
+ aigsd = 0.010772573
+ ltvfbsdoff = 0
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ lvoff = -2.8456354e-8
+ fprout = 300
+ lvsat = 0.0003
+ xrcrg1 = 12
+ xrcrg2 = 1
+ lvth0 = 1.8754806e-8
+ ijthdrev = 0.01
+ delta = 0.007595625
+ nfactor = 1
+ laigc = -6.1235169e-11
+ lpdiblc2 = 3.7903799e-9
+ rshg = 15.6
+ rnoia = 0
+ rnoib = 0
+ wtvoff = 5.5500668e-10
+ ptvfbsdoff = 0
+ pketa = -3.1399835e-15
+ ngate = 8e+20
+ ngcon = 1
+ wpclm = -9.7111111e-9
+ capmod = 2
+ wku0we = 2e-11
+ gbmin = 1e-12
+ nigbacc = 10
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ mobmod = 0
+ tnom = 25
+ toxe = 2.47e-9
+ toxm = 2.43e-9
+ lkvth0we = -2e-12
+ nigbinv = 10
+ acnqsmod = 0
+ wags = 4.2657181000000004e-8
+ rbodymod = 0
+ wcit = -3.5323584e-10
+ voff = -0.078900611
+ tvoff = -3.4914836e-5
+ acde = 0.4
+ fnoimod = 1
+ xjbvd = 1
+ xjbvs = 1
+ vsat = 84306.193
+ lk2we = -1.5e-12
+ eigbinv = 1.1
+ wint = 0
+ vth0 = 0.37693652
+ wkt1 = 1.478409e-8
+ wkt2 = -3.7001265e-9
+ wmax = 2.726e-7
+ aigc = 0.011721192
+ wmin = 1.08e-7
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ ku0we = -0.0007
+ beta0 = 13
+ leta0 = 0
+ wpdiblc2 = 4.3752159e-9
+ wua1 = -6.5376855e-17
+ wub1 = 8.5457734e-26
+ wuc1 = 1.5793115e-17
+ bigc = 0.001442
+ wwlc = 0
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ cigbacc = 0.32875
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.0874977e-12
+ cgdo = 4.5622265999999996e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.0874977e-12
+ cgso = 4.5622265999999996e-11
+ tnoimod = 0
+ cigc = 0.000625
+ toxref = 3e-9
+ dmcgt = 0
+ tcjsw = 0.000357
+ wkvth0we = 2e-12
+ cigbinv = 0.006
+ trnqsmod = 0
+ bigsd = 0.00125
+ version = 4.5
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ tempmod = 0
+ ltvoff = 1.0403103e-9
+ wvoff = -2.1121636e-9
+ k2we = 5e-5
+ wvsat = 0.002322956
+ aigbacc = 0.02
+ dsub = 0.75
+ wvth0 = 2.3985259e-9
+ dtox = 2.7e-10
+ rgatemod = 0
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ tnjtsswg = 1
+ waigc = 1.00872e-11
+ pvfbsdoff = 0
+ lku0we = 2.5e-11
+ epsrox = 3.9
+ eta0 = 0.2
+ etab = -0.2
+ lketa = 1.3109546e-8
+ aigbinv = 0.0163
+ xpart = 1
+ rdsmod = 0
+ igbmod = 1
+ egidl = 0.29734
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ pbswgd = 0.95
+ pbswgs = 0.95
+ igcmod = 1
+ poxedge = 1
+ binunit = 2
+ pvoff = 3.0483375000000002e-15
+ cdscb = 0
+ cdscd = 0
+ pvsat = 0
+ wk2we = 5e-12
+ pvth0 = -1.2529756000000001e-15
+ drout = 0.56
+ permod = 1
+ paigc = 3.0482801e-18
+ ijthsfwd = 0.01
+ )

.model nch_ss_36 nmos (
+ level = 54
+ rshg = 15.6
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ cigbacc = 0.32875
+ tnoimod = 0
+ ku0we = -0.0007
+ a0 = 2.8517872
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ beta0 = 13
+ at = 72186.119
+ cf = 7.5795e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.0061801551
+ k3 = -1.8419
+ em = 1000000.0
+ leta0 = 0
+ rgatemod = 0
+ ll = -1.18e-13
+ lw = 0
+ u0 = 0.011328434
+ tpbswg = 0.0009
+ w0 = 0
+ ua = -2.2247872e-9
+ ub = 2.0937783e-18
+ uc = 7.1203963e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 5.6700000000000005e-9
+ tnjtsswg = 1
+ ww = 0
+ xw = 3.4e-9
+ cigbinv = 0.006
+ tnom = 25
+ ppclm = 2.75592e-14
+ toxe = 2.47e-9
+ toxm = 2.43e-9
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ ptvoff = 2.8225911e-16
+ version = 4.5
+ waigsd = 3.178874e-12
+ tempmod = 0
+ dmcgt = 0
+ tcjsw = 0.000357
+ diomod = 1
+ wags = 2.560818e-7
+ aigbacc = 0.02
+ wcit = 1.8683634e-10
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 3.0174000000000004e-10
+ pku0we = -1.5e-18
+ cjswgs = 3.0174000000000004e-10
+ voff = -0.13810998
+ acde = 0.4
+ bigsd = 0.00125
+ vsat = 84306.193
+ wint = 0
+ vth0 = 0.43955442
+ wtvfbsdoff = 0
+ wkt1 = -3.7370623e-8
+ wkt2 = -4.3121065e-11
+ aigbinv = 0.0163
+ wmax = 2.726e-7
+ mjswgd = 0.85
+ mjswgs = 0.85
+ aigc = 0.011581706
+ wmin = 1.08e-7
+ wvoff = 7.1640927e-9
+ tcjswg = 0.001
+ wvsat = 0.002322956
+ ltvfbsdoff = 0
+ wvth0 = -3.3496131e-9
+ wua1 = 2.3276683e-17
+ wub1 = 1.5603072e-26
+ wuc1 = -5.1034561e-18
+ waigc = 2.6093343e-11
+ pvfbsdoff = 0
+ bigc = 0.001442
+ wwlc = 0
+ lketa = -3.8407777e-8
+ ijthsfwd = 0.01
+ cdsc = 0
+ xpart = 1
+ cgbo = 0
+ cgdl = 3.0874977e-12
+ cgdo = 4.5622265999999996e-11
+ xtid = 3
+ xtis = 3
+ poxedge = 1
+ cgsl = 3.0874977e-12
+ cgso = 4.5622265999999996e-11
+ cigc = 0.000625
+ egidl = 0.29734
+ fprout = 300
+ ptvfbsdoff = 0
+ binunit = 2
+ xrcrg1 = 12
+ xrcrg2 = 1
+ ijthsrev = 0.01
+ wtvoff = -1.1880818e-9
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ capmod = 2
+ k2we = 5e-5
+ wku0we = 2e-11
+ ppdiblc2 = 3.3310302e-16
+ dsub = 0.75
+ dtox = 2.7e-10
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ pvoff = -1.03321526e-15
+ mobmod = 0
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ cdscb = 0
+ cdscd = 0
+ pvsat = 0
+ wk2we = 5e-12
+ pvth0 = 1.2762056e-15
+ drout = 0.56
+ eta0 = 0.2
+ etab = -0.2
+ paigc = -3.9944226e-18
+ voffl = 0
+ weta0 = 0
+ pkvth0we = -1.3e-19
+ ags = -2.5047885
+ lpclm = -2.4174737e-7
+ cjd = 0.00145199
+ cit = 0.00083484714
+ cjs = 0.00145199
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 1.30529375e-8
+ k3b = 1.9326
+ njtsswg = 9
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ cgidl = 0.22
+ vfbsdoff = 0.02
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ la0 = -8.4086042e-7
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = 0.0060354098000000005
+ kt1 = -0.088256509
+ lk2 = -6.7273888e-9
+ kt2 = -0.075738087
+ ckappad = 0.6
+ ckappas = 0.6
+ llc = -1.18e-13
+ lln = 0.7
+ lu0 = -5.3539671e-10
+ mjd = 0.26
+ pdiblc1 = 0
+ pdiblc2 = 0.031716534
+ lua = 3.6483177e-18
+ mjs = 0.26
+ lub = -6.2349821e-26
+ luc = -1.6579966e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ pdiblcb = -0.3
+ njd = 1.02
+ njs = 1.02
+ pa0 = 8.661463e-14
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ pbswd = 0.8
+ pbsws = 0.8
+ nsd = 1e+20
+ pbd = 0.52
+ pat = -3.0818679e-9
+ pbs = 0.52
+ pk2 = -2.2869691e-16
+ paramchk = 1
+ pu0 = 2.4409578e-18
+ prt = 0
+ pua = -4.9144669e-25
+ pub = 1.8790045e-33
+ puc = 1.8346553e-24
+ pud = 0
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 5.8363721e-10
+ ub1 = -5.3348382e-19
+ uc1 = 8.6067289e-11
+ tpb = 0.0014
+ wa0 = -2.3569588e-7
+ ute = -1
+ wat = 0.013137708
+ pdits = 0
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 2.3848778e-9
+ wlc = 0
+ wln = 1
+ cigsd = 0.069865
+ wu0 = 4.8052813e-11
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -2.0950609e-17
+ wub = 2.8553091e-26
+ wuc = -4.8106046e-18
+ wud = 0
+ wwc = 0
+ bigbacc = 0.002588
+ wwl = 0
+ wwn = 1
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ ijthdfwd = 0.01
+ kvth0we = 0.00018
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ toxref = 3e-9
+ lintnoi = -1.5e-8
+ keta = 0.053210932
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ tnoia = 0
+ lags = 1.4146322e-6
+ ijthdrev = 0.01
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ peta0 = 0
+ lcit = 3.5040592e-10
+ wketa = -7.2433388e-9
+ kt1l = 0
+ lpdiblc2 = -5.676798e-9
+ tpbsw = 0.0019
+ cjswd = 8.774000000000001e-11
+ cjsws = 8.774000000000001e-11
+ mjswd = 0.11
+ tvfbsdoff = 0.022
+ mjsws = 0.11
+ ltvoff = -1.663256e-9
+ agidl = 9.41e-8
+ lint = 9.7879675e-9
+ lkt1 = -7.1707703e-8
+ lkt2 = -5.7687528e-9
+ lmax = 4.4741e-7
+ lmin = 2.1410000000000002e-7
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ minv = -0.3
+ lku0we = 2.5e-11
+ lua1 = 4.6540649e-17
+ lub1 = -5.3739597e-26
+ luc1 = -7.7582888e-18
+ epsrox = 3.9
+ lkvth0we = -2e-12
+ ndep = 1e+18
+ nfactor = 1
+ lwlc = 0
+ moin = 5.1
+ scref = 1e-6
+ rdsmod = 0
+ pigcd = 2.621
+ nigc = 3.083
+ igbmod = 1
+ aigsd = 0.010772573
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ acnqsmod = 0
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ lvoff = -2.4042325e-9
+ pbswgd = 0.95
+ noff = 2.7195
+ pbswgs = 0.95
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ lvsat = 0.0003
+ rbodymod = 0
+ lvth0 = -8.7970687e-9
+ igcmod = 1
+ nigbacc = 10
+ delta = 0.007595625
+ pags = -1.0314937e-13
+ laigc = 1.3898222e-13
+ ntox = -0.31099999999999994
+ pcit = -7.882386e-17
+ pclm = 2.434611
+ rnoia = 0
+ rnoib = 0
+ phin = 0.15
+ pketa = 2.46808e-15
+ ngate = 8e+20
+ nigbinv = 10
+ ngcon = 1
+ wpclm = -7.2345657e-8
+ pkt1 = 9.7367187e-15
+ pkt2 = 1.7671038e-16
+ wpdiblc2 = 6.3151306e-10
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ permod = 1
+ rbdb = 50
+ pua1 = -7.4684646e-24
+ prwb = 0
+ prwg = 0
+ pub1 = -7.978346e-34
+ puc1 = 1.3960704e-24
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ fnoimod = 1
+ rdsw = 100
+ eigbinv = 1.1
+ wkvth0we = 2e-12
+ voffcv = -0.16942
+ wpemod = 1
+ trnqsmod = 0
+ tvoff = 0.006109554
+ )

.model nch_ss_37 nmos (
+ level = 54
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ pdits = 0
+ cigsd = 0.069865
+ lkvth0we = -2e-12
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ eta0 = 0.2
+ etab = -0.2
+ ptvoff = -1.8615536e-17
+ waigsd = 3.178874e-12
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ acnqsmod = 0
+ diomod = 1
+ wtvfbsdoff = 0
+ tnoia = 0
+ pditsd = 0
+ pditsl = 0
+ rbodymod = 0
+ cjswgd = 3.0174000000000004e-10
+ pku0we = -1.5e-18
+ cjswgs = 3.0174000000000004e-10
+ a0 = -2.4455841
+ a1 = 0
+ a2 = 1
+ peta0 = 0
+ b0 = 0
+ b1 = 0
+ ltvfbsdoff = 0
+ at = 121458.51
+ cf = 7.5795e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = -0.0033973019999999996
+ k3 = -1.8419
+ em = 1000000.0
+ ll = -1.18e-13
+ wketa = 1.2169685000000001e-8
+ lw = 0
+ u0 = 0.009724212999999999
+ w0 = 0
+ ua = -2.2679307e-9
+ ub = 1.903479518e-18
+ uc = 2.5998306e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 5.6700000000000005e-9
+ ww = 0
+ xw = 3.4e-9
+ tpbsw = 0.0019
+ nfactor = 1
+ tvfbsdoff = 0.022
+ cjswd = 8.774000000000001e-11
+ cjsws = 8.774000000000001e-11
+ mjswgd = 0.85
+ mjswd = 0.11
+ mjswgs = 0.85
+ mjsws = 0.11
+ agidl = 9.41e-8
+ tcjswg = 0.001
+ wpdiblc2 = 2.0871493e-9
+ ptvfbsdoff = 0
+ nigbacc = 10
+ scref = 1e-6
+ wvfbsdoff = 0
+ pigcd = 2.621
+ lvfbsdoff = 0
+ aigsd = 0.010772573
+ fprout = 300
+ lvoff = 6.451419999999991e-11
+ nigbinv = 10
+ keta = -0.10792277
+ xrcrg1 = 12
+ xrcrg2 = 1
+ wkvth0we = 2e-12
+ lvsat = 0.000865079705
+ lvth0 = -7.861937700000001e-9
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ trnqsmod = 0
+ delta = 0.007595625
+ lcit = -3.5333293000000003e-11
+ wtvoff = 2.3786433e-10
+ laigc = -6.7426314e-12
+ kt1l = 0
+ rnoia = 0
+ rnoib = 0
+ fnoimod = 1
+ lint = 9.7879675e-9
+ pketa = -1.6280779999999998e-15
+ ngate = 8e+20
+ capmod = 2
+ eigbinv = 1.1
+ lkt1 = 5.5879381e-10
+ lkt2 = 1.6714521e-10
+ lmax = 2.1410000000000002e-7
+ ngcon = 1
+ lmin = 8.833e-8
+ wpclm = 1.5314007e-7
+ wku0we = 2e-11
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ mobmod = 0
+ rgatemod = 0
+ gbmin = 1e-12
+ tnjtsswg = 1
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ minv = -0.3
+ lua1 = -6.7367772e-18
+ lub1 = -3.8361216e-26
+ luc1 = -1.0970607e-17
+ ndep = 1e+18
+ lwlc = 0
+ moin = 5.1
+ nigc = 3.083
+ cigbacc = 0.32875
+ tnoimod = 0
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ cigbinv = 0.006
+ tvoff = -0.0028392003
+ ntox = -0.31099999999999994
+ pcit = 1.4940572e-17
+ pclm = 1.0592301
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ phin = 0.15
+ version = 4.5
+ tempmod = 0
+ pkt1 = -1.8629533e-16
+ pkt2 = -2.0087744e-16
+ ku0we = -0.0007
+ beta0 = 13
+ leta0 = 0
+ ppclm = -2.0018289e-14
+ aigbacc = 0.02
+ rbdb = 50
+ pua1 = 2.2068447e-24
+ prwb = 0
+ prwg = 0
+ pub1 = -2.7426774e-33
+ puc1 = 1.8773731e-24
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ ijthsfwd = 0.01
+ rdsw = 100
+ toxref = 3e-9
+ aigbinv = 0.0163
+ dmcgt = 0
+ tcjsw = 0.000357
+ ijthsrev = 0.01
+ rshg = 15.6
+ bigsd = 0.00125
+ ltvoff = 2.2493116e-10
+ wvoff = 1.8056166e-9
+ poxedge = 1
+ wvsat = 0.00305175308
+ ppdiblc2 = 2.596377e-17
+ wvth0 = 2.3151897e-9
+ binunit = 2
+ pvfbsdoff = 0
+ lku0we = 2.5e-11
+ waigc = 5.3999849e-12
+ tnom = 25
+ epsrox = 3.9
+ toxe = 2.47e-9
+ toxm = 2.43e-9
+ rdsmod = 0
+ lketa = -4.408530899999999e-9
+ igbmod = 1
+ xpart = 1
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ egidl = 0.29734
+ pbswgd = 0.95
+ pbswgs = 0.95
+ pkvth0we = -1.3e-19
+ wags = -2.3277778e-7
+ igcmod = 1
+ wcit = -2.5754486e-10
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ voff = -0.149810363
+ acde = 0.4
+ vfbsdoff = 0.02
+ vsat = 81628.05359999998
+ wint = 0
+ vth0 = 0.43512263300000004
+ wkt1 = 9.657879099999999e-9
+ wkt2 = 1.7463947e-9
+ wmax = 2.726e-7
+ aigc = 0.01161432
+ wmin = 1.08e-7
+ paramchk = 1
+ pvoff = 9.741822000000004e-17
+ wua1 = -2.2577864e-17
+ wub1 = 2.4820337e-26
+ wuc1 = -7.3845115e-18
+ cdscb = 0
+ cdscd = 0
+ bigc = 0.001442
+ permod = 1
+ pvsat = -1.5376888e-10
+ wwlc = 0
+ njtsswg = 9
+ wk2we = 5e-12
+ pvth0 = 8.093938e-17
+ drout = 0.56
+ ags = 4.199629600000001
+ paigc = 3.7187593e-19
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ ijthdfwd = 0.01
+ cdsc = 0
+ cjd = 0.00145199
+ cit = 0.0026629951
+ cgbo = 0
+ cjs = 0.00145199
+ clc = 1e-7
+ cle = 0.6
+ voffl = 0
+ cgdl = 3.0874977e-12
+ bvd = 8.7
+ cgdo = 4.5622265999999996e-11
+ xtid = 3
+ bvs = 8.7
+ xtis = 3
+ dlc = 1.30529375e-8
+ ckappad = 0.6
+ ckappas = 0.6
+ k3b = 1.9326
+ cgsl = 3.0874977e-12
+ cgso = 4.5622265999999996e-11
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ cigc = 0.000625
+ pdiblc1 = 0
+ pdiblc2 = 0.0095469071
+ pdiblcb = -0.3
+ weta0 = 0
+ voffcv = -0.16942
+ wpemod = 1
+ lpclm = 4.8457997e-8
+ la0 = 2.768849e-7
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.0043610641
+ kt1 = -0.43075175
+ lk2 = -4.7065454e-9
+ kt2 = -0.10387031
+ ijthdrev = 0.01
+ llc = -1.18e-13
+ lln = 0.7
+ lu0 = -1.9690617e-10
+ mjd = 0.26
+ mjs = 0.26
+ lua = 1.2751594e-17
+ lub = -2.21968369e-26
+ cgidl = 0.22
+ luc = -7.0415723e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = -2.9632335e-14
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 5.625644e-10
+ pbs = 0.52
+ pk2 = 3.1759465e-16
+ lpdiblc2 = -9.9900678e-10
+ pu0 = 4.2802262e-19
+ bigbacc = 0.002588
+ prt = 0
+ pua = 3.9870432e-24
+ pub = -6.31495433e-33
+ puc = 2.2635812e-25
+ pud = 0
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 8.3613685e-10
+ ub1 = -6.0636714e-19
+ uc1 = 1.0129155e-10
+ tpb = 0.0014
+ wa0 = 3.1523761e-7
+ kvth0we = 0.00018
+ pbswd = 0.8
+ pbsws = 0.8
+ ute = -1
+ wat = -0.0041344832
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -2.0418175e-10
+ wlc = 0
+ wln = 1
+ wu0 = 5.759279e-11
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -4.2175679e-17
+ wub = 6.73870221e-26
+ wuc = 2.8116572e-18
+ wud = 0
+ k2we = 5e-5
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ lintnoi = -1.5e-8
+ tpbswg = 0.0009
+ dsub = 0.75
+ bigbinv = 0.004953
+ dtox = 2.7e-10
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ )

.model nch_ss_38 nmos (
+ level = 54
+ dmcgt = 0
+ poxedge = 1
+ pkvth0we = -1.3e-19
+ tcjsw = 0.000357
+ pditsd = 0
+ pditsl = 0
+ noff = 2.7195
+ cjswgd = 3.0174000000000004e-10
+ pku0we = -1.5e-18
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ cjswgs = 3.0174000000000004e-10
+ binunit = 2
+ vfbsdoff = 0.02
+ ntox = -0.31099999999999994
+ pcit = 7.5496361e-18
+ pclm = 2.2357699
+ bigsd = 0.00125
+ ptvfbsdoff = 0
+ mjswgd = 0.85
+ mjswgs = 0.85
+ tcjswg = 0.001
+ phin = 0.15
+ wvoff = 4.874463324000002e-9
+ paramchk = 1
+ pkt1 = -2.4505624e-15
+ pkt2 = 3.9546557e-16
+ wvsat = 0.001769474099999998
+ wvth0 = 8.374116600000003e-9
+ pvfbsdoff = 0
+ waigc = -1.2918923e-11
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ rbdb = 50
+ pua1 = -4.7371604e-25
+ prwb = 0
+ pub1 = 4.7307687999999995e-33
+ prwg = 0
+ puc1 = -4.218097e-24
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ lketa = 3.8815738e-8
+ a0 = 0.7744856
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ ijthdfwd = 0.01
+ at = 98941.55040000001
+ cf = 7.5795e-11
+ xpart = 1
+ ef = 1.0
+ k1 = 0.274
+ k2 = -0.041338197
+ k3 = -1.8419
+ em = 1000000.0
+ rdsw = 100
+ ll = 0
+ lw = 0
+ u0 = 0.0052944609
+ w0 = 0
+ ua = -2.6695158e-9
+ ub = 2.0926996330000003e-18
+ uc = -9.6044814e-11
+ ud = 0
+ fprout = 300
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 5.6700000000000005e-9
+ ww = 0
+ xw = 3.4e-9
+ xrcrg1 = 12
+ xrcrg2 = 1
+ egidl = 0.29734
+ ijthdrev = 0.01
+ wtvoff = 2.7545299e-10
+ lpdiblc2 = 4.9724259e-14
+ rshg = 15.6
+ njtsswg = 9
+ capmod = 2
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ wku0we = 2e-11
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = -0.0010813536
+ mobmod = 0
+ pdiblcb = -0.3
+ ags = 4.199629600000001
+ pvoff = -1.910533700000002e-16
+ cjd = 0.00145199
+ cit = 0.0011085924
+ cjs = 0.00145199
+ clc = 1e-7
+ cle = 0.6
+ cdscb = 0
+ cdscd = 0
+ bvd = 8.7
+ tnom = 25
+ bvs = 8.7
+ dlc = 3.26497e-9
+ pvsat = -3.323489999999998e-11
+ k3b = 1.9326
+ lkvth0we = -2e-12
+ wk2we = 5e-12
+ toxe = 2.47e-9
+ dwb = 0
+ dwc = 0
+ toxm = 2.43e-9
+ dwg = 0
+ dwj = 0
+ pvth0 = -4.886005e-16
+ drout = 0.56
+ paigc = 2.0938533e-18
+ bigbacc = 0.002588
+ la0 = -2.5801646e-8
+ voffl = 0
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.00224447035
+ kt1 = -0.62571779
+ kt2 = -0.068117715
+ lk2 = -1.1401013e-9
+ llc = 0
+ lln = 1
+ lu0 = 2.1949052e-10
+ mjd = 0.26
+ acnqsmod = 0
+ mjs = 0.26
+ lua = 5.0500592e-17
+ lub = -3.9983527e-26
+ luc = 4.4304811e-18
+ lud = 0
+ laigsd = 1.06572e-17
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ kvth0we = 0.00018
+ weta0 = 4.2794074e-8
+ pa0 = 2.9413877e-15
+ wetab = -1.5859302e-8
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 5.166446900000001e-10
+ pbs = 0.52
+ pk2 = 2.316472e-16
+ lpclm = -6.2136744e-8
+ pu0 = -4.6164555e-17
+ wags = -2.3277778e-7
+ prt = 0
+ pua = -3.0159915e-24
+ pub = 1.3943639e-33
+ puc = 2.394639e-25
+ pud = 0
+ lintnoi = -1.5e-8
+ rbodymod = 0
+ wcit = -1.7891793699999998e-10
+ bigbinv = 0.004953
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 7.2026227e-10
+ vtsswgd = 4.2
+ ub1 = -6.260082000000002e-19
+ vtsswgs = 4.2
+ uc1 = -2.7209866e-10
+ cgidl = 0.22
+ tpb = 0.0014
+ wa0 = -3.1291358e-8
+ voff = -0.11849200800000002
+ ute = -1
+ wat = -0.00364597396
+ acde = 0.4
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 7.1015279e-10
+ wlc = 0
+ wln = 1
+ wu0 = 5.532584400000001e-10
+ xgl = -1.09e-8
+ xgw = 0
+ wua = 3.2324691e-17
+ wub = -1.4627000299999995e-26
+ wuc = 2.6722336e-18
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ vsat = 72365.62299999999
+ wint = 0
+ vth0 = 0.2829285080000001
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ wkt1 = 3.3745826e-8
+ wkt2 = -4.5976799e-9
+ wmax = 2.726e-7
+ aigc = 0.011905208
+ wmin = 1.08e-7
+ pbswd = 0.8
+ pbsws = 0.8
+ wpdiblc2 = 2.3634934e-9
+ wua1 = 5.9387403e-18
+ wub1 = -5.4684426e-26
+ wuc1 = 5.7460914e-17
+ pdits = 0
+ bigc = 0.001442
+ cigsd = 0.069865
+ wwlc = 0
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ cdsc = 0
+ nfactor = 1
+ toxref = 3e-9
+ cgbo = 0
+ cgdl = 3.0874977e-12
+ cgdo = 4.5622265999999996e-11
+ xtid = 3
+ xtis = 3
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ cgsl = 3.0874977e-12
+ cgso = 4.5622265999999996e-11
+ cigc = 0.000625
+ wkvth0we = 2e-12
+ tnoia = 0
+ peta0 = -4.0226429e-15
+ trnqsmod = 0
+ petab = 1.4907744e-15
+ wketa = 2.7230814999999998e-8
+ tpbsw = 0.0019
+ ltvoff = 1.3417313e-10
+ nigbacc = 10
+ tvfbsdoff = 0.022
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ cjswd = 8.774000000000001e-11
+ cjsws = 8.774000000000001e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ k2we = 5e-5
+ nigbinv = 10
+ dsub = 0.75
+ rgatemod = 0
+ lku0we = 2.5e-11
+ dtox = 2.7e-10
+ tnjtsswg = 1
+ epsrox = 3.9
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ rdsmod = 0
+ eta0 = -0.13238438
+ etab = 0.18670848
+ igbmod = 1
+ scref = 1e-6
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ pigcd = 2.621
+ aigsd = 0.010772573
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ fnoimod = 1
+ pbswgd = 0.95
+ pbswgs = 0.95
+ eigbinv = 1.1
+ lvoff = -2.8794112000000013e-9
+ igcmod = 1
+ lvsat = 0.0017357541499999996
+ lvth0 = 6.444309499999999e-9
+ delta = 0.007595625
+ laigc = -3.4086068e-11
+ rnoia = 0
+ rnoib = 0
+ pketa = -3.0438220100000003e-15
+ ngate = 8e+20
+ paigsd = -2.9413875e-24
+ ngcon = 1
+ cigbacc = 0.32875
+ wpclm = -8.3073835e-8
+ gbmin = 1e-12
+ tnoimod = 0
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ permod = 1
+ cigbinv = 0.006
+ ijthsfwd = 0.01
+ voffcv = -0.16942
+ wpemod = 1
+ version = 4.5
+ keta = -0.56775528
+ tempmod = 0
+ ijthsrev = 0.01
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 1.1078059e-10
+ tvoff = -0.0018736893
+ aigbacc = 0.02
+ kt1l = 0
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ lint = 0
+ lkt1 = 1.8885602e-8
+ lkt2 = -3.1935983e-9
+ lmax = 8.833e-8
+ lmin = 5.233e-8
+ tpbswg = 0.0009
+ ku0we = -0.0007
+ aigbinv = 0.0163
+ beta0 = 13
+ lpe0 = 9.2e-8
+ ppdiblc2 = -1.2574432e-20
+ lpeb = 2.5e-7
+ leta0 = 3.1244132e-8
+ letab = -3.6350598e-8
+ wtvfbsdoff = 0
+ minv = -0.3
+ ppclm = 2.1858187e-15
+ lua1 = 4.1554342e-18
+ lub1 = -3.6515003e-26
+ luc1 = 2.4128073e-17
+ ndep = 1e+18
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ ptvoff = -2.2148869e-17
+ lwlc = 0
+ moin = 5.1
+ ltvfbsdoff = 0
+ waigsd = 3.1789053e-12
+ nigc = 3.083
+ diomod = 1
+ )

.model nch_ss_39 nmos (
+ level = 54
+ wkt1 = 7.160945e-9
+ wkt2 = 1.1625249e-8
+ wmax = 2.726e-7
+ aigc = 0.011615807
+ wmin = 1.08e-7
+ fnoimod = 1
+ eigbinv = 1.1
+ wua1 = -1.0774777e-16
+ wub1 = 2.8568729000000003e-25
+ wuc1 = 2.134869e-17
+ bigc = 0.001442
+ wwlc = 0
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ scref = 1e-6
+ ijthsfwd = 0.01
+ cdsc = 0
+ fprout = 300
+ pigcd = 2.621
+ cgbo = 0
+ aigsd = 0.010772573
+ cgdl = 3.0874977e-12
+ cgdo = 4.5622265999999996e-11
+ xtid = 3
+ xtis = 3
+ xrcrg1 = 12
+ xrcrg2 = 1
+ cgsl = 3.0874977e-12
+ cgso = 4.5622265999999996e-11
+ cigc = 0.000625
+ lvoff = -6.4884398999999995e-9
+ cigbacc = 0.32875
+ lvsat = -0.0029471140999999994
+ wtvoff = 7.91509e-11
+ lvth0 = 6.355232699999999e-9
+ ijthsrev = 0.01
+ tnoimod = 0
+ delta = 0.007595625
+ laigc = -1.730084e-11
+ rnoia = 0
+ rnoib = 0
+ cigbinv = 0.006
+ dmcg = 3.1e-8
+ capmod = 2
+ dmci = 3.1e-8
+ dmdg = 0
+ wku0we = 2e-11
+ pketa = 5.517686e-15
+ ngate = 8e+20
+ a0 = 19.191807
+ a1 = 0
+ a2 = 1
+ ngcon = 1
+ b0 = 0
+ b1 = 0
+ mobmod = 0
+ wpclm = -5.2664346e-8
+ at = 93149.89199999998
+ cf = 7.5795e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = -0.055713829
+ k3 = -1.8419
+ em = 1000000.0
+ k2we = 5e-5
+ ll = 0
+ lw = 0
+ u0 = 0.0032278555
+ w0 = 0
+ ua = -2.3710013e-9
+ ub = 1.4550579529999998e-18
+ uc = -1.4785261e-10
+ ud = 0
+ version = 4.5
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 5.6700000000000005e-9
+ ww = 0
+ xw = 3.4e-9
+ dsub = 0.75
+ dtox = 2.7e-10
+ gbmin = 1e-12
+ tempmod = 0
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ eta0 = 1.1504337
+ aigbacc = 0.02
+ etab = -1.3364008
+ pkvth0we = -1.3e-19
+ aigbinv = 0.0163
+ tvoff = -0.0045522389
+ vfbsdoff = 0.02
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ paramchk = 1
+ ku0we = -0.0007
+ beta0 = 13
+ leta0 = -4.3159315e-8
+ poxedge = 1
+ letab = 5.198974e-8
+ ppclm = 4.2206835e-16
+ binunit = 2
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ ijthdfwd = 0.01
+ toxref = 3e-9
+ dmcgt = 0
+ keta = 0.47864502999999997
+ tcjsw = 0.000357
+ ijthdrev = 0.01
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 4.8801133e-10
+ ltvoff = 2.8952901e-10
+ kt1l = 0
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ bigsd = 0.00125
+ lint = 0
+ wvoff = -2.2288246e-9
+ lkt1 = 1.0413925e-8
+ lkt2 = 8.1983323e-9
+ lmax = 5.233e-8
+ lmin = 4.333e-8
+ wvsat = -0.012853907800000001
+ lku0we = 2.5e-11
+ pvfbsdoff = 0
+ lpe0 = 9.2e-8
+ wvth0 = -1.0255132099999999e-8
+ lpeb = 2.5e-7
+ epsrox = 3.9
+ waigc = 4.0939876e-11
+ minv = -0.3
+ lua1 = -3.9796071e-17
+ lub1 = 8.382587100000001e-26
+ luc1 = 1.26018728e-18
+ rdsmod = 0
+ lkvth0we = -2e-12
+ ndep = 1e+18
+ igbmod = 1
+ lwlc = 0
+ lketa = -2.18754807e-8
+ moin = 5.1
+ njtsswg = 9
+ xpart = 1
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ nigc = 3.083
+ pbswgd = 0.95
+ pbswgs = 0.95
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ acnqsmod = 0
+ egidl = 0.29734
+ igcmod = 1
+ ckappad = 0.6
+ ckappas = 0.6
+ noff = 2.7195
+ pdiblc1 = 0
+ pdiblc2 = -0.0010804963
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ pdiblcb = -0.3
+ rbodymod = 0
+ ntox = -0.31099999999999994
+ pcit = -2.7955777e-17
+ pclm = 1.0542662
+ ags = 4.199629600000001
+ bigbacc = 0.002588
+ phin = 0.15
+ cjd = 0.00145199
+ cit = -0.0053953827
+ cjs = 0.00145199
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 3.26497e-9
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ pkt1 = -9.0863924e-16
+ pkt2 = -5.454643e-16
+ dwg = 0
+ dwj = 0
+ kvth0we = 0.00018
+ wpdiblc2 = 2.3632766e-9
+ permod = 1
+ pvoff = 2.2093735000000008e-16
+ lintnoi = -1.5e-8
+ la0 = -1.0940063e-6
+ cdscb = 0
+ cdscd = 0
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.0019085555799999996
+ bigbinv = 0.004953
+ kt1 = -0.47965441
+ kt2 = -0.26453031
+ lk2 = -3.0631458e-10
+ vtsswgd = 4.2
+ pvsat = 8.149221800000001e-10
+ vtsswgs = 4.2
+ llc = 0
+ lln = 1
+ lu0 = 3.3935358e-10
+ wk2we = 5e-12
+ pvth0 = 5.91897254e-16
+ mjd = 0.26
+ mjs = 0.26
+ lua = 3.3186753e-17
+ lub = -3.0003129999999985e-27
+ luc = 7.435334e-18
+ lud = 0
+ rbdb = 50
+ pua1 = 6.1201017e-24
+ prwb = 0
+ lwc = 0
+ pub1 = -1.50107919e-32
+ prwg = 0
+ drout = 0.56
+ lwl = 0
+ puc1 = -2.1235877e-24
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 1.2471671e-13
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ nsd = 1e+20
+ pvag = 1.2
+ pbd = 0.52
+ pat = 6.070153999999999e-11
+ pbs = 0.52
+ pk2 = 1.8168527e-16
+ paigc = -1.0299571e-18
+ pu0 = -1.3197203999999988e-18
+ prt = 0
+ pua = 6.5377716e-24
+ pub = -1.101976303e-32
+ rdsw = 100
+ puc = -3.076481e-25
+ pud = 0
+ voffl = 0
+ rsh = 17.5
+ tcj = 0.00076
+ voffcv = -0.16942
+ wpemod = 1
+ ua1 = 1.4780468e-9
+ ub1 = -2.7008499e-18
+ uc1 = 1.2217521e-10
+ tpb = 0.0014
+ wa0 = -2.130866e-6
+ weta0 = -1.5669611e-7
+ ute = -1
+ wetab = 4.0317659e-8
+ wat = 0.0042150943
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 1.5715655e-9
+ wlc = 0
+ wln = 1
+ wu0 = -2.19928297e-10
+ lpclm = 6.3904735e-9
+ xgl = -1.09e-8
+ wkvth0we = 2e-12
+ xgw = 0
+ wua = -1.3239536e-16
+ wub = 1.9940967600000001e-25
+ wuc = 1.2105201e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ cgidl = 0.22
+ trnqsmod = 0
+ rshg = 15.6
+ wtvfbsdoff = 0
+ nfactor = 1
+ pbswd = 0.8
+ pbsws = 0.8
+ tpbswg = 0.0009
+ ltvfbsdoff = 0
+ rgatemod = 0
+ tnjtsswg = 1
+ pdits = 0
+ tnom = 25
+ cigsd = 0.069865
+ toxe = 2.47e-9
+ ptvoff = -1.0763348e-17
+ toxm = 2.43e-9
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ waigsd = 3.1788545e-12
+ nigbacc = 10
+ pk2we = -1e-19
+ diomod = 1
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ ptvfbsdoff = 0
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 3.0174000000000004e-10
+ pku0we = -1.5e-18
+ cjswgs = 3.0174000000000004e-10
+ wags = -2.3277778e-7
+ tnoia = 0
+ nigbinv = 10
+ wcit = 4.3324313999999997e-10
+ peta0 = 7.5477876e-15
+ petab = -1.7674893e-15
+ voff = -0.056267378999999965
+ wketa = -1.20381479e-7
+ acde = 0.4
+ tvfbsdoff = 0.022
+ tpbsw = 0.0019
+ mjswgd = 0.85
+ mjswgs = 0.85
+ vsat = 153104.713
+ wint = 0
+ cjswd = 8.774000000000001e-11
+ cjsws = 8.774000000000001e-11
+ vth0 = 0.284464339
+ tcjswg = 0.001
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ )

.model nch_ss_40 nmos (
+ level = 54
+ wkt1 = -2.5038067e-8
+ wkt2 = -1.1473225e-8
+ wmax = 2.726e-7
+ aigc = 0.011144932
+ wmin = 1.08e-7
+ fnoimod = 1
+ eigbinv = 1.1
+ wua1 = 1.9140234e-16
+ wub1 = -2.5776439e-25
+ wuc1 = -2.8394855000000005e-17
+ bigc = 0.001442
+ wwlc = 0
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ scref = 1e-6
+ ijthsfwd = 0.01
+ cdsc = 0
+ fprout = 300
+ pigcd = 2.621
+ cgbo = 0
+ aigsd = 0.010772574
+ cgdl = 3.0874977e-12
+ cgdo = 4.5622265999999996e-11
+ xtid = 3
+ xtis = 3
+ xrcrg1 = 12
+ xrcrg2 = 1
+ cgsl = 3.0874977e-12
+ cgso = 4.5622265999999996e-11
+ cigc = 0.000625
+ lvoff = -1.8639393000000007e-9
+ cigbacc = 0.32875
+ lvsat = 0.00614940452
+ wtvoff = -7.2128996e-10
+ lvth0 = 2.1645048000000004e-9
+ ijthsrev = 0.01
+ tnoimod = 0
+ delta = 0.007595625
+ laigc = 5.7720314e-12
+ rnoia = 0
+ rnoib = 0
+ cigbinv = 0.006
+ dmcg = 3.1e-8
+ capmod = 2
+ dmci = 3.1e-8
+ dmdg = 0
+ wku0we = 2e-11
+ pketa = -8.4677334e-15
+ ngate = 8e+20
+ a0 = -5.925916599999999
+ a1 = 0
+ a2 = 1
+ ngcon = 1
+ b0 = 0
+ b1 = 0
+ mobmod = 0
+ wpclm = -7.2101286e-7
+ at = 144965.742
+ cf = 7.5795e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.017523130999999997
+ k3 = -1.8419
+ em = 1000000.0
+ k2we = 5e-5
+ ll = 0
+ lw = 0
+ u0 = 0.012982557999999998
+ w0 = 0
+ ua = -5.589164400000002e-10
+ ub = 8.937269600000036e-20
+ uc = 3.9457239999999995e-10
+ ud = 0
+ version = 4.5
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 5.6700000000000005e-9
+ ww = 0
+ xw = 3.4e-9
+ dsub = 0.75
+ dtox = 2.7e-10
+ gbmin = 1e-12
+ tempmod = 0
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ eta0 = -0.30390379700000003
+ aigbacc = 0.02
+ etab = -0.74723747
+ laigsd = -1.5325105e-17
+ pkvth0we = -1.3e-19
+ aigbinv = 0.0163
+ tvoff = 0.0062987975
+ vfbsdoff = 0.02
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ paramchk = 1
+ ku0we = -0.0007
+ beta0 = 13
+ leta0 = 2.8103219e-8
+ poxedge = 1
+ letab = 2.3120738e-8
+ ppclm = 3.3171145e-14
+ binunit = 2
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ ijthdfwd = 0.01
+ toxref = 3e-9
+ dmcgt = 0
+ keta = -0.51478944
+ tcjsw = 0.000357
+ ijthdrev = 0.01
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 1.741214e-10
+ ltvoff = -2.4217179e-10
+ kt1l = 0
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ bigsd = 0.00125
+ lint = 0
+ wvoff = 1.85924831e-8
+ lkt1 = -1.4940467e-9
+ lkt2 = -1.1864945e-9
+ lmax = 4.333e-8
+ lmin = 3.6e-8
+ wvsat = 0.0259582414
+ lku0we = 2.5e-11
+ pvfbsdoff = 0
+ lpe0 = 9.2e-8
+ wvth0 = -1.4766607e-8
+ lpeb = 2.5e-7
+ epsrox = 3.9
+ waigc = 5.1623453e-11
+ minv = -0.3
+ lua1 = 6.0050187e-18
+ lub1 = 4.0140646999999995e-27
+ luc1 = 5.7838555e-18
+ rdsmod = 0
+ lkvth0we = -2e-12
+ ndep = 1e+18
+ igbmod = 1
+ lwlc = 0
+ lketa = 2.6802806000000003e-8
+ moin = 5.1
+ njtsswg = 9
+ xpart = 1
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ nigc = 3.083
+ pbswgd = 0.95
+ pbswgs = 0.95
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ acnqsmod = 0
+ egidl = 0.29734
+ igcmod = 1
+ ckappad = 0.6
+ ckappas = 0.6
+ noff = 2.7195
+ pdiblc1 = 0
+ pdiblc2 = -0.0010804963
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ pdiblcb = -0.3
+ rbodymod = 0
+ ntox = -0.31099999999999994
+ pcit = -9.987879999999998e-18
+ pclm = 4.6708343
+ ags = 4.199629600000001
+ bigbacc = 0.002588
+ phin = 0.15
+ paigsd = 4.2297301e-24
+ cjd = 0.00145199
+ cit = 0.0010105263
+ cjs = 0.00145199
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 3.26497e-9
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ pkt1 = 6.6911236e-16
+ pkt2 = 5.863609e-16
+ dwg = 0
+ dwj = 0
+ kvth0we = 0.00018
+ wpdiblc2 = 2.3632766e-9
+ permod = 1
+ pvoff = -7.993068399999999e-16
+ lintnoi = -1.5e-8
+ la0 = 1.3676219000000002e-7
+ cdscb = 0
+ cdscd = 0
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.00444752332
+ bigbinv = 0.004953
+ kt1 = -0.23663458
+ kt2 = -0.073003235
+ lk2 = -3.894925700000001e-9
+ vtsswgd = 4.2
+ pvsat = -1.08687436e-9
+ vtsswgs = 4.2
+ llc = 0
+ lln = 1
+ lu0 = -1.3862676e-10
+ wk2we = 5e-12
+ pvth0 = 8.1295839e-16
+ mjd = 0.26
+ mjs = 0.26
+ lua = -5.56054081e-17
+ lub = 6.391826569999999e-26
+ luc = -1.91434719e-17
+ lud = 0
+ rbdb = 50
+ pua1 = -8.5382538e-24
+ prwb = 0
+ lwc = 0
+ pub1 = 1.16183448e-32
+ prwg = 0
+ drout = 0.56
+ lwl = 0
+ puc1 = 3.138452e-25
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = -7.5523402e-14
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ nsd = 1e+20
+ pvag = 1.2
+ pbd = 0.52
+ pat = 5.3899479999999974e-11
+ pbs = 0.52
+ pk2 = 5.0756697e-16
+ paigc = -1.5534524e-18
+ pu0 = -6.852166199999999e-18
+ prt = 0
+ pua = -2.8276596999999977e-25
+ pub = -6.331388000000253e-35
+ rdsw = 100
+ puc = 2.5547617e-24
+ pud = 0
+ voffl = 0
+ rsh = 17.5
+ tcj = 0.00076
+ voffcv = -0.16942
+ wpemod = 1
+ ua1 = 5.4333072e-10
+ ub1 = -1.07203754e-18
+ uc1 = 2.985545e-11
+ tpb = 0.0014
+ wa0 = 1.9556670799999998e-6
+ weta0 = 9.9276847e-8
+ ute = -1
+ wetab = 3.9258957e-9
+ wat = 0.0043539224999999985
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -5.0790816e-9
+ wlc = 0
+ wln = 1
+ wu0 = -1.0702157e-10
+ lpclm = -1.70821362e-7
+ xgl = -1.09e-8
+ wkvth0we = 2e-12
+ xgw = 0
+ wua = 6.799270000000015e-18
+ wub = -2.4191335000000008e-26
+ wuc = -4.6311215e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ cgidl = 0.22
+ trnqsmod = 0
+ rshg = 15.6
+ wtvfbsdoff = 0
+ nfactor = 1
+ pbswd = 0.8
+ pbsws = 0.8
+ tpbswg = 0.0009
+ ltvfbsdoff = 0
+ rgatemod = 0
+ tnjtsswg = 1
+ pdits = 0
+ tnom = 25
+ cigsd = 0.069865
+ toxe = 2.47e-9
+ ptvoff = 2.8458255e-17
+ toxm = 2.43e-9
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ waigsd = 3.1787682e-12
+ nigbacc = 10
+ pk2we = -1e-19
+ diomod = 1
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ ptvfbsdoff = 0
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 3.0174000000000004e-10
+ pku0we = -1.5e-18
+ cjswgs = 3.0174000000000004e-10
+ wags = -2.3277778e-7
+ tnoia = 0
+ nigbinv = 10
+ wcit = 6.655421999999997e-11
+ peta0 = -4.9948868e-15
+ petab = 1.5707054e-17
+ voff = -0.150644936
+ wketa = 1.65035329e-7
+ acde = 0.4
+ tvfbsdoff = 0.022
+ tpbsw = 0.0019
+ mjswgd = 0.85
+ mjswgs = 0.85
+ vsat = -32538.627999999982
+ wint = 0
+ cjswd = 8.774000000000001e-11
+ cjsws = 8.774000000000001e-11
+ vth0 = 0.369989347
+ tcjswg = 0.001
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ )

.model nch_tt_1 nmos (
+ level = 54
+ fprout = 300
+ xrcrg1 = 12
+ xrcrg2 = 1
+ ags = 0.8675
+ wtvoff = 0
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ tvoff = 0.0019109629
+ keta = -0.06
+ cjd = 0.001357
+ cit = 0.0001
+ cjs = 0.001357
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 9.8024918e-9
+ xjbvd = 1
+ k3b = 1.9326
+ xjbvs = 1
+ lk2we = -1.5e-12
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ tvfbsdoff = 0.022
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 0
+ capmod = 2
+ la0 = 0
+ kt1l = 0
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = 0
+ kt1 = -0.200226
+ kt2 = -0.05325
+ wku0we = 2e-11
+ wkvth0we = 2e-12
+ llc = 0
+ ku0we = -0.0007
+ lln = 1
+ lu0 = 0
+ mjd = 0.26
+ mjs = 0.26
+ beta0 = 13
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ leta0 = 0
+ njs = 1.02
+ pa0 = 0
+ mobmod = 0
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 0
+ pbs = 0.52
+ lint = 6.5375218e-9
+ trnqsmod = 0
+ pu0 = 0
+ prt = 0
+ pud = 0
+ lkt1 = 0
+ lmax = 2.001e-5
+ lmin = 8.9991e-6
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 1.2299687e-9
+ ub1 = -7.2455506e-19
+ uc1 = 3.028e-11
+ dlcig = 2.5e-9
+ tpb = 0.0014
+ lpe0 = 9.2e-8
+ njtsswg = 9
+ bgidl = 2320000000.0
+ lpeb = 2.5e-7
+ wa0 = 0
+ ute = -1.007
+ wat = 0
+ web = 6843.8
+ wec = -25529.0
+ wlc = 0
+ wln = 1
+ wu0 = 0
+ xgl = -1.09e-8
+ xgw = 0
+ wud = 0
+ wwc = 0
+ minv = -0.3
+ wwl = 0
+ wwn = 1
+ xtsswgd = 0.18
+ wvfbsdoff = 0
+ xtsswgs = 0.18
+ lvfbsdoff = 0
+ lub1 = 0
+ ndep = 1e+18
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.018555248
+ lwlc = 0
+ rgatemod = 0
+ dmcgt = 0
+ pdiblcb = -0.3
+ moin = 5.1
+ tcjsw = 0.000357
+ tnjtsswg = 1
+ nigc = 3.083
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ bigsd = 0.00125
+ bigbacc = 0.002588
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ wvoff = 0
+ ntox = 1
+ pcit = 0
+ kvth0we = 0.00018
+ pclm = 1.4
+ wvsat = 0
+ wvth0 = 0
+ lintnoi = -1.5e-8
+ bigbinv = 0.004953
+ phin = 0.15
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ pkt1 = 0
+ a0 = 3.25
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 72000
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.024601254
+ k3 = -1.8419
+ em = 1000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.01567
+ w0 = 0
+ ua = -1.8237726e-9
+ ub = 2.103696e-18
+ xpart = 1
+ uc = 7.33e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 6e-9
+ toxref = 3e-9
+ rbdb = 50
+ prwb = 0
+ prwg = 0
+ pub1 = 0
+ egidl = 0.29734
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ rdsw = 100
+ ijthsfwd = 0.01
+ ltvoff = 0
+ nfactor = 1
+ rshg = 15.6
+ ijthsrev = 0.01
+ pvoff = 0
+ lku0we = 2.5e-11
+ cdscb = 0
+ cdscd = 0
+ epsrox = 3.9
+ pvsat = 0
+ wk2we = 5e-12
+ pvth0 = 0
+ drout = 0.56
+ nigbacc = 10
+ rdsmod = 0
+ igbmod = 1
+ voffl = 0
+ tnom = 25
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ weta0 = 0
+ pbswgd = 0.95
+ pbswgs = 0.95
+ nigbinv = 10
+ igcmod = 1
+ cgidl = 0.22
+ wags = 0
+ wcit = 0
+ voff = -0.1128204
+ fnoimod = 1
+ pbswd = 0.8
+ pbsws = 0.8
+ acde = 0.4
+ pkvth0we = -1.3e-19
+ eigbinv = 1.1
+ vsat = 102860
+ wint = 0
+ vth0 = 0.34911089
+ wkt1 = 0
+ pvfbsdoff = 0
+ wmax = 0.00090001
+ aigc = 0.011769394
+ wmin = 9e-6
+ pdits = 0
+ vfbsdoff = 0.02
+ permod = 1
+ cigsd = 0.069865
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ bigc = 0.001442
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ paramchk = 1
+ wwlc = 0
+ cigbacc = 0.32875
+ voffcv = -0.16942
+ wpemod = 1
+ cdsc = 0
+ tnoia = 0
+ tnoimod = 0
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ peta0 = 0
+ cigbinv = 0.006
+ tpbsw = 0.0019
+ ijthdfwd = 0.01
+ cjswd = 8.2e-11
+ cjsws = 8.2e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ version = 4.5
+ tempmod = 0
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ tpbswg = 0.0009
+ ijthdrev = 0.01
+ aigbacc = 0.02
+ k2we = 5e-5
+ dsub = 0.75
+ dtox = 2.7e-10
+ scref = 1e-6
+ ptvoff = 0
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ pigcd = 2.621
+ aigsd = 0.01077322
+ lvoff = 0
+ eta0 = 0.3
+ aigbinv = 0.0163
+ diomod = 1
+ etab = -0.25
+ wtvfbsdoff = 0
+ lvsat = 0
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 2.82e-10
+ pku0we = -1.5e-18
+ lvth0 = 0
+ cjswgs = 2.82e-10
+ lkvth0we = -2e-12
+ delta = 0.007595625
+ ltvfbsdoff = 0
+ rnoia = 0
+ rnoib = 0
+ mjswgd = 0.85
+ mjswgs = 0.85
+ acnqsmod = 0
+ ngate = 8e+20
+ tcjswg = 0.001
+ ngcon = 1
+ poxedge = 1
+ rbodymod = 0
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ binunit = 2
+ ptvfbsdoff = 0
+ )

.model nch_tt_2 nmos (
+ level = 54
+ wtvoff = 0
+ cgidl = 0.22
+ ijthdfwd = 0.01
+ capmod = 2
+ pbswd = 0.8
+ pbsws = 0.8
+ wku0we = 2e-11
+ rshg = 15.6
+ cigbacc = 0.32875
+ mobmod = 0
+ pvfbsdoff = 0
+ ijthdrev = 0.01
+ tnoimod = 0
+ pdits = 0
+ lpdiblc2 = -5.8501673e-10
+ cigsd = 0.069865
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ cigbinv = 0.006
+ tnom = 25
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ version = 4.5
+ tnoia = 0
+ tempmod = 0
+ lkvth0we = -2e-12
+ peta0 = 0
+ tpbsw = 0.0019
+ aigbacc = 0.02
+ wags = 0
+ cjswd = 8.2e-11
+ cjsws = 8.2e-11
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ wcit = 0
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ acnqsmod = 0
+ voff = -0.11120139
+ acde = 0.4
+ vsat = 102860
+ wint = 0
+ rbodymod = 0
+ aigbinv = 0.0163
+ vth0 = 0.34336703
+ wkt1 = 0
+ wmax = 0.00090001
+ aigc = 0.01178613
+ wmin = 9e-6
+ scref = 1e-6
+ pigcd = 2.621
+ toxref = 3e-9
+ aigsd = 0.01077322
+ bigc = 0.001442
+ wwlc = 0
+ lvoff = -1.4554874e-8
+ poxedge = 1
+ cdsc = 0
+ lvsat = 0
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ lvth0 = 5.1637332e-8
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ delta = 0.007595625
+ binunit = 2
+ laigc = -1.5044982e-10
+ rnoia = 0
+ rnoib = 0
+ ltvoff = -1.4627394e-10
+ a0 = 3.4752469
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ ngate = 8e+20
+ at = 61592.494
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.026088843
+ k3 = -1.8419
+ em = 1000000.0
+ ngcon = 1
+ ll = 0
+ lw = 0
+ u0 = 0.015891951
+ w0 = 0
+ ua = -1.7995884e-9
+ ub = 2.1046515e-18
+ uc = 7.3387901e-11
+ ud = 0
+ wkvth0we = 2e-12
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 6e-9
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ lku0we = 2.5e-11
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ trnqsmod = 0
+ epsrox = 3.9
+ k2we = 5e-5
+ rdsmod = 0
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ dsub = 0.75
+ dtox = 2.7e-10
+ igbmod = 1
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ ags = 0.87104901
+ pbswgd = 0.95
+ pbswgs = 0.95
+ eta0 = 0.3
+ cjd = 0.001357
+ rgatemod = 0
+ etab = -0.25
+ cit = -2.3830864e-5
+ cjs = 0.001357
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 9.8024918e-9
+ tnjtsswg = 1
+ k3b = 1.9326
+ igcmod = 1
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ tvoff = 0.0019272336
+ la0 = -2.0249698e-6
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = 0.093563481
+ kt1 = -0.19577666
+ lk2 = -1.337342e-8
+ kt2 = -0.051823539
+ xjbvd = 1
+ llc = 0
+ xjbvs = 1
+ lln = 1
+ tvfbsdoff = 0.022
+ lk2we = -1.5e-12
+ lu0 = -1.9953361e-9
+ mjd = 0.26
+ lua = -2.1741579e-16
+ mjs = 0.26
+ lub = -8.5898229e-27
+ luc = -7.902321e-19
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njtsswg = 9
+ njd = 1.02
+ njs = 1.02
+ pa0 = 0
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 0
+ pbs = 0.52
+ pu0 = 0
+ xtsswgd = 0.18
+ prt = 0
+ pud = 0
+ xtsswgs = 0.18
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 1.2713861e-9
+ ub1 = -7.4616446e-19
+ ku0we = -0.0007
+ uc1 = 2.5703642e-11
+ ckappad = 0.6
+ ckappas = 0.6
+ beta0 = 13
+ tpb = 0.0014
+ wa0 = 0
+ leta0 = 0
+ pdiblc1 = 0
+ pdiblc2 = 0.018620322
+ pdiblcb = -0.3
+ ute = -1.0077691
+ wat = 0
+ web = 6843.8
+ wec = -25529.0
+ wlc = 0
+ wln = 1
+ wu0 = 0
+ xgl = -1.09e-8
+ xgw = 0
+ permod = 1
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ bigbacc = 0.002588
+ voffcv = -0.16942
+ wpemod = 1
+ dmcgt = 0
+ tcjsw = 0.000357
+ kvth0we = 0.00018
+ lintnoi = -1.5e-8
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ keta = -0.059896633
+ ijthsfwd = 0.01
+ bigsd = 0.00125
+ lags = -3.1905621e-8
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 1.1132395e-9
+ wvoff = 0
+ kt1l = 0
+ tpbswg = 0.0009
+ wvsat = 0
+ wvth0 = 0
+ ijthsrev = 0.01
+ lint = 6.5375218e-9
+ lkt1 = -3.9999573e-8
+ lkt2 = -1.2823887e-8
+ wtvfbsdoff = 0
+ lmax = 8.9991e-6
+ lmin = 8.9908e-7
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ ptvoff = 0
+ lketa = -9.2926692e-10
+ xpart = 1
+ ltvfbsdoff = 0
+ minv = -0.3
+ lua1 = -3.7234224e-16
+ lub1 = 1.9426851e-25
+ luc1 = 4.1141459e-17
+ nfactor = 1
+ diomod = 1
+ ndep = 1e+18
+ lute = 6.9145309e-9
+ egidl = 0.29734
+ lwlc = 0
+ moin = 5.1
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 2.82e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.82e-10
+ nigc = 3.083
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ mjswgd = 0.85
+ mjswgs = 0.85
+ nigbacc = 10
+ ptvfbsdoff = 0
+ tcjswg = 0.001
+ ntox = 1
+ pkvth0we = -1.3e-19
+ pcit = 0
+ pclm = 1.4
+ pvoff = 0
+ nigbinv = 10
+ phin = 0.15
+ cdscb = 0
+ cdscd = 0
+ vfbsdoff = 0.02
+ pvsat = 0
+ wk2we = 5e-12
+ pkt1 = 0
+ pvth0 = 0
+ drout = 0.56
+ voffl = 0
+ fprout = 300
+ paramchk = 1
+ rbdb = 50
+ prwb = 0
+ prwg = 0
+ pub1 = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ fnoimod = 1
+ weta0 = 0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ eigbinv = 1.1
+ rdsw = 100
+ )

.model nch_tt_3 nmos (
+ level = 54
+ ku0we = -0.0007
+ beta0 = 13
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ leta0 = 0
+ ijthsrev = 0.01
+ kvth0we = 0.00018
+ lintnoi = -1.5e-8
+ k2we = 5e-5
+ bigbinv = 0.004953
+ dlcig = 2.5e-9
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ bgidl = 2320000000.0
+ dsub = 0.75
+ wvfbsdoff = 0
+ dtox = 2.7e-10
+ lvfbsdoff = 0
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ eta0 = 0.3
+ dmcgt = 0
+ etab = -0.25
+ tcjsw = 0.000357
+ bigsd = 0.00125
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ wvoff = 0
+ pkvth0we = -1.3e-19
+ nfactor = 1
+ wvsat = 0
+ wvth0 = 0
+ vfbsdoff = 0.02
+ lketa = -2.6515603e-8
+ toxref = 3e-9
+ xpart = 1
+ nigbacc = 10
+ paramchk = 1
+ egidl = 0.29734
+ nigbinv = 10
+ keta = -0.031147941
+ ltvoff = -6.4393769e-10
+ ijthdfwd = 0.01
+ lags = 4.0889306e-7
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = -1.1051822e-10
+ kt1l = 0
+ lku0we = 2.5e-11
+ fnoimod = 1
+ ijthdrev = 0.01
+ epsrox = 3.9
+ eigbinv = 1.1
+ pvoff = 0
+ lint = 6.5375218e-9
+ cdscb = 0
+ cdscd = 0
+ lkt1 = -1.7764368e-8
+ lkt2 = -1.1493547e-8
+ lmax = 8.9908e-7
+ lpdiblc2 = 3.0380287e-9
+ pvsat = 0
+ lmin = 4.4908e-7
+ rdsmod = 0
+ wk2we = 5e-12
+ pvth0 = 0
+ drout = 0.56
+ igbmod = 1
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ minv = -0.3
+ voffl = 0
+ lua1 = -1.0281867e-16
+ lub1 = 1.8552992e-26
+ luc1 = 3.7680622e-18
+ pbswgd = 0.95
+ pbswgs = 0.95
+ ndep = 1e+18
+ weta0 = 0
+ lwlc = 0
+ igcmod = 1
+ moin = 5.1
+ a0 = 1.288
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ cigbacc = 0.32875
+ at = 219598.22
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.025010322
+ k3 = -1.8419
+ em = 1000000.0
+ ll = 0
+ nigc = 3.083
+ lw = 0
+ u0 = 0.015390444
+ w0 = 0
+ ua = -1.9429424e-9
+ ub = 2.1566e-18
+ uc = 9.3717778e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 6e-9
+ lkvth0we = -2e-12
+ cgidl = 0.22
+ tnoimod = 0
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ cigbinv = 0.006
+ acnqsmod = 0
+ pbswd = 0.8
+ pbsws = 0.8
+ ntox = 1
+ pcit = 0
+ pclm = 1.4
+ pvfbsdoff = 0
+ rbodymod = 0
+ version = 4.5
+ permod = 1
+ phin = 0.15
+ tempmod = 0
+ pdits = 0
+ cigsd = 0.069865
+ pkt1 = 0
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ aigbacc = 0.02
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ voffcv = -0.16942
+ wpemod = 1
+ rbdb = 50
+ prwb = 0
+ pub1 = 0
+ prwg = 0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ tnoia = 0
+ rdsw = 100
+ aigbinv = 0.0163
+ peta0 = 0
+ tpbsw = 0.0019
+ wtvfbsdoff = 0
+ cjswd = 8.2e-11
+ cjsws = 8.2e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ tpbswg = 0.0009
+ rshg = 15.6
+ ltvfbsdoff = 0
+ wkvth0we = 2e-12
+ poxedge = 1
+ trnqsmod = 0
+ ptvoff = 0
+ binunit = 2
+ scref = 1e-6
+ pigcd = 2.621
+ aigsd = 0.01077322
+ tnom = 25
+ diomod = 1
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ ptvfbsdoff = 0
+ lvoff = -1.3768912e-8
+ pditsd = 0
+ rgatemod = 0
+ pditsl = 0
+ cjswgd = 2.82e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.82e-10
+ tnjtsswg = 1
+ lvsat = 0
+ lvth0 = 7.4115504e-9
+ delta = 0.007595625
+ laigc = -5.5724245e-11
+ rnoia = 0
+ rnoib = 0
+ mjswgd = 0.85
+ mjswgs = 0.85
+ wags = 0
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ wcit = 0
+ tcjswg = 0.001
+ ngate = 8e+20
+ voff = -0.1120845
+ acde = 0.4
+ ngcon = 1
+ vsat = 102860
+ wint = 0
+ vth0 = 0.39305892
+ gbmin = 1e-12
+ wkt1 = 0
+ jswgd = 1.28e-13
+ wmax = 0.00090001
+ jswgs = 1.28e-13
+ aigc = 0.011679696
+ wmin = 9e-6
+ ags = 0.3757696
+ cjd = 0.001357
+ cit = 0.0013511778
+ cjs = 0.001357
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 9.8024918e-9
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ fprout = 300
+ dwg = 0
+ dwj = 0
+ njtsswg = 9
+ bigc = 0.001442
+ xrcrg1 = 12
+ xrcrg2 = 1
+ wwlc = 0
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ la0 = -7.832e-8
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.047061618
+ kt1 = -0.22076004
+ kt2 = -0.053318302
+ lk2 = -1.2413537e-8
+ llc = 0
+ cdsc = 0
+ lln = 1
+ lu0 = -1.5489956e-9
+ ckappad = 0.6
+ ckappas = 0.6
+ mjd = 0.26
+ mjs = 0.26
+ lua = -8.9830708e-17
+ lub = -5.4824e-26
+ luc = -1.8883822e-17
+ lud = 0
+ lwc = 0
+ cgbo = 0
+ wtvoff = 0
+ lwl = 0
+ lwn = 1
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ pdiblc1 = 0
+ pdiblc2 = 0.014549485
+ njd = 1.02
+ xtis = 3
+ njs = 1.02
+ pa0 = 0
+ pdiblcb = -0.3
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 0
+ pbs = 0.52
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ pu0 = 0
+ tvoff = 0.0024864064
+ prt = 0
+ pud = 0
+ tvfbsdoff = 0.022
+ rsh = 17.5
+ tcj = 0.00076
+ ijthsfwd = 0.01
+ xjbvd = 1
+ ua1 = 9.685506e-10
+ ub1 = -5.4873129e-19
+ xjbvs = 1
+ uc1 = 6.7696222e-11
+ lk2we = -1.5e-12
+ tpb = 0.0014
+ capmod = 2
+ wa0 = 0
+ ute = -1
+ wat = 0
+ web = 6843.8
+ wec = -25529.0
+ wlc = 0
+ wln = 1
+ wku0we = 2e-11
+ wu0 = 0
+ xgl = -1.09e-8
+ xgw = 0
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ bigbacc = 0.002588
+ mobmod = 0
+ )

.model nch_tt_4 nmos (
+ level = 54
+ minv = -0.3
+ lua1 = -3.0475764e-17
+ pk2we = -1e-19
+ lub1 = -2.9971927e-26
+ luc1 = -4.3987511e-18
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ ndep = 1e+18
+ rgatemod = 0
+ lwlc = 0
+ moin = 5.1
+ tnjtsswg = 1
+ tnoia = 0
+ nigc = 3.083
+ peta0 = 0
+ poxedge = 1
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ tpbsw = 0.0019
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ binunit = 2
+ cjswd = 8.2e-11
+ cjsws = 8.2e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ ntox = 1
+ pcit = 0
+ pclm = 1.5439223
+ phin = 0.15
+ pkt1 = 0
+ toxref = 3e-9
+ scref = 1e-6
+ jtsswgd = 2.3e-7
+ pigcd = 2.621
+ jtsswgs = 2.3e-7
+ aigsd = 0.01077322
+ rbdb = 50
+ prwb = 0
+ pub1 = 0
+ prwg = 0
+ lvoff = -6.3216134e-9
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ rdsw = 100
+ lvsat = 0
+ lvth0 = -4.690878e-9
+ delta = 0.007595625
+ ltvoff = -1.206053e-10
+ laigc = -1.9935708e-11
+ rnoia = 0
+ rnoib = 0
+ ijthsfwd = 0.01
+ ngate = 8e+20
+ njtsswg = 9
+ ngcon = 1
+ rshg = 15.6
+ lku0we = 2.5e-11
+ ags = 0.054315598
+ epsrox = 3.9
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ cjd = 0.001357
+ cit = 0.00073144105
+ ijthsrev = 0.01
+ cjs = 0.001357
+ clc = 1e-7
+ cle = 0.6
+ gbmin = 1e-12
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 1.30529375e-8
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ k3b = 1.9326
+ ckappad = 0.6
+ ckappas = 0.6
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ rdsmod = 0
+ pdiblc1 = 0
+ pdiblc2 = 0.027331777
+ pdiblcb = -0.3
+ igbmod = 1
+ la0 = -2.4730306e-7
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.016865258
+ kt1 = -0.23920434
+ kt2 = -0.070668297
+ lk2 = -9.6174482e-9
+ llc = -1.18e-13
+ lln = 0.7
+ lu0 = -6.2433887e-10
+ mjd = 0.26
+ mjs = 0.26
+ lua = -1.0757894e-17
+ lub = -4.7838952e-26
+ luc = -6.6488035e-18
+ lud = 0
+ pbswgd = 0.95
+ pbswgs = 0.95
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ tnom = 25
+ njd = 1.02
+ njs = 1.02
+ pa0 = 0
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 0
+ pbs = 0.52
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ pu0 = 0
+ igcmod = 1
+ prt = 0
+ pud = 0
+ bigbacc = 0.002588
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 8.041349e-10
+ ub1 = -4.3844738e-19
+ uc1 = 8.6257162e-11
+ tpb = 0.0014
+ wa0 = 0
+ ute = -1
+ wat = 0
+ web = 6843.8
+ wec = -25529.0
+ kvth0we = 0.00018
+ wlc = 0
+ wln = 1
+ wu0 = 0
+ xgl = -1.09e-8
+ xgw = 0
+ tvoff = 0.0012970146
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ tvfbsdoff = 0.022
+ lintnoi = -1.5e-8
+ xjbvd = 1
+ xjbvs = 1
+ wags = 0
+ lk2we = -1.5e-12
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ wcit = 0
+ voff = -0.12901018
+ acde = 0.4
+ pkvth0we = -1.3e-19
+ ku0we = -0.0007
+ beta0 = 13
+ vsat = 102860
+ wint = 0
+ permod = 1
+ leta0 = 0
+ vth0 = 0.42056443
+ wkt1 = 0
+ wmax = 0.00090001
+ aigc = 0.011598359
+ wmin = 9e-6
+ vfbsdoff = 0.02
+ a0 = 1.6720524
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 150970.13
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.018655575
+ k3 = -1.8419
+ em = 1000000.0
+ dlcig = 2.5e-9
+ ll = -1.18e-13
+ wvfbsdoff = 0
+ lw = 0
+ u0 = 0.013288952
+ bgidl = 2320000000.0
+ w0 = 0
+ lvfbsdoff = 0
+ ua = -2.1226533e-9
+ ub = 2.1407249e-18
+ uc = 6.5910917e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 6e-9
+ voffcv = -0.16942
+ wpemod = 1
+ bigc = 0.001442
+ paramchk = 1
+ wwlc = 0
+ wtvfbsdoff = 0
+ dmcgt = 0
+ tcjsw = 0.000357
+ nfactor = 1
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ ltvfbsdoff = 0
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ ijthdfwd = 0.01
+ bigsd = 0.00125
+ tpbswg = 0.0009
+ wvoff = 0
+ nigbacc = 10
+ wvsat = 0
+ wvth0 = 0
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ ijthdrev = 0.01
+ ptvfbsdoff = 0
+ lpdiblc2 = -2.58618e-9
+ ptvoff = 0
+ nigbinv = 10
+ k2we = 5e-5
+ dsub = 0.75
+ lketa = -2.2644187e-8
+ dtox = 2.7e-10
+ xpart = 1
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ diomod = 1
+ pditsd = 0
+ pditsl = 0
+ egidl = 0.29734
+ cjswgd = 2.82e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.82e-10
+ eta0 = 0.3
+ etab = -0.25
+ fnoimod = 1
+ eigbinv = 1.1
+ lkvth0we = -2e-12
+ mjswgd = 0.85
+ mjswgs = 0.85
+ tcjswg = 0.001
+ acnqsmod = 0
+ rbodymod = 0
+ pvoff = 0
+ cigbacc = 0.32875
+ cdscb = 0
+ cdscd = 0
+ pvsat = 0
+ wk2we = 5e-12
+ pvth0 = 0
+ drout = 0.56
+ tnoimod = 0
+ fprout = 300
+ voffl = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ cigbinv = 0.006
+ weta0 = 0
+ lpclm = -6.3325799e-8
+ wtvoff = 0
+ version = 4.5
+ cgidl = 0.22
+ tempmod = 0
+ keta = -0.039946614
+ capmod = 2
+ lags = 5.5033282e-7
+ wku0we = 2e-11
+ aigbacc = 0.02
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 1.6216594e-10
+ pbswd = 0.8
+ mobmod = 0
+ pbsws = 0.8
+ kt1l = 0
+ wkvth0we = 2e-12
+ pvfbsdoff = 0
+ lint = 9.7879675e-9
+ trnqsmod = 0
+ pdits = 0
+ lkt1 = -9.6488734e-9
+ lkt2 = -3.8595493e-9
+ aigbinv = 0.0163
+ lmax = 4.4908e-7
+ cigsd = 0.069865
+ lmin = 2.1577e-7
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ laigsd = -8.1082969e-17
+ )

.model nch_tt_5 nmos (
+ level = 54
+ nigbinv = 10
+ bigsd = 0.00125
+ wags = 0
+ wcit = 0
+ acnqsmod = 0
+ wvoff = 0
+ voff = -0.15746310460000001
+ acde = 0.4
+ wvsat = 0
+ vsat = 102521.2852
+ wvth0 = 0
+ rbodymod = 0
+ wint = 0
+ vth0 = 0.4365613742
+ wkt1 = 0
+ wmax = 0.00090001
+ aigc = 0.011526753
+ wmin = 9e-6
+ fnoimod = 1
+ eigbinv = 1.1
+ toxref = 3e-9
+ lketa = -1.1430034e-8
+ xpart = 1
+ bigc = 0.001442
+ wwlc = 0
+ egidl = 0.29734
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ ltvoff = 1.4850105e-11
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ cigbacc = 0.32875
+ tnoimod = 0
+ lku0we = 2.5e-11
+ cigbinv = 0.006
+ epsrox = 3.9
+ wkvth0we = 2e-12
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ pvoff = 0
+ rdsmod = 0
+ trnqsmod = 0
+ cdscb = 0
+ cdscd = 0
+ igbmod = 1
+ pvsat = 0
+ version = 4.5
+ wk2we = 5e-12
+ pvth0 = 0
+ k2we = 5e-5
+ drout = 0.56
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ tempmod = 0
+ dsub = 0.75
+ dtox = 2.7e-10
+ pbswgd = 0.95
+ pbswgs = 0.95
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ voffl = 0
+ igcmod = 1
+ aigbacc = 0.02
+ weta0 = 0
+ eta0 = 0.3
+ rgatemod = 0
+ etab = -0.25
+ lpclm = -2.4377173e-8
+ tnjtsswg = 1
+ cgidl = 0.22
+ aigbinv = 0.0163
+ pbswd = 0.8
+ pbsws = 0.8
+ pvfbsdoff = 0
+ permod = 1
+ wtvfbsdoff = 0
+ pdits = 0
+ cigsd = 0.069865
+ dvt0w = 0
+ dvt1w = 0
+ poxedge = 1
+ dvt2w = 0
+ ltvfbsdoff = 0
+ voffcv = -0.16942
+ wpemod = 1
+ binunit = 2
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ tnoia = 0
+ peta0 = 0
+ wketa = 0
+ keta = -0.093093889
+ ptvfbsdoff = 0
+ tpbsw = 0.0019
+ ijthsfwd = 0.01
+ cjswd = 8.2e-11
+ cjsws = 8.2e-11
+ a0 = 0.66068814
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ mjswd = 0.11
+ lags = 3.3904274e-13
+ mjsws = 0.11
+ agidl = 9.41e-8
+ tpbswg = 0.0009
+ at = 79499.116
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = -0.016112078
+ k3 = -1.8419
+ em = 1000000.0
+ jswd = 1.28e-13
+ ll = -1.18e-13
+ jsws = 1.28e-13
+ lw = 0
+ u0 = 0.011286872
+ w0 = 0
+ lcit = 8.4591162e-11
+ ua = -2.2893587e-9
+ ub = 2.089788886e-18
+ uc = 4.5969231e-11
+ ud = 0
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 6e-9
+ kt1l = 0
+ ijthsrev = 0.01
+ lint = 9.7879675e-9
+ ptvoff = 0
+ lkt1 = -3.3075226e-9
+ lkt2 = -6.0180086e-10
+ lmax = 2.1577e-7
+ lmin = 9e-8
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ scref = 1e-6
+ diomod = 1
+ pigcd = 2.621
+ minv = -0.3
+ aigsd = 0.01077322
+ lua1 = 7.6861327e-18
+ lub1 = -5.2342256e-26
+ luc1 = -4.2210821e-18
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 2.82e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.82e-10
+ ndep = 1e+18
+ lvoff = -3.1806260000000004e-10
+ njtsswg = 9
+ lwlc = 0
+ moin = 5.1
+ lvsat = 7.148430000000002e-5
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ lvth0 = -8.0662159e-9
+ nigc = 3.083
+ delta = 0.007595625
+ mjswgd = 0.85
+ mjswgs = 0.85
+ laigc = -4.8268328e-12
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.02163037
+ pdiblcb = -0.3
+ tcjswg = 0.001
+ rnoia = 0
+ rnoib = 0
+ ags = 2.6625264
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ cjd = 0.001357
+ cit = 0.001099094
+ cjs = 0.001357
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 1.30529375e-8
+ pketa = 0
+ ngate = 8e+20
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ ngcon = 1
+ pkvth0we = -1.3e-19
+ ntox = 1
+ pcit = 0
+ pclm = 1.3593316
+ bigbacc = 0.002588
+ la0 = -3.3904685e-8
+ gbmin = 1e-12
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.0017848735
+ kt1 = -0.26925814
+ kt2 = -0.086107863
+ lk2 = -2.2814734e-9
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ llc = -1.18e-13
+ lln = 0.7
+ phin = 0.15
+ lu0 = -2.0189995e-10
+ mjd = 0.26
+ mjs = 0.26
+ lua = 2.4416942e-17
+ lub = -3.7091512499999996e-26
+ luc = -2.4411077e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ vfbsdoff = 0.02
+ njd = 1.02
+ njs = 1.02
+ pa0 = 0
+ nsd = 1e+20
+ kvth0we = 0.00018
+ pbd = 0.52
+ pat = 0
+ pbs = 0.52
+ pkt1 = 0
+ pu0 = 0
+ prt = 0
+ fprout = 300
+ pub = 0
+ pud = 0
+ lintnoi = -1.5e-8
+ rsh = 17.5
+ xrcrg1 = 12
+ xrcrg2 = 1
+ tcj = 0.00076
+ ua1 = 6.2327283e-10
+ ub1 = -3.3242687e-19
+ uc1 = 8.5415128e-11
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ tpb = 0.0014
+ wa0 = 0
+ ute = -1
+ paramchk = 1
+ wat = 0
+ web = 6843.8
+ wec = -25529.0
+ wlc = 0
+ wln = 1
+ wu0 = 0
+ rbdb = 50
+ xgl = -1.09e-8
+ prwb = 0
+ pub1 = 0
+ prwg = 0
+ xgw = 0
+ wub = 0
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ rbpb = 50
+ rbpd = 50
+ wtvoff = 0
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ rdsw = 100
+ tvfbsdoff = 0.022
+ tvoff = 0.00065504585
+ capmod = 2
+ ijthdfwd = 0.01
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ wku0we = 2e-11
+ mobmod = 0
+ rshg = 15.6
+ ku0we = -0.0007
+ beta0 = 13
+ leta0 = 0
+ ijthdrev = 0.01
+ nfactor = 1
+ lpdiblc2 = -1.3831831e-9
+ wvfbsdoff = 0
+ dlcig = 2.5e-9
+ lvfbsdoff = 0
+ bgidl = 2320000000.0
+ laigsd = 3.3904273e-17
+ tnom = 25
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ nigbacc = 10
+ dmcgt = 0
+ tcjsw = 0.000357
+ lkvth0we = -2e-12
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ )

.model nch_tt_6 nmos (
+ level = 54
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ vfbsdoff = 0.02
+ toxref = 3e-9
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.0069155858
+ scref = 1e-6
+ pdiblcb = -0.3
+ pigcd = 2.621
+ aigsd = 0.01077322
+ paramchk = 1
+ lvoff = -2.06441089e-9
+ ags = 2.66253
+ lvsat = 0.0015664268699999999
+ ltvoff = 1.0839662e-10
+ lvth0 = 2.2492931699999996e-9
+ bigbacc = 0.002588
+ cjd = 0.001357
+ cit = 0.00031861111
+ cjs = 0.001357
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ delta = 0.007595625
+ dlc = 3.26497e-9
+ k3b = 1.9326
+ laigc = -2.2427226e-11
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ keta = -0.52835722
+ rnoia = 0
+ rnoib = 0
+ ijthdfwd = 0.01
+ kvth0we = 0.00018
+ la0 = 3.0288889e-8
+ jsd = 6.11e-7
+ lintnoi = -1.5e-8
+ jss = 6.11e-7
+ lat = -0.00038029214
+ kt1 = -0.40872879
+ kt2 = -0.10088778
+ lk2 = -4.8654938e-10
+ lku0we = 2.5e-11
+ pketa = 0
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ ngate = 8e+20
+ bigbinv = 0.004953
+ llc = 0
+ lln = 1
+ lu0 = 1.0283078e-10
+ lcit = 1.5795656e-10
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ mjd = 0.26
+ mjs = 0.26
+ lua = 3.5218789e-17
+ lub = -1.9869262700000004e-26
+ luc = 2.2716666e-18
+ lud = 0
+ epsrox = 3.9
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ ngcon = 1
+ njd = 1.02
+ njs = 1.02
+ kt1l = 0
+ pa0 = 0
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 0
+ pbs = 0.52
+ pu0 = 0.0
+ prt = 0
+ pub = 0
+ puc = 0
+ pud = 0
+ rdsmod = 0
+ ijthdrev = 0.01
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ rsh = 17.5
+ jswgs = 1.28e-13
+ lint = 0
+ tcj = 0.00076
+ igbmod = 1
+ ua1 = 8.897383e-10
+ ub1 = -8.0235504e-19
+ uc1 = -6.3390556e-11
+ tpb = 0.0014
+ lkt1 = 9.8027184e-9
+ lkt2 = 7.8751111e-10
+ wa0 = 0
+ lpdiblc2 = 6.6256944e-15
+ lmax = 9e-8
+ ute = -1
+ wat = 0
+ web = 6843.8
+ pscbe1 = 1000000000.0
+ wec = -25529.0
+ pscbe2 = 1e-20
+ lmin = 5.4e-8
+ wlc = 0
+ wln = 1
+ wu0 = 0.0
+ xgl = -1.09e-8
+ xgw = 0
+ wub = 0
+ wuc = 0
+ wud = 0
+ lpe0 = 9.2e-8
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ pbswgd = 0.95
+ lpeb = 2.5e-7
+ pbswgs = 0.95
+ minv = -0.3
+ igcmod = 1
+ lua1 = -1.7361621e-17
+ lub1 = -8.1690078e-27
+ luc1 = 9.7666522e-18
+ ndep = 1e+18
+ lwlc = 0
+ moin = 5.1
+ nigc = 3.083
+ tvfbsdoff = 0.022
+ nfactor = 1
+ lkvth0we = -2e-12
+ tvoff = -0.00034012981
+ wtvfbsdoff = 0
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ acnqsmod = 0
+ ltvfbsdoff = 0
+ permod = 1
+ ntox = 1
+ pcit = 0.0
+ ku0we = -0.0007
+ pclm = 1.2209944
+ beta0 = 13
+ rbodymod = 0
+ leta0 = 3.0288889e-9
+ nigbacc = 10
+ letab = -2.2684433e-8
+ phin = 0.15
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ pkt1 = 0
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ voffcv = -0.16942
+ wpemod = 1
+ nigbinv = 10
+ ptvfbsdoff = 0
+ rbdb = 50
+ prwb = 0
+ pub1 = 0
+ prwg = 0
+ dmcgt = 0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ tcjsw = 0.000357
+ rdsw = 100
+ fnoimod = 1
+ eigbinv = 1.1
+ bigsd = 0.00125
+ tpbswg = 0.0009
+ wvoff = 0
+ rshg = 15.6
+ wkvth0we = 2e-12
+ wvsat = 0.0
+ wvth0 = 0.0
+ ptvoff = 0
+ trnqsmod = 0
+ cigbacc = 0.32875
+ diomod = 1
+ lketa = 2.9484719e-8
+ xpart = 1
+ pditsd = 0
+ pditsl = 0
+ tnoimod = 0
+ cjswgd = 2.82e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.82e-10
+ tnom = 25
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ egidl = 0.29734
+ a0 = -0.02222221999999996
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ rgatemod = 0
+ at = 64556.761
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = -0.035207015
+ k3 = -1.8419
+ em = 1000000.0
+ cigbinv = 0.006
+ ll = 0
+ lw = 0
+ u0 = 0.0080450556
+ tnjtsswg = 1
+ w0 = 0
+ ua = -2.404272e-9
+ ub = 1.906573466e-18
+ uc = -4.166667e-12
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 6e-9
+ mjswgd = 0.85
+ mjswgs = 0.85
+ tcjswg = 0.001
+ version = 4.5
+ wags = 0
+ tempmod = 0
+ wcit = 0.0
+ voff = -0.138884931
+ acde = 0.4
+ aigbacc = 0.02
+ vsat = 86617.64
+ wint = 0
+ vth0 = 0.326821916
+ pvoff = 0
+ wkt1 = 0
+ wmax = 0.00090001
+ aigc = 0.011713991
+ wmin = 9e-6
+ cdscb = 0
+ cdscd = 0
+ pvsat = 0.0
+ wk2we = 5e-12
+ pvth0 = 0.0
+ fprout = 300
+ drout = 0.56
+ xrcrg1 = 12
+ xrcrg2 = 1
+ aigbinv = 0.0163
+ voffl = 0
+ bigc = 0.001442
+ wwlc = 0
+ wtvoff = 0
+ weta0 = 0
+ lpclm = -1.1373478e-8
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ cgidl = 0.22
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ capmod = 2
+ wku0we = 2e-11
+ ijthsfwd = 0.01
+ poxedge = 1
+ mobmod = 0
+ pbswd = 0.8
+ pvfbsdoff = 0
+ pbsws = 0.8
+ binunit = 2
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ ijthsrev = 0.01
+ pdits = 0
+ cigsd = 0.069865
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ k2we = 5e-5
+ dsub = 0.75
+ dtox = 2.7e-10
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ eta0 = 0.26777778
+ etab = -0.0086762422
+ tnoia = 0
+ peta0 = 0
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ wketa = 0
+ tpbsw = 0.0019
+ cjswd = 8.2e-11
+ cjsws = 8.2e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ pkvth0we = -1.3e-19
+ njtsswg = 9
+ )

.model nch_tt_7 nmos (
+ level = 54
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ ltvoff = -2.4740506e-10
+ aigbacc = 0.02
+ rdsw = 100
+ ijthsfwd = 0.01
+ lku0we = 2.5e-11
+ aigbinv = 0.0163
+ epsrox = 3.9
+ rshg = 15.6
+ rdsmod = 0
+ igbmod = 1
+ ijthsrev = 0.01
+ pvoff = 0
+ cdscb = 0
+ cdscd = 0
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ pvsat = 0.0
+ wk2we = 5e-12
+ pvth0 = 0.0
+ drout = 0.56
+ pbswgd = 0.95
+ pbswgs = 0.95
+ igcmod = 1
+ poxedge = 1
+ wtvfbsdoff = 0
+ voffl = 0
+ tnom = 25
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ weta0 = 0
+ binunit = 2
+ lpclm = -7.2871722e-8
+ ltvfbsdoff = 0
+ cgidl = 0.22
+ wags = 0
+ wcit = 0.0
+ pvfbsdoff = 0
+ permod = 1
+ pbswd = 0.8
+ pbsws = 0.8
+ voff = -0.112415764
+ pkvth0we = -1.3e-19
+ acde = 0.4
+ ptvfbsdoff = 0
+ vsat = 86759.482
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ wint = 0
+ vth0 = 0.324717597
+ wkt1 = 0
+ wmax = 0.00090001
+ aigc = 0.011692671
+ pdits = 0
+ wmin = 9e-6
+ vfbsdoff = 0.02
+ cigsd = 0.069865
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ voffcv = -0.16942
+ wpemod = 1
+ wub1 = 0.0
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ bigc = 0.001442
+ paramchk = 1
+ wwlc = 0
+ tnoia = 0
+ cdsc = 0
+ cgbo = 0
+ njtsswg = 9
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ peta0 = 0
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ tpbsw = 0.0019
+ ijthdfwd = 0.01
+ tpbswg = 0.0009
+ ckappad = 0.6
+ cjswd = 8.2e-11
+ ckappas = 0.6
+ cjsws = 8.2e-11
+ mjswd = 0.11
+ pdiblc1 = 0
+ pdiblc2 = 0.0069157
+ mjsws = 0.11
+ agidl = 9.41e-8
+ pdiblcb = -0.3
+ ptvoff = 0
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ ijthdrev = 0.01
+ bigbacc = 0.002588
+ diomod = 1
+ k2we = 5e-5
+ dsub = 0.75
+ scref = 1e-6
+ dtox = 2.7e-10
+ pditsd = 0
+ pditsl = 0
+ kvth0we = 0.00018
+ cjswgd = 2.82e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.82e-10
+ ags = 2.66253
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ pigcd = 2.621
+ aigsd = 0.01077322
+ cjd = 0.001357
+ cit = -0.0027423847
+ cjs = 0.001357
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ lintnoi = -1.5e-8
+ dlc = 3.26497e-9
+ bigbinv = 0.004953
+ k3b = 1.9326
+ lvoff = -3.599622200000001e-9
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ eta0 = 0.35179556
+ etab = -1.0973583
+ lvsat = 0.0015582000999999996
+ mjswgd = 0.85
+ mjswgs = 0.85
+ lvth0 = 2.3713433000000004e-9
+ la0 = -3.1577778e-7
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = 0.0075786667
+ lkvth0we = -2e-12
+ kt1 = 0.010917511
+ kt2 = -0.10990444
+ lk2 = -1.5787889e-9
+ delta = 0.007595625
+ tcjswg = 0.001
+ llc = 0
+ laigc = -2.1190647e-11
+ lln = 1
+ lu0 = 5.4692711e-10
+ mjd = 0.26
+ mjs = 0.26
+ lua = 7.8730998e-17
+ lub = -4.3148946000000005e-26
+ luc = 1.578889e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 0
+ rnoia = 0
+ rnoib = 0
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 0.0
+ pbs = 0.52
+ pu0 = 0.0
+ prt = 0
+ pub = 0
+ puc = 0
+ pud = 0
+ acnqsmod = 0
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 3.744227e-10
+ ngate = 8e+20
+ ub1 = -1.4506222e-18
+ uc1 = -1.6722222e-10
+ tpb = 0.0014
+ ngcon = 1
+ wa0 = 0
+ ute = -1
+ wat = 0.0
+ web = 6843.8
+ wec = -25529.0
+ wlc = 0
+ wln = 1
+ wu0 = 0.0
+ xgl = -1.09e-8
+ xgw = 0
+ wub = 0
+ wuc = 0
+ wud = 0
+ rbodymod = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ a0 = 5.9444444
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = -72666.667
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = -0.016375299
+ k3 = -1.8419
+ em = 1000000.0
+ fprout = 300
+ ll = 0
+ lw = 0
+ u0 = 0.00038822222
+ nfactor = 1
+ w0 = 0
+ ua = -3.1544825e-9
+ ub = 2.30794738e-18
+ uc = 7.77778e-12
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 6e-9
+ xrcrg1 = 12
+ xrcrg2 = 1
+ wtvoff = 0
+ tvfbsdoff = 0.022
+ nigbacc = 10
+ capmod = 2
+ tvoff = 0.0057943818
+ wku0we = 2e-11
+ keta = 0.088888889
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ mobmod = 0
+ nigbinv = 10
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 3.3549431e-10
+ kt1l = 0
+ ku0we = -0.0007
+ wkvth0we = 2e-12
+ beta0 = 13
+ leta0 = -1.8441422e-9
+ letab = 4.0459126e-8
+ lint = 0
+ trnqsmod = 0
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ lkt1 = -1.4536767e-8
+ lkt2 = 1.3104778e-9
+ lmax = 5.4e-8
+ lmin = 4.5e-8
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ lpe0 = 9.2e-8
+ fnoimod = 1
+ lpeb = 2.5e-7
+ eigbinv = 1.1
+ minv = -0.3
+ lua1 = 1.2526683e-17
+ lub1 = 2.9430489e-26
+ luc1 = 1.5788889e-17
+ ndep = 1e+18
+ dmcgt = 0
+ rgatemod = 0
+ lwlc = 0
+ tcjsw = 0.000357
+ moin = 5.1
+ tnjtsswg = 1
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ nigc = 3.083
+ bigsd = 0.00125
+ noff = 2.7195
+ cigbacc = 0.32875
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ wvoff = 0
+ tnoimod = 0
+ ntox = 1
+ pcit = 0.0
+ pclm = 2.281309
+ wvsat = 0.0
+ wvth0 = 0.0
+ cigbinv = 0.006
+ phin = 0.15
+ toxref = 3e-9
+ pkt1 = 0
+ lketa = -6.3155556e-9
+ version = 4.5
+ xpart = 1
+ tempmod = 0
+ egidl = 0.29734
+ rbdb = 50
+ prwb = 0
+ pub1 = 0.0
+ prwg = 0
+ )

.model nch_tt_8 nmos (
+ level = 54
+ ngate = 8e+20
+ ngcon = 1
+ wpclm = 0
+ rdsmod = 0
+ wkvth0we = 2e-12
+ wtvfbsdoff = 0
+ igbmod = 1
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ trnqsmod = 0
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ nigbacc = 10
+ ltvfbsdoff = 0
+ pbswgd = 0.95
+ pbswgs = 0.95
+ k2we = 5e-5
+ igcmod = 1
+ dsub = 0.75
+ dtox = 2.7e-10
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ nigbinv = 10
+ rgatemod = 0
+ eta0 = -0.001232
+ etab = -0.88502038
+ tnjtsswg = 1
+ tvfbsdoff = 0.022
+ ptvfbsdoff = 0
+ tvoff = 0.0030235155
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ fnoimod = 1
+ permod = 1
+ eigbinv = 1.1
+ ku0we = -0.0007
+ beta0 = 13
+ leta0 = 1.5454208e-8
+ letab = 3.0054568e-8
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ ppclm = 0
+ voffcv = -0.16942
+ wpemod = 1
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ cigbacc = 0.32875
+ dmcgt = 0
+ tnoimod = 0
+ tcjsw = 0.000357
+ cigbinv = 0.006
+ tpbswg = 0.0009
+ keta = 0.44888889
+ ijthsfwd = 0.01
+ bigsd = 0.00125
+ version = 4.5
+ wvoff = 0
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 3.0392239e-10
+ tempmod = 0
+ kt1l = 0
+ ptvoff = 0
+ wvsat = 0.0
+ wvth0 = 0.0
+ ijthsrev = 0.01
+ lint = 0
+ aigbacc = 0.02
+ lkt1 = -3.9088498e-9
+ lkt2 = 1.6072e-9
+ diomod = 1
+ lmax = 4.5e-8
+ lmin = 3.6e-8
+ lpe0 = 9.2e-8
+ pditsd = 0
+ pditsl = 0
+ lketa = -2.3955556e-8
+ lpeb = 2.5e-7
+ cjswgd = 2.82e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.82e-10
+ xpart = 1
+ minv = -0.3
+ aigbinv = 0.0163
+ lua1 = 7.1708778e-18
+ lub1 = -2.3942999e-26
+ luc1 = -1.63268e-17
+ egidl = 0.29734
+ ndep = 1e+18
+ lwlc = 0
+ mjswgd = 0.85
+ mjswgs = 0.85
+ moin = 5.1
+ nigc = 3.083
+ tcjswg = 0.001
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ poxedge = 1
+ pkvth0we = -1.3e-19
+ ntox = 1
+ pcit = 0.0
+ pclm = 2.10165423
+ binunit = 2
+ pvoff = 0
+ fprout = 300
+ phin = 0.15
+ cdscb = 0
+ cdscd = 0
+ vfbsdoff = 0.02
+ pvsat = 0.0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ wk2we = 5e-12
+ pvth0 = 0.0
+ drout = 0.56
+ pkt1 = 0
+ voffl = 0
+ wtvoff = 0
+ paramchk = 1
+ weta0 = 0
+ rbdb = 50
+ prwb = 0
+ pub1 = 0.0
+ prwg = 0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ lpclm = -6.406864000000001e-8
+ rdsw = 100
+ capmod = 2
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ cgidl = 0.22
+ wku0we = 2e-11
+ mobmod = 0
+ ijthdfwd = 0.01
+ a0 = 3.6555556
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 123237.73
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.024156861
+ k3 = -1.8419
+ em = 1000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.0044833333
+ pvfbsdoff = 0
+ w0 = 0
+ ua = -2.2580401200000003e-9
+ ub = 1.5627388499999998e-18
+ uc = 2.4e-10
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 6e-9
+ pbswd = 0.8
+ pbsws = 0.8
+ rshg = 15.6
+ ijthdrev = 0.01
+ pdits = 0
+ njtsswg = 9
+ cigsd = 0.069865
+ laigsd = -2.1777778e-17
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ ckappad = 0.6
+ ckappas = 0.6
+ pk2we = -1e-19
+ tnom = 25
+ pdiblc1 = 0
+ pdiblc2 = 0.0069157
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ pdiblcb = -0.3
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ tnoia = 0
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ peta0 = 0
+ lkvth0we = -2e-12
+ bigbacc = 0.002588
+ tpbsw = 0.0019
+ wags = 0
+ cjswd = 8.2e-11
+ cjsws = 8.2e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ wcit = 0.0
+ kvth0we = 0.00018
+ acnqsmod = 0
+ voff = -0.039834349000000005
+ acde = 0.4
+ lintnoi = -1.5e-8
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ vsat = 85481.92200000002
+ rbodymod = 0
+ vtsswgs = 4.2
+ wint = 0
+ vth0 = 0.35076130299999997
+ toxref = 3e-9
+ wkt1 = 0
+ ags = 2.66253
+ wmax = 0.00090001
+ aigc = 0.011387162
+ wmin = 9e-6
+ cjd = 0.001357
+ cit = -0.0020980598
+ cjs = 0.001357
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 3.26497e-9
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ scref = 1e-6
+ wub1 = 0.0
+ pigcd = 2.621
+ aigsd = 0.010773221
+ la0 = -2.0362223e-7
+ bigc = 0.001442
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.0020206488
+ kt1 = -0.20597876
+ kt2 = -0.11596
+ lk2 = -3.5648647e-9
+ wwlc = 0
+ llc = 0
+ lvoff = -7.156111900000001e-9
+ lln = 1
+ lu0 = 3.4626667e-10
+ mjd = 0.26
+ mjs = 0.26
+ lua = 3.4805321000000004e-17
+ lub = -6.633731000000002e-27
+ luc = -9.7999999e-18
+ lud = 0
+ ltvoff = -1.1163261e-10
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 0
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 0.0
+ pbs = 0.52
+ pk2 = 0
+ lvsat = 0.0016208003899999999
+ cdsc = 0
+ pu0 = 0.0
+ lvth0 = 1.0952018800000002e-9
+ prt = 0
+ cgbo = 0
+ pua = 0
+ pub = 0
+ puc = 0
+ pud = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ delta = 0.007595625
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 4.8372486e-10
+ ub1 = -3.6136738e-19
+ cigc = 0.000625
+ laigc = -6.2207351e-12
+ uc1 = 4.882e-10
+ tpb = 0.0014
+ wa0 = 0
+ rnoia = 0
+ rnoib = 0
+ nfactor = 1
+ ute = -1
+ wat = 0.0
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 0
+ wlc = 0
+ lku0we = 2.5e-11
+ wln = 1
+ wu0 = 0.0
+ xgl = -1.09e-8
+ xgw = 0
+ wua = 0
+ wub = 0
+ wuc = 0
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ epsrox = 3.9
+ )

.model nch_tt_9 nmos (
+ level = 54
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ ptvfbsdoff = 0
+ voffl = 0
+ minv = -0.3
+ lub1 = 0
+ weta0 = 0
+ ndep = 1e+18
+ wetab = -1.0073378e-8
+ lwlc = 0
+ moin = 5.1
+ nigc = 3.083
+ cgidl = 0.22
+ lkvth0we = -2e-12
+ njtsswg = 9
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ pvfbsdoff = 0
+ noic = 45200000.0
+ permod = 1
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ acnqsmod = 0
+ pbswd = 0.8
+ pbsws = 0.8
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.018557155
+ pdiblcb = -0.3
+ ntox = 1
+ pcit = 0
+ pclm = 1.4152454
+ rbodymod = 0
+ phin = 0.15
+ voffcv = -0.16942
+ wpemod = 1
+ pdits = 0
+ cigsd = 0.069865
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ pkt1 = 0
+ bigbacc = 0.002588
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ kvth0we = 0.00018
+ rbdb = 50
+ prwb = 0
+ pub1 = 0
+ prwg = 0
+ wpdiblc2 = -1.7177628e-11
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ lintnoi = -1.5e-8
+ tnoia = 0
+ bigbinv = 0.004953
+ rdsw = 100
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ peta0 = 0
+ tpbswg = 0.0009
+ wketa = 3.3422159e-8
+ tpbsw = 0.0019
+ cjswd = 8.2e-11
+ cjsws = 8.2e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ ags = 0.87683314
+ ptvoff = 0
+ cjd = 0.001357
+ cit = 4.8708935e-5
+ cjs = 0.001357
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ wkvth0we = 2e-12
+ bvs = 8.7
+ rshg = 15.6
+ waigsd = 3.0716751e-12
+ dlc = 9.8024918e-9
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ trnqsmod = 0
+ diomod = 1
+ la0 = 0
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = 0
+ kt1 = -0.19515831
+ kt2 = -0.052853133
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 2.82e-10
+ llc = 0
+ pku0we = -1.5e-18
+ lln = 1
+ cjswgs = 2.82e-10
+ lu0 = 0
+ mjd = 0.26
+ mjs = 0.26
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ scref = 1e-6
+ njd = 1.02
+ njs = 1.02
+ pa0 = 0
+ nfactor = 1
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 0
+ pbs = 0.52
+ pigcd = 2.621
+ aigsd = 0.010772879
+ pu0 = 0
+ prt = 0
+ pud = 0
+ tnom = 25
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 1.311952e-9
+ toxe = 2.43e-9
+ ub1 = -8.0649865e-19
+ toxm = 2.43e-9
+ lvoff = 0
+ uc1 = 3.0375074e-11
+ mjswgd = 0.85
+ mjswgs = 0.85
+ tpb = 0.0014
+ rgatemod = 0
+ wa0 = -2.5183444e-7
+ ute = -0.96248296
+ wat = 0
+ tnjtsswg = 1
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -3.7920026e-9
+ lvsat = 0
+ wlc = 0
+ tcjswg = 0.001
+ wln = 1
+ wu0 = -2.6190782e-10
+ xgl = -1.09e-8
+ xgw = 0
+ lvth0 = 0
+ wua = -4.0765791e-17
+ wub = 4.0599742e-26
+ wuc = -7.8572347e-18
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ delta = 0.007595625
+ nigbacc = 10
+ rnoia = 0
+ rnoib = 0
+ wags = -8.4054279e-8
+ wcit = 4.6192733e-10
+ ngate = 8e+20
+ voff = -0.11308442
+ ngcon = 1
+ wpclm = -1.3730014e-7
+ acde = 0.4
+ nigbinv = 10
+ vsat = 103058.98
+ wint = 0
+ gbmin = 1e-12
+ vth0 = 0.35034845
+ fprout = 300
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ wkt1 = -4.5639654e-8
+ wkt2 = -3.5741805e-9
+ wmax = 9e-6
+ xrcrg1 = 12
+ xrcrg2 = 1
+ aigc = 0.011766468
+ wmin = 9e-7
+ wtvoff = -8.3463378e-10
+ wua1 = -7.3834184e-16
+ wub1 = 7.3798399e-25
+ wuc1 = -8.5623711e-19
+ fnoimod = 1
+ bigc = 0.001442
+ wute = -4.0092044e-7
+ eigbinv = 1.1
+ wwlc = 0
+ tvfbsdoff = 0.022
+ capmod = 2
+ cdsc = 0
+ cgbo = 0
+ wku0we = 2e-11
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ tvoff = 0.0020036382
+ cigc = 0.000625
+ mobmod = 0
+ xjbvd = 1
+ ijthsfwd = 0.01
+ xjbvs = 1
+ lk2we = -1.5e-12
+ cigbacc = 0.32875
+ ku0we = -0.0007
+ beta0 = 13
+ leta0 = 0
+ tnoimod = 0
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ ijthsrev = 0.01
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ cigbinv = 0.006
+ dlcig = 2.5e-9
+ k2we = 5e-5
+ bgidl = 2320000000.0
+ dsub = 0.75
+ dtox = 2.7e-10
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ a0 = 3.277963
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ version = 4.5
+ at = 72000
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.025022307
+ k3 = -1.8419
+ em = 1000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.015699082
+ dmcgt = 0
+ w0 = 0
+ tempmod = 0
+ ua = -1.8192461e-9
+ ub = 2.0991879e-18
+ uc = 7.4172444e-11
+ ud = 0
+ eta0 = 0.3
+ tcjsw = 0.000357
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ alpha0 = 2e-10
+ ww = 0
+ alpha1 = 3.6
+ xw = 6e-9
+ etab = -0.24888148
+ aigbacc = 0.02
+ bigsd = 0.00125
+ wvoff = 2.3777201e-9
+ pkvth0we = -1.3e-19
+ aigbinv = 0.0163
+ wvsat = -0.0017920539
+ wvth0 = -1.1145485e-8
+ toxref = 3e-9
+ waigc = 2.6350949e-11
+ vfbsdoff = 0.02
+ xpart = 1
+ paramchk = 1
+ ltvoff = 0
+ egidl = 0.29734
+ poxedge = 1
+ binunit = 2
+ wtvfbsdoff = 0
+ keta = -0.063711099
+ lku0we = 2.5e-11
+ ijthdfwd = 0.01
+ epsrox = 3.9
+ ltvfbsdoff = 0
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 0
+ rdsmod = 0
+ kt1l = 0
+ igbmod = 1
+ ijthdrev = 0.01
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ pvoff = 0
+ lint = 6.5375218e-9
+ pbswgd = 0.95
+ cdscb = 0
+ cdscd = 0
+ pbswgs = 0.95
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ lkt1 = 0
+ pvsat = 0
+ lmax = 2.001e-5
+ wk2we = 5e-12
+ pvth0 = 0
+ lmin = 8.9991e-6
+ drout = 0.56
+ igcmod = 1
+ )

.model nch_tt_10 nmos (
+ level = 54
+ xrcrg1 = 12
+ xrcrg2 = 1
+ cgidl = 0.22
+ vfbsdoff = 0.02
+ wtvoff = -8.9580408e-10
+ nfactor = 1
+ pbswd = 0.8
+ pbsws = 0.8
+ paramchk = 1
+ capmod = 2
+ wku0we = 2e-11
+ mobmod = 0
+ pdits = 0
+ cigsd = 0.069865
+ nigbacc = 10
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ ijthdfwd = 0.01
+ keta = -0.064075044
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ nigbinv = 10
+ lags = -6.3328546e-8
+ wtvfbsdoff = 0
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 1.1337416e-9
+ tnoia = 0
+ laigsd = 1.1048614e-17
+ ijthdrev = 0.01
+ kt1l = 0
+ peta0 = 0
+ ltvfbsdoff = 0
+ lpdiblc2 = -6.1589259e-10
+ wketa = 3.7630763e-8
+ lint = 6.5375218e-9
+ tpbsw = 0.0019
+ lkt1 = -4.5537316e-8
+ lkt2 = -1.2972142e-8
+ cjswd = 8.2e-11
+ lmax = 8.9991e-6
+ cjsws = 8.2e-11
+ lmin = 8.9908e-7
+ fnoimod = 1
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ lpe0 = 9.2e-8
+ eigbinv = 1.1
+ lpeb = 2.5e-7
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ minv = -0.3
+ lua1 = -4.3996966e-16
+ lub1 = 2.6060002e-25
+ luc1 = 3.9191378e-17
+ ndep = 1e+18
+ lute = -3.7058959e-8
+ lwlc = 0
+ ptvfbsdoff = 0
+ moin = 5.1
+ lkvth0we = -2e-12
+ nigc = 3.083
+ scref = 1e-6
+ pigcd = 2.621
+ aigsd = 0.010772879
+ cigbacc = 0.32875
+ acnqsmod = 0
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ lvoff = -1.4242682e-8
+ toxref = 3e-9
+ tnoimod = 0
+ pags = 2.8299487e-13
+ rbodymod = 0
+ lvsat = 0
+ lvth0 = 5.1255324e-8
+ ntox = 1
+ pcit = -1.846418e-16
+ pclm = 1.4152454
+ cigbinv = 0.006
+ delta = 0.007595625
+ laigc = -1.4938914e-10
+ tvfbsdoff = 0.022
+ rnoia = 0
+ rnoib = 0
+ phin = 0.15
+ pkt1 = 4.9872912e-14
+ pkt2 = 1.3351872e-15
+ pketa = -3.7835355e-14
+ version = 4.5
+ ngate = 8e+20
+ ltvoff = -2.0733557e-10
+ ngcon = 1
+ tempmod = 0
+ wpclm = -1.3730014e-7
+ wpdiblc2 = -4.8108443e-11
+ gbmin = 1e-12
+ rbdb = 50
+ pua1 = 6.0905252e-22
+ prwb = 0
+ prwg = 0
+ pub1 = -5.9738158e-31
+ jswgd = 1.28e-13
+ puc1 = 1.7562426e-23
+ jswgs = 1.28e-13
+ rbpb = 50
+ rbpd = 50
+ aigbacc = 0.02
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ pute = 3.9602525e-13
+ lku0we = 2.5e-11
+ rdsw = 100
+ wvfbsdoff = 0
+ epsrox = 3.9
+ lvfbsdoff = 0
+ rdsmod = 0
+ aigbinv = 0.0163
+ igbmod = 1
+ wkvth0we = 2e-12
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ pbswgd = 0.95
+ pbswgs = 0.95
+ rshg = 15.6
+ trnqsmod = 0
+ tvoff = 0.0020267011
+ igcmod = 1
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ poxedge = 1
+ ku0we = -0.0007
+ beta0 = 13
+ tnom = 25
+ rgatemod = 0
+ leta0 = 0
+ binunit = 2
+ tnjtsswg = 1
+ toxe = 2.43e-9
+ paigsd = -9.9503825e-23
+ toxm = 2.43e-9
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ permod = 1
+ wags = -1.1553313e-7
+ wcit = 4.8246591e-10
+ dmcgt = 0
+ tcjsw = 0.000357
+ voff = -0.11150014
+ acde = 0.4
+ voffcv = -0.16942
+ wpemod = 1
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ vsat = 103058.98
+ wint = 0
+ vth0 = 0.34464708
+ wkt1 = -5.1187253e-8
+ wkt2 = -3.7226997e-9
+ wmax = 9e-6
+ aigc = 0.011783086
+ bigsd = 0.00125
+ wmin = 9e-7
+ wvoff = 2.6904676e-9
+ wua1 = -8.0608962e-16
+ wub1 = 8.0443355e-25
+ wuc1 = -2.8097884e-18
+ wvsat = -0.0017920539
+ wvth0 = -1.1528173e-8
+ bigc = 0.001442
+ wute = -4.4497219e-7
+ wwlc = 0
+ waigc = 2.7413515e-11
+ tpbswg = 0.0009
+ njtsswg = 9
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ lketa = 3.2718606e-9
+ xtsswgd = 0.18
+ cgsl = 3.31989e-12
+ ijthsfwd = 0.01
+ cgso = 4.90562e-11
+ xtsswgs = 0.18
+ cigc = 0.000625
+ xpart = 1
+ ckappad = 0.6
+ ckappas = 0.6
+ ptvoff = 5.4992103e-16
+ pdiblc1 = 0
+ pdiblc2 = 0.018625664
+ pdiblcb = -0.3
+ waigsd = 3.0716862e-12
+ egidl = 0.29734
+ diomod = 1
+ ijthsrev = 0.01
+ pditsd = 0
+ pditsl = 0
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ cjswgd = 2.82e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.82e-10
+ ags = 0.88387747
+ bigbacc = 0.002588
+ cjd = 0.001357
+ cit = -7.7402473e-5
+ cjs = 0.001357
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 9.8024918e-9
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ k2we = 5e-5
+ kvth0we = 0.00018
+ dsub = 0.75
+ dtox = 2.7e-10
+ mjswgd = 0.85
+ mjswgs = 0.85
+ pvfbsdoff = 0
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ la0 = -2.0592205e-6
+ lintnoi = -1.5e-8
+ ppdiblc2 = 2.7806803e-16
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = 0.094482725
+ tcjswg = 0.001
+ kt1 = -0.19009298
+ lk2 = -1.3154073e-8
+ kt2 = -0.051410181
+ bigbinv = 0.004953
+ llc = 0
+ vtsswgd = 4.2
+ lln = 1
+ vtsswgs = 4.2
+ lu0 = -1.9964409e-9
+ mjd = 0.26
+ lua = -2.2049077e-16
+ mjs = 0.26
+ lub = -1.5408759e-27
+ luc = 1.1211784e-18
+ lud = 0
+ pvoff = -2.8116001e-15
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 3.0846188e-13
+ eta0 = 0.3
+ nsd = 1e+20
+ pbd = 0.52
+ pat = -8.2787187e-9
+ pbs = 0.52
+ pk2 = -1.9754424e-15
+ cdscb = 0
+ cdscd = 0
+ etab = -0.24888148
+ pu0 = 9.9503831e-18
+ pvsat = 0
+ prt = 0
+ pua = 2.7693259e-23
+ pub = -6.3482817e-32
+ puc = -1.7214163e-23
+ pud = 0
+ wk2we = 5e-12
+ pvth0 = 3.4403639e-15
+ drout = 0.56
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 1.3608919e-9
+ ub1 = -8.3548641e-19
+ uc1 = 2.6015633e-11
+ paigc = -9.5524673e-18
+ tpb = 0.0014
+ wa0 = -2.8614611e-7
+ ute = -0.95836072
+ wat = 0.00092088084
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -3.5722648e-9
+ voffl = 0
+ wlc = 0
+ wln = 1
+ wu0 = -2.6301465e-10
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -4.3846243e-17
+ wub = 4.7661234e-26
+ wuc = -5.9424224e-18
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ a0 = 3.5070197
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ weta0 = 0
+ pkvth0we = -1.3e-19
+ at = 61490.242
+ cf = 8.15e-11
+ wetab = -1.0073378e-8
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.026485497
+ k3 = -1.8419
+ em = 1000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.015921155
+ fprout = 300
+ w0 = 0
+ ua = -1.7947198e-9
+ ub = 2.0993593e-18
+ uc = 7.4047731e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 6e-9
+ )

.model nch_tt_11 nmos (
+ level = 54
+ ku0we = -0.0007
+ beta0 = 13
+ wku0we = 2e-11
+ leta0 = 0
+ rbdb = 50
+ mobmod = 0
+ pua1 = 9.7840116e-23
+ prwb = 0
+ prwg = 0
+ pub1 = -1.2240721e-31
+ puc1 = -3.5940917e-24
+ a0 = 1.2386098
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ wtvfbsdoff = 0
+ at = 220073.87
+ cf = 8.15e-11
+ rbpb = 50
+ rbpd = 50
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.025732723
+ k3 = -1.8419
+ rbps = 50
+ em = 1000000.0
+ rbsb = 50
+ pvag = 1.2
+ ll = 0
+ lw = 0
+ u0 = 0.015421688
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ w0 = 0
+ ua = -1.9419497e-9
+ ub = 2.1613601e-18
+ uc = 9.7509556e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 6e-9
+ rdsw = 100
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ ijthsfwd = 0.01
+ ltvfbsdoff = 0
+ dmcgt = 0
+ tcjsw = 0.000357
+ laigsd = -9.7335958e-18
+ ijthsrev = 0.01
+ rshg = 15.6
+ njtsswg = 9
+ bigsd = 0.00125
+ ptvfbsdoff = 0
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ wvoff = -7.7864574e-9
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.014827337
+ pdiblcb = -0.3
+ wvsat = -0.0017920539
+ ppdiblc2 = 2.4623293e-15
+ tnom = 25
+ wvth0 = -1.2261894e-9
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ waigc = -9.5733062e-12
+ lketa = -3.0044615e-8
+ bigbacc = 0.002588
+ xpart = 1
+ wags = 1.2460313e-6
+ kvth0we = 0.00018
+ toxref = 3e-9
+ egidl = 0.29734
+ pkvth0we = -1.3e-19
+ wcit = 1.5976377e-10
+ ags = 0.23741392
+ cjd = 0.001357
+ cit = 0.0013334381
+ voff = -0.11121991
+ lintnoi = -1.5e-8
+ cjs = 0.001357
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ acde = 0.4
+ dlc = 9.8024918e-9
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ k3b = 1.9326
+ vtsswgs = 4.2
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ vsat = 103058.98
+ wint = 0
+ vfbsdoff = 0.02
+ vth0 = 0.39319507
+ wkt1 = 1.7828643e-8
+ wkt2 = -3.7425887e-9
+ wmax = 9e-6
+ la0 = -4.0335612e-8
+ aigc = 0.011680759
+ wmin = 9e-7
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.0466567
+ kt1 = -0.22273968
+ lk2 = -1.2484105e-8
+ kt2 = -0.052902736
+ llc = 0
+ lln = 1
+ lu0 = -1.5519156e-9
+ mjd = 0.26
+ ltvoff = -6.7137092e-10
+ lua = -8.9456155e-17
+ mjs = 0.26
+ lub = -5.6721601e-26
+ luc = -1.9759846e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = -3.420874e-13
+ nsd = 1e+20
+ pbd = 0.52
+ pat = -3.6466881e-9
+ pbs = 0.52
+ pk2 = 6.3553328e-16
+ pvfbsdoff = 0
+ paramchk = 1
+ pu0 = 2.6298232e-17
+ wua1 = -2.3169366e-16
+ wub1 = 2.7075449e-25
+ prt = 0
+ wuc1 = 2.096158e-17
+ pua = -3.3732216e-24
+ pub = 1.7089792e-32
+ puc = 7.8894695e-24
+ pud = 0
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 9.9427719e-10
+ bigc = 0.001442
+ ub1 = -5.7879508e-19
+ uc1 = 6.536871e-11
+ pvoff = 6.5128631e-15
+ tpb = 0.0014
+ wwlc = 0
+ wa0 = 4.4480813e-7
+ ute = -1
+ wat = -0.0042836479
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -6.5059453e-9
+ cdscb = 0
+ cdscd = 0
+ lku0we = 2.5e-11
+ wlc = 0
+ wln = 1
+ wu0 = -2.8138302e-10
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -8.9400845e-18
+ wub = -4.2869787e-26
+ pvsat = 0
+ wuc = -3.4148751e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ epsrox = 3.9
+ cdsc = 0
+ wk2we = 5e-12
+ pvth0 = -5.7284018e-15
+ drout = 0.56
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ ijthdfwd = 0.01
+ cgsl = 3.31989e-12
+ paigc = 2.3365803e-17
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ rdsmod = 0
+ nfactor = 1
+ voffl = 0
+ igbmod = 1
+ weta0 = 0
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ wetab = -1.0073378e-8
+ pbswgd = 0.95
+ pbswgs = 0.95
+ ijthdrev = 0.01
+ igcmod = 1
+ cgidl = 0.22
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ lpdiblc2 = 2.7646188e-9
+ nigbacc = 10
+ k2we = 5e-5
+ pbswd = 0.8
+ pbsws = 0.8
+ dsub = 0.75
+ dtox = 2.7e-10
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ nigbinv = 10
+ paigsd = 8.7660773e-23
+ eta0 = 0.3
+ pdits = 0
+ etab = -0.24888148
+ cigsd = 0.069865
+ lkvth0we = -2e-12
+ permod = 1
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ pk2we = -1e-19
+ fnoimod = 1
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ acnqsmod = 0
+ eigbinv = 1.1
+ voffcv = -0.16942
+ wpemod = 1
+ tnoia = 0
+ rbodymod = 0
+ peta0 = 0
+ wketa = -4.0591301e-8
+ tpbsw = 0.0019
+ cjswd = 8.2e-11
+ cjsws = 8.2e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ cigbacc = 0.32875
+ wpdiblc2 = -2.5023346e-9
+ tnoimod = 0
+ tpbswg = 0.0009
+ cigbinv = 0.006
+ scref = 1e-6
+ ptvoff = 2.4706364e-16
+ pigcd = 2.621
+ keta = -0.026640801
+ aigsd = 0.010772879
+ waigsd = 3.0714759e-12
+ version = 4.5
+ lvoff = -1.4492081e-8
+ lags = 5.1202402e-7
+ wkvth0we = 2e-12
+ tempmod = 0
+ jswd = 1.28e-13
+ diomod = 1
+ jsws = 1.28e-13
+ lcit = -1.2190653e-10
+ lvsat = 0
+ kt1l = 0
+ lvth0 = 8.0476154e-9
+ pditsd = 0
+ pditsl = 0
+ trnqsmod = 0
+ cjswgd = 2.82e-10
+ tvfbsdoff = 0.022
+ pku0we = -1.5e-18
+ cjswgs = 2.82e-10
+ delta = 0.007595625
+ laigc = -5.8318716e-11
+ aigbacc = 0.02
+ lint = 6.5375218e-9
+ rnoia = 0
+ rnoib = 0
+ lkt1 = -1.6481753e-8
+ lkt2 = -1.1643768e-8
+ lmax = 8.9908e-7
+ lmin = 4.4908e-7
+ pketa = 3.1782283e-14
+ mjswgd = 0.85
+ lpe0 = 9.2e-8
+ ngate = 8e+20
+ mjswgs = 0.85
+ lpeb = 2.5e-7
+ ngcon = 1
+ wpclm = -1.3730014e-7
+ aigbinv = 0.0163
+ tcjswg = 0.001
+ minv = -0.3
+ rgatemod = 0
+ lua1 = -1.1368255e-16
+ lub1 = 3.2144732e-26
+ luc1 = 4.1671397e-18
+ gbmin = 1e-12
+ tnjtsswg = 1
+ ndep = 1e+18
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ lwlc = 0
+ moin = 5.1
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ nigc = 3.083
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ poxedge = 1
+ fprout = 300
+ xrcrg1 = 12
+ xrcrg2 = 1
+ pags = -9.2879744e-13
+ ntox = 1
+ pcit = 1.025631e-16
+ binunit = 2
+ pclm = 1.4152454
+ tvoff = 0.0025480892
+ wtvoff = -5.5551488e-10
+ xjbvd = 1
+ phin = 0.15
+ xjbvs = 1
+ lk2we = -1.5e-12
+ pkt1 = -1.1551235e-14
+ pkt2 = 1.3528884e-15
+ capmod = 2
+ )

.model nch_tt_12 nmos (
+ level = 54
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ ptvfbsdoff = 0
+ cigbacc = 0.32875
+ laigsd = -9.015225e-17
+ wkvth0we = 2e-12
+ tnoia = 0
+ tnoimod = 0
+ trnqsmod = 0
+ peta0 = 0
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ wketa = 1.7936379e-8
+ tpbsw = 0.0019
+ a0 = 1.7327189
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ cigbinv = 0.006
+ at = 153009.14
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.019241707
+ k3 = -1.8419
+ em = 1000000.0
+ cjswd = 8.2e-11
+ ll = -1.18e-13
+ cjsws = 8.2e-11
+ lw = 0
+ u0 = 0.013315621
+ w0 = 0
+ mjswd = 0.11
+ ua = -2.1226101e-9
+ ub = 2.1428106e-18
+ uc = 6.8443458e-11
+ ud = 0
+ mjsws = 0.11
+ agidl = 9.41e-8
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 6e-9
+ k2we = 5e-5
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ dsub = 0.75
+ dtox = 2.7e-10
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ version = 4.5
+ rgatemod = 0
+ tnjtsswg = 1
+ tempmod = 0
+ eta0 = 0.3
+ etab = -0.24888148
+ aigbacc = 0.02
+ scref = 1e-6
+ pigcd = 2.621
+ aigsd = 0.010772879
+ toxref = 3e-9
+ lvoff = -6.0911145e-9
+ aigbinv = 0.0163
+ lvsat = 0
+ lvth0 = -4.941492e-9
+ tvfbsdoff = 0.022
+ delta = 0.007595625
+ laigc = -1.9233809e-11
+ rnoia = 0
+ rnoib = 0
+ ltvoff = -1.0250882e-10
+ pketa = 6.0301037e-15
+ ngate = 8e+20
+ ngcon = 1
+ wpclm = -2.8227848e-7
+ poxedge = 1
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ lku0we = 2.5e-11
+ wvfbsdoff = 0
+ epsrox = 3.9
+ lvfbsdoff = 0
+ binunit = 2
+ rdsmod = 0
+ ijthsfwd = 0.01
+ igbmod = 1
+ keta = -0.041938217
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ lags = 4.5664516e-7
+ pbswgd = 0.95
+ pbswgs = 0.95
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 1.6914929e-10
+ ijthsrev = 0.01
+ igcmod = 1
+ kt1l = 0
+ tvoff = 0.0012552207
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ lint = 9.7879675e-9
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ lkt1 = -9.5958544e-9
+ lkt2 = -3.7159363e-9
+ lmax = 4.4908e-7
+ lmin = 2.1577e-7
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ ku0we = -0.0007
+ paigsd = 8.167794e-23
+ ppdiblc2 = -2.773275e-15
+ beta0 = 13
+ minv = -0.3
+ lua1 = -3.2594611e-17
+ lub1 = -2.740043e-26
+ leta0 = 0
+ luc1 = -3.5163101e-18
+ ndep = 1e+18
+ ppclm = 6.379047e-14
+ lwlc = 0
+ permod = 1
+ moin = 5.1
+ dlcig = 2.5e-9
+ nigc = 3.083
+ bgidl = 2320000000.0
+ njtsswg = 9
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ pkvth0we = -1.3e-19
+ dmcgt = 0
+ voffcv = -0.16942
+ ckappad = 0.6
+ wpemod = 1
+ ckappas = 0.6
+ tcjsw = 0.000357
+ pdiblc1 = 0
+ pdiblc2 = 0.026288388
+ pags = 8.4375107e-13
+ pdiblcb = -0.3
+ ntox = 1
+ pcit = -6.2892012e-17
+ pclm = 1.5752657
+ vfbsdoff = 0.02
+ phin = 0.15
+ bigsd = 0.00125
+ pkt1 = -4.7748923e-16
+ pkt2 = -1.2933793e-15
+ bigbacc = 0.002588
+ wvoff = 1.1733398e-8
+ paramchk = 1
+ wvsat = -0.0017920539
+ kvth0we = 0.00018
+ wvth0 = -1.9374896e-8
+ tpbswg = 0.0009
+ rbdb = 50
+ pua1 = 1.9082335e-23
+ prwb = 0
+ prwg = 0
+ pub1 = -2.3158905e-32
+ puc1 = -7.9472634e-24
+ waigc = 5.7897385e-11
+ lintnoi = -1.5e-8
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ rdsw = 100
+ ags = 0.36327497
+ lketa = -2.3313752e-8
+ ijthdfwd = 0.01
+ ptvoff = -1.6297696e-16
+ xpart = 1
+ cjd = 0.001357
+ cit = 0.00067194759
+ cjs = 0.001357
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ waigsd = 3.0714895e-12
+ dlc = 1.30529375e-8
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ egidl = 0.29734
+ diomod = 1
+ la0 = -2.5774361e-7
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.017148219
+ pditsd = 0
+ pditsl = 0
+ kt1 = -0.23838945
+ ijthdrev = 0.01
+ lk2 = -9.6280577e-9
+ kt2 = -0.070920535
+ cjswgd = 2.82e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.82e-10
+ llc = -1.18e-13
+ lln = 0.7
+ rshg = 15.6
+ lu0 = -6.2524579e-10
+ mjd = 0.26
+ lua = -9.9655811e-18
+ mjs = 0.26
+ lub = -4.8559819e-26
+ luc = -6.9707629e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 9.4027643e-14
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 2.5483517e-9
+ lpdiblc2 = -2.2782436e-9
+ pbs = 0.52
+ pk2 = 9.5548939e-17
+ pu0 = 8.1677938e-18
+ prt = 0
+ pua = -7.1355685e-24
+ pub = 6.4921301e-33
+ puc = 2.8995668e-24
+ pud = 0
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 8.0998641e-10
+ ub1 = -4.4346517e-19
+ uc1 = 8.2831095e-11
+ mjswgd = 0.85
+ mjswgs = 0.85
+ tpb = 0.0014
+ wa0 = -5.4636242e-7
+ nfactor = 1
+ pvfbsdoff = 0
+ ute = -1
+ wat = -0.018363284
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -5.2787082e-9
+ tcjswg = 0.001
+ wlc = 0
+ wln = 1
+ wu0 = -2.4017748e-10
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -3.8929611e-19
+ wub = -1.8784192e-26
+ wuc = -2.2808063e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ tnom = 25
+ pvoff = -2.0758734e-15
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ cdscb = 0
+ cdscd = 0
+ lkvth0we = -2e-12
+ pvsat = 0
+ wk2we = 5e-12
+ pvth0 = 2.2570293e-15
+ drout = 0.56
+ paigc = -6.3213007e-18
+ nigbacc = 10
+ voffl = 0
+ acnqsmod = 0
+ wags = -2.7824881e-6
+ fprout = 300
+ weta0 = 0
+ wetab = -1.0073378e-8
+ wcit = 5.3579813e-10
+ xrcrg1 = 12
+ xrcrg2 = 1
+ lpclm = -7.0408907e-8
+ voff = -0.13031302
+ rbodymod = 0
+ nigbinv = 10
+ acde = 0.4
+ cgidl = 0.22
+ vsat = 103058.98
+ wtvoff = 3.7639557e-10
+ wint = 0
+ vth0 = 0.42271577
+ wkt1 = -7.3389616e-9
+ wkt2 = 2.2716562e-9
+ wmax = 9e-6
+ wtvfbsdoff = 0
+ aigc = 0.01159193
+ wmin = 9e-7
+ capmod = 2
+ pbswd = 0.8
+ pbsws = 0.8
+ ltvfbsdoff = 0
+ fnoimod = 1
+ wua1 = -5.2698704e-17
+ wub1 = 4.5190152e-26
+ wku0we = 2e-11
+ wuc1 = 3.0855152e-17
+ eigbinv = 1.1
+ wpdiblc2 = 9.3967661e-9
+ bigc = 0.001442
+ mobmod = 0
+ wwlc = 0
+ pdits = 0
+ cigsd = 0.069865
+ cdsc = 0
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ )

.model nch_tt_13 nmos (
+ level = 54
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ lint = 9.7879675e-9
+ bigsd = 0.00125
+ lkt1 = -3.621126e-9
+ lkt2 = -5.6046527e-10
+ lmax = 2.1577e-7
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ lmin = 9e-8
+ wvoff = -2.233608000000001e-9
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ wvsat = -0.00035982647999999954
+ minv = -0.3
+ wvth0 = -5.862617e-9
+ lua1 = 8.0644671e-18
+ lub1 = -5.2760301e-26
+ luc1 = -4.6427809e-18
+ ags = 2.5274682
+ ndep = 1e+18
+ waigc = 3.6164887e-11
+ cjd = 0.001357
+ cit = 0.0010410649
+ cjs = 0.001357
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ lwlc = 0
+ dlc = 1.30529375e-8
+ k3b = 1.9326
+ moin = 5.1
+ lkvth0we = -2e-12
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ nigc = 3.083
+ lketa = -1.0074554e-8
+ xpart = 1
+ la0 = -3.95931149e-8
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.0018760989
+ toxref = 3e-9
+ kt1 = -0.26670569
+ lk2 = -2.2996724e-9
+ kt2 = -0.085875374
+ llc = -1.18e-13
+ lln = 0.7
+ a0 = 0.69883298
+ a1 = 0
+ a2 = 1
+ lu0 = -1.9939706e-10
+ b0 = 0
+ b1 = 0
+ acnqsmod = 0
+ mjd = 0.26
+ lua = 2.3685126e-17
+ mjs = 0.26
+ lub = -3.581049857e-26
+ luc = -1.971816e-18
+ lud = 0
+ at = 80629.42
+ cf = 8.15e-11
+ lwc = 0
+ noff = 2.7195
+ lwl = 0
+ lwn = 1
+ ef = 1.0
+ k1 = 0.274
+ k2 = -0.015489977
+ k3 = -1.8419
+ em = 1000000.0
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ njd = 1.02
+ njs = 1.02
+ nfactor = 1
+ pa0 = 5.1229998e-14
+ egidl = 0.29734
+ ll = -1.18e-13
+ lw = 0
+ u0 = 0.01129738
+ w0 = 0
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 8.2157566e-10
+ pbs = 0.52
+ ua = -2.2820921e-9
+ ub = 2.0823870489000003e-18
+ uc = 4.4751766e-11
+ ud = 0
+ pk2 = 1.6389978e-16
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 6e-9
+ pu0 = -2.2541017e-17
+ prt = 0
+ pua = 6.5907354e-24
+ pub = -1.1536808500000001e-32
+ puc = -4.2264406e-24
+ pud = 0
+ pags = -3.4153056e-19
+ rbodymod = 0
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 6.1728936e-10
+ ub1 = -3.2327621e-19
+ uc1 = 8.8169819e-11
+ ntox = 1
+ pcit = -6.0109378e-17
+ pclm = 1.3619854
+ tpb = 0.0014
+ wa0 = -3.4353242e-7
+ ute = -1
+ wat = -0.010179511
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -5.6026458e-9
+ wlc = 0
+ wln = 1
+ wu0 = -9.4638093e-11
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -6.5442869e-17
+ wub = 6.6660889e-26
+ wuc = 1.0964484e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ ltvoff = 4.8985213e-12
+ phin = 0.15
+ pvfbsdoff = 0
+ nigbacc = 10
+ pkt1 = 2.8243122e-15
+ pkt2 = -3.7226831e-16
+ wpdiblc2 = -7.3538749e-9
+ lku0we = 2.5e-11
+ pvoff = 8.711494700000001e-16
+ rbdb = 50
+ pua1 = -3.4072796e-24
+ prwb = 0
+ prwg = 0
+ pub1 = 3.7649133e-33
+ epsrox = 3.9
+ puc1 = 3.7978198e-24
+ cdscb = 0
+ cdscd = 0
+ rbpb = 50
+ rbpd = 50
+ nigbinv = 10
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ pvsat = -3.0219949000000006e-10
+ wk2we = 5e-12
+ pvth0 = -5.940435999999998e-16
+ rdsw = 100
+ drout = 0.56
+ rdsmod = 0
+ igbmod = 1
+ paigc = -1.7357437e-18
+ voffl = 0
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ pbswgd = 0.95
+ pbswgs = 0.95
+ weta0 = 0
+ wetab = -1.0073378e-8
+ wkvth0we = 2e-12
+ fnoimod = 1
+ lpclm = -2.540677e-8
+ igcmod = 1
+ eigbinv = 1.1
+ rshg = 15.6
+ trnqsmod = 0
+ cgidl = 0.22
+ pbswd = 0.8
+ pbsws = 0.8
+ paigsd = -5.1229584e-23
+ rgatemod = 0
+ tnom = 25
+ cigbacc = 0.32875
+ tnjtsswg = 1
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ permod = 1
+ pdits = 0
+ cigsd = 0.069865
+ tnoimod = 0
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ cigbinv = 0.006
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ wags = 1.2163338e-6
+ voffcv = -0.16942
+ wpemod = 1
+ wcit = 5.2261028e-10
+ tnoia = 0
+ voff = -0.1572150866
+ version = 4.5
+ acde = 0.4
+ tempmod = 0
+ peta0 = 0
+ vsat = 102561.23895
+ wint = 0
+ vth0 = 0.4372123399
+ wketa = 1.0437078e-7
+ wkt1 = -2.298731e-8
+ wkt2 = -2.0937989e-9
+ tpbsw = 0.0019
+ wmax = 9e-6
+ aigc = 0.011522737
+ wmin = 9e-7
+ cjswd = 8.2e-11
+ aigbacc = 0.02
+ cjsws = 8.2e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ wua1 = 5.3887147e-17
+ wub1 = -8.2410881e-26
+ wuc1 = -2.4808749e-17
+ tpbswg = 0.0009
+ bigc = 0.001442
+ wwlc = 0
+ aigbinv = 0.0163
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ ptvoff = 8.9623963e-17
+ ijthsfwd = 0.01
+ scref = 1e-6
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ waigsd = 3.0721194e-12
+ pigcd = 2.621
+ aigsd = 0.010772879
+ diomod = 1
+ lvoff = -4.1479246e-10
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 2.82e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.82e-10
+ lvsat = 0.00010503966000000005
+ tvfbsdoff = 0.022
+ ijthsrev = 0.01
+ lvth0 = -8.000254980000001e-9
+ poxedge = 1
+ delta = 0.007595625
+ laigc = -4.6341008e-12
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ binunit = 2
+ rnoia = 0
+ rnoib = 0
+ mjswgd = 0.85
+ mjswgs = 0.85
+ k2we = 5e-5
+ pketa = -1.2207451e-14
+ tcjswg = 0.001
+ ngate = 8e+20
+ dsub = 0.75
+ ngcon = 1
+ dtox = 2.7e-10
+ wpclm = -2.3899735e-8
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ ppdiblc2 = 7.6111026e-16
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ eta0 = 0.3
+ etab = -0.24888148
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ fprout = 300
+ wtvfbsdoff = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ pkvth0we = -1.3e-19
+ ltvfbsdoff = 0
+ wtvoff = -8.2076521e-10
+ tvoff = 0.00074618122
+ vfbsdoff = 0.02
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ capmod = 2
+ njtsswg = 9
+ wku0we = 2e-11
+ paramchk = 1
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ ku0we = -0.0007
+ mobmod = 0
+ beta0 = 13
+ leta0 = 0
+ ckappad = 0.6
+ ptvfbsdoff = 0
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.022446923
+ pdiblcb = -0.3
+ ppclm = 9.2725546e-15
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ ijthdfwd = 0.01
+ keta = -0.10468292
+ bigbacc = 0.002588
+ laigsd = 3.9592657e-17
+ lags = 3.7696529e-13
+ dmcgt = 0
+ tcjsw = 0.000357
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 9.1265533e-11
+ kvth0we = 0.00018
+ ijthdrev = 0.01
+ kt1l = 0
+ lintnoi = -1.5e-8
+ lpdiblc2 = -1.4676946e-9
+ bigbinv = 0.004953
+ )

.model nch_tt_14 nmos (
+ level = 54
+ poxedge = 1
+ binunit = 2
+ scref = 1e-6
+ toxref = 3e-9
+ pigcd = 2.621
+ aigsd = 0.010772879
+ wags = 1.2163302e-6
+ lvoff = -2.0518068800000008e-9
+ pkvth0we = -1.3e-19
+ wcit = 1.5125736e-10
+ tvfbsdoff = 0.022
+ voff = -0.13980004150000003
+ lvsat = 0.0015075818900000004
+ lvth0 = 2.23756691e-9
+ acde = 0.4
+ delta = 0.007595625
+ vsat = 87640.57610000002
+ laigc = -2.2637509e-11
+ wint = 0
+ vfbsdoff = 0.02
+ vth0 = 0.3282993353
+ ltvoff = 1.2509019e-10
+ wkt1 = 8.3830806e-8
+ wkt2 = 1.6147625e-8
+ rnoia = 0
+ rnoib = 0
+ wmax = 9e-6
+ aigc = 0.011714263
+ wmin = 9e-7
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ pketa = 8.4378567e-15
+ ngate = 8e+20
+ paramchk = 1
+ ngcon = 1
+ wpclm = 3.4675908e-7
+ wua1 = -1.154179e-16
+ wub1 = 3.1505286e-27
+ wuc1 = 9.7519251e-17
+ lku0we = 2.5e-11
+ a0 = -0.035582299999999956
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ bigc = 0.001442
+ gbmin = 1e-12
+ epsrox = 3.9
+ at = 65883.509
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = -0.034587969
+ k3 = -1.8419
+ wvfbsdoff = 0
+ em = 1000000.0
+ wwlc = 0
+ jswgd = 1.28e-13
+ lvfbsdoff = 0
+ jswgs = 1.28e-13
+ ll = 0
+ lw = 0
+ u0 = 0.0078765756
+ w0 = 0
+ ua = -2.421907e-9
+ ub = 1.9130826320999997e-18
+ uc = 4.338735e-12
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 6e-9
+ rdsmod = 0
+ cdsc = 0
+ igbmod = 1
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ ijthdfwd = 0.01
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ pbswgd = 0.95
+ pbswgs = 0.95
+ njtsswg = 9
+ igcmod = 1
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ ijthdrev = 0.01
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.006833075
+ pdiblcb = -0.3
+ tvoff = -0.00053245355
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ lpdiblc2 = 7.1362462e-15
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ k2we = 5e-5
+ paigsd = 1.5255572e-23
+ dsub = 0.75
+ dtox = 2.7e-10
+ ku0we = -0.0007
+ bigbacc = 0.002588
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ beta0 = 13
+ leta0 = 2.6128654e-9
+ letab = -2.2297043e-8
+ permod = 1
+ kvth0we = 0.00018
+ ppclm = -2.5569374e-14
+ eta0 = 0.27220356
+ etab = -0.011678893
+ lkvth0we = -2e-12
+ dlcig = 2.5e-9
+ lintnoi = -1.5e-8
+ bgidl = 2320000000.0
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ acnqsmod = 0
+ voffcv = -0.16942
+ wpemod = 1
+ dmcgt = 0
+ tcjsw = 0.000357
+ rbodymod = 0
+ bigsd = 0.00125
+ ags = 2.5274722
+ wvoff = 8.241506600000007e-9
+ cjd = 0.001357
+ cit = 0.00030181593
+ cjs = 0.001357
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 3.26497e-9
+ tpbswg = 0.0009
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ wvsat = -0.0092125549
+ nfactor = 1
+ wvth0 = -1.3305709099999998e-8
+ wpdiblc2 = 7.4309162e-10
+ waigc = -2.4473999e-12
+ la0 = 2.94419216e-8
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.00048998333
+ kt1 = -0.41803712
+ lk2 = -5.0446112e-10
+ kt2 = -0.10268076
+ llc = 0
+ lln = 1
+ lu0 = 1.2215857e-10
+ mjd = 0.26
+ lua = 3.6827721e-17
+ mjs = 0.26
+ lub = -1.9895881809999996e-26
+ luc = 1.827009e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ ptvoff = -1.5034232e-16
+ njd = 1.02
+ njs = 1.02
+ pa0 = 7.627786000000002e-15
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 9.8787885e-10
+ pbs = 0.52
+ pk2 = 1.6131306e-16
+ waigsd = 3.0714121e-12
+ lketa = 2.8547804e-8
+ pu0 = -1.7406607e-16
+ prt = 0
+ pua = -1.4490045e-23
+ xpart = 1
+ pub = 2.3973370000000036e-34
+ puc = 4.0045874e-24
+ pud = 0
+ rsh = 17.5
+ keta = -0.51555907
+ tcj = 0.00076
+ ua1 = 9.0255397e-10
+ ub1 = -8.0270486e-19
+ uc1 = -7.4218809e-11
+ diomod = 1
+ tpb = 0.0014
+ nigbacc = 10
+ wa0 = 1.203209e-7
+ egidl = 0.29734
+ ute = -1
+ wat = -0.011948694
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -5.5751276e-9
+ pditsd = 0
+ pditsl = 0
+ wlc = 0
+ wln = 1
+ wkvth0we = 2e-12
+ wu0 = 1.5173305e-9
+ cjswgd = 2.82e-10
+ pku0we = -1.5e-18
+ xgl = -1.09e-8
+ cjswgs = 2.82e-10
+ xgw = 0
+ wua = 1.5882075e-16
+ wub = -5.862147e-26
+ wuc = -7.6599643e-17
+ wud = 0
+ wwc = 0
+ jswd = 1.28e-13
+ wwl = 0
+ wwn = 1
+ jsws = 1.28e-13
+ lcit = 1.6075494e-10
+ kt1l = 0
+ trnqsmod = 0
+ nigbinv = 10
+ lint = 0
+ mjswgd = 0.85
+ mjswgs = 0.85
+ lkt1 = 1.0604028e-8
+ lkt2 = 1.0192413e-9
+ pvfbsdoff = 0
+ lmax = 9e-8
+ tcjswg = 0.001
+ lmin = 5.4e-8
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ minv = -0.3
+ rgatemod = 0
+ lua1 = -1.8750406e-17
+ wtvfbsdoff = 0
+ lub1 = -7.6940068e-27
+ luc1 = 1.062175e-17
+ pvoff = -1.135113399999999e-16
+ tnjtsswg = 1
+ fnoimod = 1
+ ndep = 1e+18
+ eigbinv = 1.1
+ cdscb = 0
+ cdscd = 0
+ lwlc = 0
+ moin = 5.1
+ pvsat = 5.299570200000001e-10
+ wk2we = 5e-12
+ pvth0 = 1.0560707800000005e-16
+ ltvfbsdoff = 0
+ drout = 0.56
+ nigc = 3.083
+ paigc = 1.8938113e-18
+ fprout = 300
+ voffl = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ weta0 = -3.9858587e-8
+ wetab = 2.7041872e-8
+ lpclm = -8.5343289e-9
+ wtvoff = 1.7320676e-9
+ cigbacc = 0.32875
+ ntox = 1
+ pcit = -2.5202203e-17
+ pclm = 1.1824913
+ cgidl = 0.22
+ ptvfbsdoff = 0
+ tnoimod = 0
+ phin = 0.15
+ capmod = 2
+ pkt1 = -7.2165907e-15
+ pkt2 = -2.0869621e-15
+ wku0we = 2e-11
+ cigbinv = 0.006
+ pbswd = 0.8
+ pbsws = 0.8
+ mobmod = 0
+ rbdb = 50
+ pua1 = 1.2507395e-23
+ prwb = 0
+ prwg = 0
+ pub1 = -4.2778592e-33
+ puc1 = -7.7010123e-24
+ version = 4.5
+ pdits = 0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ cigsd = 0.069865
+ tempmod = 0
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ rdsw = 100
+ ijthsfwd = 0.01
+ aigbacc = 0.02
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ laigsd = -1.6939346e-18
+ tnoia = 0
+ ijthsrev = 0.01
+ rshg = 15.6
+ peta0 = 3.7467072e-15
+ aigbinv = 0.0163
+ petab = -3.4888335e-15
+ wketa = -1.1526014e-7
+ tpbsw = 0.0019
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ cjswd = 8.2e-11
+ cjsws = 8.2e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ ppdiblc2 = -4.5980291e-21
+ tnom = 25
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ )

.model nch_tt_15 nmos (
+ level = 54
+ fnoimod = 1
+ ltvoff = -2.8596488e-10
+ eigbinv = 1.1
+ pvfbsdoff = 0
+ lku0we = 2.5e-11
+ epsrox = 3.9
+ pvoff = 8.85540199999999e-16
+ cdscb = 0
+ cdscd = 0
+ rdsmod = 0
+ cigbacc = 0.32875
+ pvsat = -2.8119773e-9
+ igbmod = 1
+ wk2we = 5e-12
+ pvth0 = -7.348170000000001e-16
+ drout = 0.56
+ ijthsfwd = 0.01
+ paigc = 1.0773556e-18
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ tnoimod = 0
+ voffl = 0
+ pbswgd = 0.95
+ pbswgs = 0.95
+ keta = 0.067264197
+ cigbinv = 0.006
+ weta0 = 3.2678994e-7
+ igcmod = 1
+ wetab = -1.4667966e-7
+ lpclm = -8.0899178e-8
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 3.2711574e-10
+ ijthsrev = 0.01
+ kt1l = 0
+ cgidl = 0.22
+ version = 4.5
+ a0 = 5.6809619
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = -88751.793
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = -0.014951152
+ k3 = -1.8419
+ em = 1000000.0
+ ll = 0
+ tempmod = 0
+ lw = 0
+ lint = 0
+ u0 = 0.00039525646
+ w0 = 0
+ ua = -3.0786989e-9
+ ub = 2.197681248e-18
+ uc = -5.08518e-12
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 6e-9
+ lkt1 = -1.5973163e-8
+ lkt2 = 1.223943e-9
+ lmax = 5.4e-8
+ lmin = 4.5e-8
+ paigsd = -3.180948e-23
+ pbswd = 0.8
+ lpe0 = 9.2e-8
+ pbsws = 0.8
+ lpeb = 2.5e-7
+ aigbacc = 0.02
+ minv = -0.3
+ permod = 1
+ lua1 = 1.293984e-17
+ lub1 = 3.71094339e-26
+ luc1 = 1.702510023e-17
+ ndep = 1e+18
+ pdits = 0
+ lwlc = 0
+ cigsd = 0.069865
+ moin = 5.1
+ aigbinv = 0.0163
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ nigc = 3.083
+ voffcv = -0.16942
+ wpemod = 1
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ pkvth0we = -1.3e-19
+ tnoia = 0
+ ntox = 1
+ pcit = 7.5457403e-17
+ pclm = 2.4301611
+ peta0 = -1.7518907e-14
+ petab = 6.5870154e-15
+ vfbsdoff = 0.02
+ wketa = 1.9475197e-7
+ poxedge = 1
+ tpbsw = 0.0019
+ phin = 0.15
+ cjswd = 8.2e-11
+ cjsws = 8.2e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ binunit = 2
+ pkt1 = 1.293618e-14
+ pkt2 = 7.7933247e-16
+ tpbswg = 0.0009
+ paramchk = 1
+ rbdb = 50
+ pua1 = -3.7208869e-24
+ prwb = 0
+ prwg = 0
+ pub1 = -6.9156579e-32
+ puc1 = -1.1133321e-23
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ ptvoff = 3.472697e-16
+ waigsd = 3.0722235e-12
+ rdsw = 100
+ ijthdfwd = 0.01
+ scref = 1e-6
+ diomod = 1
+ pigcd = 2.621
+ aigsd = 0.010772879
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ pditsd = 0
+ pditsl = 0
+ lvoff = -3.6979500799999987e-9
+ cjswgd = 2.82e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.82e-10
+ tvfbsdoff = 0.022
+ lvsat = 0.0018704337899999998
+ ijthdrev = 0.01
+ lvth0 = 2.4529352400000003e-9
+ rshg = 15.6
+ delta = 0.007595625
+ laigc = -2.1310273e-11
+ wtvfbsdoff = 0
+ mjswgd = 0.85
+ mjswgs = 0.85
+ rnoia = 0
+ rnoib = 0
+ tcjswg = 0.001
+ ltvfbsdoff = 0
+ pketa = -9.5428465e-15
+ ngate = 8e+20
+ ngcon = 1
+ wpclm = -1.3405624e-6
+ njtsswg = 9
+ tnom = 25
+ wvfbsdoff = 0
+ gbmin = 1e-12
+ lvfbsdoff = 0
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ jswgd = 1.28e-13
+ toxe = 2.43e-9
+ jswgs = 1.28e-13
+ toxm = 2.43e-9
+ ckappad = 0.6
+ lkvth0we = -2e-12
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.0068331981
+ pdiblcb = -0.3
+ fprout = 300
+ ptvfbsdoff = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ acnqsmod = 0
+ wags = 1.2163302e-6
+ wcit = -1.5842531e-9
+ wtvoff = -6.84745e-9
+ bigbacc = 0.002588
+ rbodymod = 0
+ voff = -0.111418263
+ acde = 0.4
+ vsat = 81384.50940000001
+ tvoff = 0.0065547027
+ kvth0we = 0.00018
+ wint = 0
+ vth0 = 0.324586088
+ wkt1 = -2.6363076e-7
+ wkt2 = -3.3271248e-8
+ xjbvd = 1
+ xjbvs = 1
+ wmax = 9e-6
+ lk2we = -1.5e-12
+ capmod = 2
+ aigc = 0.011691379
+ wmin = 9e-7
+ lintnoi = -1.5e-8
+ bigbinv = 0.004953
+ wku0we = 2e-11
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ mobmod = 0
+ ku0we = -0.0007
+ wua1 = 1.6438006e-16
+ wub1 = 1.12174916e-24
+ wuc1 = 1.56696984e-16
+ beta0 = 13
+ wpdiblc2 = 7.4301235e-10
+ leta0 = 1.0110619e-10
+ letab = 3.9727723e-8
+ bigc = 0.001442
+ wwlc = 0
+ ppclm = 7.229527e-14
+ cdsc = 0
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ laigsd = 3.532034e-18
+ dmcgt = 0
+ wkvth0we = 2e-12
+ tcjsw = 0.000357
+ nfactor = 1
+ ags = 2.5274722
+ trnqsmod = 0
+ cjd = 0.001357
+ cit = -0.0025664738
+ cjs = 0.001357
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ dlc = 3.26497e-9
+ k3b = 1.9326
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ bigsd = 0.00125
+ k2we = 5e-5
+ wvoff = -8.983524000000003e-9
+ la0 = -3.0211764e-7
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = 0.0084788642
+ dsub = 0.75
+ kt1 = 0.040190302
+ lk2 = -1.6433965e-9
+ kt2 = -0.1062101
+ dtox = 2.7e-10
+ llc = 0
+ lln = 1
+ lu0 = 5.5607508e-10
+ mjd = 0.26
+ nigbacc = 10
+ lua = 7.492165e-17
+ mjs = 0.26
+ lub = -3.6402602300000003e-26
+ luc = 2.373596e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ wvsat = 0.048407002000000005
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ njd = 1.02
+ njs = 1.02
+ pa0 = -1.230232e-13
+ rgatemod = 0
+ wvth0 = 1.1843679999999776e-9
+ nsd = 1e+20
+ pbd = 0.52
+ pat = -8.1071789e-9
+ pbs = 0.52
+ pk2 = 5.8185614e-16
+ tnjtsswg = 1
+ pu0 = -8.2386575e-17
+ prt = 0
+ pua = 3.4306982e-23
+ pub = -6.0757564e-32
+ puc = -7.1571349e-24
+ pud = 0
+ waigc = 1.1629424e-11
+ eta0 = 0.31550975
+ rsh = 17.5
+ etab = -1.0810714
+ tcj = 0.00076
+ ua1 = 3.5617042e-10
+ ub1 = -1.575178019e-18
+ uc1 = -1.8462139999999999e-10
+ tpb = 0.0014
+ wa0 = 2.372924e-6
+ ute = -1
+ wat = 0.14486265
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -1.282587e-8
+ nigbinv = 10
+ lketa = -5.2559457e-9
+ toxref = 3e-9
+ wlc = 0
+ wln = 1
+ wu0 = -6.3350354e-11
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -6.825073e-16
+ wub = 9.9305604e-25
+ wuc = 1.1584384e-16
+ wud = 0
+ wwc = 0
+ xpart = 1
+ wwl = 0
+ wwn = 1
+ egidl = 0.29734
+ )

.model nch_tt_16 nmos (
+ level = 54
+ pketa = 8.7750313e-15
+ pkt1 = -9.3484796e-16
+ pkt2 = 1.5926682e-15
+ ngate = 8e+20
+ lku0we = 2.5e-11
+ ngcon = 1
+ wpclm = -1.03603352e-6
+ epsrox = 3.9
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ wpdiblc2 = 7.4301235e-10
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ rdsmod = 0
+ bigbacc = 0.002588
+ rbdb = 50
+ pua1 = -1.9060214e-23
+ prwb = 0
+ prwg = 0
+ pub1 = 4.8488331000000005e-32
+ puc1 = 1.47310838e-23
+ igbmod = 1
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ rdsw = 100
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ kvth0we = 0.00018
+ pbswgd = 0.95
+ pbswgs = 0.95
+ lintnoi = -1.5e-8
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ igcmod = 1
+ wkvth0we = 2e-12
+ rshg = 15.6
+ trnqsmod = 0
+ tvoff = 0.002919136
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ paigsd = 4.3875156e-23
+ ku0we = -0.0007
+ permod = 1
+ beta0 = 13
+ rgatemod = 0
+ leta0 = 1.5743207e-8
+ tnom = 25
+ letab = 3.0329695e-8
+ tnjtsswg = 1
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ nfactor = 1
+ ppclm = 5.7373356e-14
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ voffcv = -0.16942
+ wpemod = 1
+ a0 = 3.2177147
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 125884.31
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.025015951
+ k3 = -1.8419
+ em = 1000000.0
+ ll = 0
+ lw = 0
+ ags = 2.5274722
+ u0 = 0.0045836023
+ w0 = 0
+ ua = -2.19661343e-9
+ ub = 1.4860819409999996e-18
+ uc = 2.2595638e-10
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ wags = 1.2163302e-6
+ xl = 4e-9
+ ww = 0
+ xw = 6e-9
+ cjd = 0.001357
+ cit = -0.0023198349
+ cjs = 0.001357
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dmcgt = 0
+ dlc = 3.26497e-9
+ wcit = 1.9973064e-9
+ tcjsw = 0.000357
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ nigbacc = 10
+ voff = -0.04075972859999999
+ acde = 0.4
+ la0 = -1.8141853e-7
+ vsat = 80550.4817
+ wint = 0
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.0020383049
+ vth0 = 0.3550252606
+ kt1 = -0.20813859
+ lk2 = -3.6017846e-9
+ kt2 = -0.11042259
+ llc = 0
+ lln = 1
+ lu0 = 3.5084613e-10
+ wkt1 = 1.9451446e-8
+ wkt2 = -4.9869936e-8
+ mjd = 0.26
+ bigsd = 0.00125
+ lua = 3.1699464000000005e-17
+ mjs = 0.26
+ lub = -1.5342368999999952e-27
+ luc = -8.94744e-18
+ lud = 0
+ wmax = 9e-6
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ aigc = 0.011397597
+ wmin = 9e-7
+ njs = 1.02
+ pa0 = -1.9996651e-13
+ nsd = 1e+20
+ nigbinv = 10
+ pbd = 0.52
+ pat = 1.590101e-10
+ pbs = 0.52
+ pk2 = 3.3250012e-16
+ tpbswg = 0.0009
+ pu0 = -4.1242647e-17
+ prt = 0
+ pua = 2.7971342e-23
+ pub = -4.5926045000000006e-32
+ puc = -7.6781524e-24
+ pud = 0
+ wvoff = 8.333983999999995e-9
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 4.3071269e-10
+ ub1 = -2.19332361e-19
+ uc1 = 5.294111900000001e-10
+ wua1 = 4.7742754e-16
+ tpb = 0.0014
+ wub1 = -1.27916739e-24
+ wuc1 = -3.71148e-16
+ wvsat = 0.044412627999999996
+ wa0 = 3.9431957e-6
+ wvth0 = -3.840119699999998e-8
+ ute = -1
+ wat = -0.023835087
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -7.7369724e-9
+ bigc = 0.001442
+ wlc = 0
+ wln = 1
+ wu0 = -9.0302236e-10
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -5.5320853e-16
+ wub = 6.903720200000001e-25
+ wuc = 1.2647685e-16
+ wud = 0
+ wwlc = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ waigc = -9.3979847e-11
+ ptvoff = -3.4317401e-17
+ waigsd = 3.0706789e-12
+ fnoimod = 1
+ cdsc = 0
+ eigbinv = 1.1
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ lketa = -2.4929909e-8
+ xtis = 3
+ ijthsfwd = 0.01
+ diomod = 1
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ xpart = 1
+ wtvfbsdoff = 0
+ cigc = 0.000625
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 2.82e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.82e-10
+ egidl = 0.29734
+ ltvfbsdoff = 0
+ ijthsrev = 0.01
+ mjswgd = 0.85
+ mjswgs = 0.85
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ cigbacc = 0.32875
+ pvfbsdoff = 0
+ tcjswg = 0.001
+ tnoimod = 0
+ k2we = 5e-5
+ dsub = 0.75
+ dtox = 2.7e-10
+ ptvfbsdoff = 0
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ cigbinv = 0.006
+ pvoff = 3.698261999999959e-17
+ cdscb = 0
+ cdscd = 0
+ eta0 = -0.003716791
+ etab = -0.88927493
+ pvsat = -2.6162530499999997e-9
+ wk2we = 5e-12
+ pvth0 = 1.20487516e-15
+ drout = 0.56
+ version = 4.5
+ fprout = 300
+ paigc = 6.2522098e-18
+ tempmod = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ voffl = 0
+ weta0 = 2.2378028e-8
+ pkvth0we = -1.3e-19
+ wetab = 3.831648e-8
+ aigbacc = 0.02
+ wtvoff = 9.4004181e-10
+ lpclm = -7.043921000000001e-8
+ cgidl = 0.22
+ vfbsdoff = 0.02
+ capmod = 2
+ aigbinv = 0.0163
+ wku0we = 2e-11
+ mobmod = 0
+ pbswd = 0.8
+ pbsws = 0.8
+ paramchk = 1
+ pdits = 0
+ cigsd = 0.069865
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ poxedge = 1
+ ijthdfwd = 0.01
+ laigsd = -2.6649547e-17
+ pk2we = -1e-19
+ keta = 0.46877367
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ binunit = 2
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ tnoia = 0
+ lcit = 3.1503043e-10
+ ijthdrev = 0.01
+ kt1l = 0
+ peta0 = -2.6027237e-15
+ petab = -2.4777955e-15
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ wketa = -1.7908228e-7
+ tpbsw = 0.0019
+ lint = 0
+ cjswd = 8.2e-11
+ cjsws = 8.2e-11
+ lkt1 = -3.805047e-9
+ lkt2 = 1.4303548e-9
+ mjswd = 0.11
+ lmax = 4.5e-8
+ mjsws = 0.11
+ agidl = 9.41e-8
+ lmin = 3.6e-8
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ minv = -0.3
+ lua1 = 9.2872684e-18
+ lub1 = -2.93270018e-26
+ luc1 = -1.796249619e-17
+ ndep = 1e+18
+ lwlc = 0
+ lkvth0we = -2e-12
+ moin = 5.1
+ toxref = 3e-9
+ nigc = 3.083
+ scref = 1e-6
+ pigcd = 2.621
+ aigsd = 0.01077288
+ acnqsmod = 0
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ lvoff = -7.160218279999998e-9
+ tvfbsdoff = 0.022
+ njtsswg = 9
+ rbodymod = 0
+ lvsat = 0.001911301613
+ lvth0 = 9.6141603e-10
+ ntox = 1
+ ltvoff = -1.0782211e-10
+ pcit = -1.0003901e-16
+ pclm = 2.21669238
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ delta = 0.007595625
+ laigc = -6.9149623e-12
+ ckappad = 0.6
+ ckappas = 0.6
+ rnoia = 0
+ rnoib = 0
+ pdiblc1 = 0
+ pdiblc2 = 0.0068331981
+ phin = 0.15
+ pdiblcb = -0.3
+ )

.model nch_tt_17 nmos (
+ level = 54
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ pbswgd = 0.95
+ xtis = 3
+ pbswgs = 0.95
+ ijthdfwd = 0.01
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ aigbinv = 0.0163
+ cigc = 0.000625
+ voffl = 0
+ igcmod = 1
+ weta0 = -1.09928e-7
+ wetab = 2.7482e-8
+ ijthdrev = 0.01
+ cgidl = 0.22
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ poxedge = 1
+ k2we = 5e-5
+ pbswd = 0.8
+ pbsws = 0.8
+ dsub = 0.75
+ permod = 1
+ dtox = 2.7e-10
+ binunit = 2
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ pdits = 0
+ eta0 = 0.42133333
+ cigsd = 0.069865
+ etab = -0.29033333
+ lkvth0we = -2e-12
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ voffcv = -0.16942
+ wpemod = 1
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ acnqsmod = 0
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ tnoia = 0
+ rbodymod = 0
+ peta0 = 0
+ wketa = -3.7974654e-8
+ tpbsw = 0.0019
+ cjswd = 8.2e-11
+ tpbswg = 0.0009
+ cjsws = 8.2e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ wtvfbsdoff = 0
+ a0 = 2.2098167
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 72000
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.016686228
+ k3 = -1.8419
+ em = 1000000.0
+ wpdiblc2 = -6.449088e-9
+ ll = 0
+ lw = 0
+ u0 = 0.0155465
+ w0 = 0
+ ua = -1.7855187e-9
+ ub = 2.0636167e-18
+ uc = 7.8391667e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ptvoff = 0
+ ww = 0
+ xw = 6e-9
+ njtsswg = 9
+ ltvfbsdoff = 0
+ waigsd = 3.0876027e-12
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ diomod = 1
+ scref = 1e-6
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.025656394
+ pigcd = 2.621
+ pdiblcb = -0.3
+ pditsd = 0
+ pditsl = 0
+ aigsd = 0.010772862
+ cjswgd = 2.82e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.82e-10
+ keta = 0.015093331
+ tvfbsdoff = 0.022
+ lvoff = 0
+ wkvth0we = 2e-12
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lvsat = 0
+ lcit = 0
+ lvth0 = 0
+ ptvfbsdoff = 0
+ kt1l = 0
+ mjswgd = 0.85
+ mjswgs = 0.85
+ trnqsmod = 0
+ delta = 0.007595625
+ bigbacc = 0.002588
+ tcjswg = 0.001
+ rnoia = 0
+ rnoib = 0
+ lint = 6.5375218e-9
+ kvth0we = 0.00018
+ lkt1 = 0
+ lmax = 2.001e-5
+ lmin = 8.9991e-6
+ ngate = 8e+20
+ lintnoi = -1.5e-8
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ ngcon = 1
+ bigbinv = 0.004953
+ wpclm = 5.7423639e-7
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ rgatemod = 0
+ minv = -0.3
+ lub1 = 0
+ gbmin = 1e-12
+ tnjtsswg = 1
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ ndep = 1e+18
+ lwlc = 0
+ moin = 5.1
+ fprout = 300
+ nigc = 3.083
+ xrcrg1 = 12
+ xrcrg2 = 1
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ wtvoff = 9.3503662e-10
+ ntox = 1
+ pcit = 0
+ pclm = 0.629885
+ tvoff = 5.0359625e-5
+ capmod = 2
+ nfactor = 1
+ wku0we = 2e-11
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ phin = 0.15
+ mobmod = 0
+ pkt1 = 0
+ ku0we = -0.0007
+ beta0 = 13
+ leta0 = 0
+ nigbacc = 10
+ rbdb = 50
+ prwb = 0
+ prwg = 0
+ pub1 = 0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ ags = 0.65720097
+ dlcig = 2.5e-9
+ rdsw = 100
+ bgidl = 2320000000.0
+ cjd = 0.001357
+ cit = 6.2896875e-5
+ cjs = 0.001357
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 9.8024918e-9
+ ijthsfwd = 0.01
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ nigbinv = 10
+ la0 = 0
+ jsd = 6.11e-7
+ dmcgt = 0
+ jss = 6.11e-7
+ lat = 0
+ kt1 = -0.28314411
+ kt2 = -0.074391698
+ tcjsw = 0.000357
+ llc = 0
+ lln = 1
+ lu0 = 0
+ mjd = 0.26
+ mjs = 0.26
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 0
+ ijthsrev = 0.01
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 0
+ pbs = 0.52
+ rshg = 15.6
+ pu0 = 0
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ prt = 0
+ pud = 0
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = -6.8749055e-10
+ ub1 = 1.0341951e-18
+ uc1 = 4.5339833e-11
+ fnoimod = 1
+ bigsd = 0.00125
+ tpb = 0.0014
+ wa0 = 7.159061e-7
+ eigbinv = 1.1
+ ute = -2.01925
+ wat = 0
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 3.760485e-9
+ wlc = 0
+ wln = 1
+ wu0 = -1.23669e-10
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -7.132277e-17
+ wub = 7.28273e-26
+ wuc = -1.167985e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ wvoff = 1.0181215e-9
+ wvsat = -0.0045771271
+ wvth0 = -8.7727395e-9
+ tnom = 25
+ toxe = 2.43e-9
+ waigc = 5.0140497e-11
+ toxm = 2.43e-9
+ toxref = 3e-9
+ cigbacc = 0.32875
+ xpart = 1
+ tnoimod = 0
+ wags = 1.1493247e-7
+ egidl = 0.29734
+ pkvth0we = -1.3e-19
+ wcit = 4.4907306e-10
+ cigbinv = 0.006
+ voff = -0.11158375
+ ltvoff = 0
+ acde = 0.4
+ vsat = 106133.02
+ vfbsdoff = 0.02
+ wint = 0
+ pvfbsdoff = 0
+ vth0 = 0.34772953
+ wkt1 = 3.4075481e-8
+ wkt2 = 1.5939759e-8
+ wmax = 9e-7
+ aigc = 0.011740211
+ wmin = 5.4e-7
+ version = 4.5
+ tempmod = 0
+ lku0we = 2.5e-11
+ epsrox = 3.9
+ paramchk = 1
+ wua1 = 1.0731531e-15
+ wub1 = -9.2968455e-25
+ wuc1 = -1.4414309e-17
+ aigbacc = 0.02
+ rdsmod = 0
+ bigc = 0.001442
+ pvoff = 0
+ wute = 5.565105e-7
+ wwlc = 0
+ igbmod = 1
+ cdscb = 0
+ cdscd = 0
+ pvsat = 0
+ wk2we = 5e-12
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ pvth0 = 0
+ cdsc = 0
+ drout = 0.56
+ )

.model nch_tt_18 nmos (
+ level = 54
+ kt1l = 0
+ nigbacc = 10
+ tvoff = -0.0002433276
+ paigsd = 1.3573222e-22
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ lint = 6.5375218e-9
+ lkt1 = 8.6246405e-8
+ lkt2 = 5.1456509e-9
+ lmax = 8.9991e-6
+ lmin = 8.9908e-7
+ permod = 1
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ nigbinv = 10
+ ags = 0.61161289
+ ku0we = -0.0007
+ ppdiblc2 = 1.9760389e-14
+ beta0 = 13
+ cjd = 0.001357
+ leta0 = 0
+ cit = -0.00011782923
+ cjs = 0.001357
+ minv = -0.3
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ lua1 = 1.38467e-15
+ lub1 = -1.4892591e-24
+ luc1 = 1.0686128e-16
+ dlc = 9.8024918e-9
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ ndep = 1e+18
+ lute = 1.0068051e-6
+ lwlc = 0
+ moin = 5.1
+ dlcig = 2.5e-9
+ voffcv = -0.16942
+ wpemod = 1
+ bgidl = 2320000000.0
+ la0 = -1.1479603e-6
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ nigc = 3.083
+ lat = 0.085345067
+ kt1 = -0.2927377
+ lk2 = -1.3507419e-8
+ kt2 = -0.074964073
+ llc = 0
+ lln = 1
+ lu0 = -2.0004396e-9
+ fnoimod = 1
+ mjd = 0.26
+ lua = -1.5028094e-16
+ mjs = 0.26
+ lub = -1.4426347e-25
+ luc = -5.2935673e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = -5.1713984e-13
+ eigbinv = 1.1
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 0
+ pbs = 0.52
+ pk2 = -1.6553107e-15
+ pu0 = 1.3573224e-17
+ prt = 0
+ noff = 2.7195
+ pua = -3.5916841e-23
+ pub = 6.5823852e-32
+ puc = 3.1761344e-23
+ pud = 0
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ pkvth0we = -1.3e-19
+ dmcgt = 0
+ rsh = 17.5
+ tcjsw = 0.000357
+ tcj = 0.00076
+ ua1 = -8.4151391e-10
+ ub1 = 1.1998524e-18
+ uc1 = 3.3453151e-11
+ tpb = 0.0014
+ wa0 = 7.7343e-7
+ pags = -1.4569295e-13
+ ute = -2.1312417
+ wtvfbsdoff = 0
+ wat = 0
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 3.944613e-9
+ wlc = 0
+ wln = 1
+ ntox = 1
+ wu0 = -1.2517881e-10
+ pcit = -6.2947523e-16
+ xgl = -1.09e-8
+ pclm = 0.629885
+ xgw = 0
+ wua = -6.7327571e-17
+ wub = 6.5505403e-26
+ wuc = -1.5212814e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ vfbsdoff = 0.02
+ tpbswg = 0.0009
+ bigsd = 0.00125
+ ltvfbsdoff = 0
+ phin = 0.15
+ cigbacc = 0.32875
+ wvoff = 8.2208115e-10
+ pkt1 = -6.952314e-14
+ pkt2 = -1.5079533e-14
+ paramchk = 1
+ tnoimod = 0
+ wvsat = -0.0045771271
+ wvth0 = -9.0760901e-9
+ ptvoff = -2.0299898e-15
+ waigsd = 3.0875876e-12
+ waigc = 5.030718e-11
+ rbdb = 50
+ pua1 = -1.044071e-21
+ prwb = 0
+ prwg = 0
+ pub1 = 9.8799081e-31
+ cigbinv = 0.006
+ puc1 = -4.3746501e-23
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ pute = -5.4971558e-13
+ diomod = 1
+ rdsw = 100
+ ptvfbsdoff = 0
+ lketa = -1.3350472e-7
+ ijthdfwd = 0.01
+ pditsd = 0
+ xpart = 1
+ pditsl = 0
+ cjswgd = 2.82e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.82e-10
+ version = 4.5
+ tempmod = 0
+ egidl = 0.29734
+ mjswgd = 0.85
+ mjswgs = 0.85
+ ijthdrev = 0.01
+ aigbacc = 0.02
+ a0 = 2.3375097
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ rshg = 15.6
+ at = 62506.667
+ cf = 8.15e-11
+ tcjswg = 0.001
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.018188722
+ k3 = -1.8419
+ em = 1000000.0
+ pvfbsdoff = 0
+ ll = 0
+ lw = 0
+ u0 = 0.015769018
+ lpdiblc2 = -2.2119558e-8
+ w0 = 0
+ ua = -1.7688022e-9
+ ub = 2.0796638e-18
+ uc = 8.4279951e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 6e-9
+ aigbinv = 0.0163
+ tnom = 25
+ pvoff = 1.7624031e-15
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ cdscb = 0
+ cdscd = 0
+ fprout = 300
+ pvsat = 0
+ lkvth0we = -2e-12
+ wk2we = 5e-12
+ pvth0 = 2.7271227e-15
+ drout = 0.56
+ xrcrg1 = 12
+ xrcrg2 = 1
+ paigc = -1.4984839e-18
+ voffl = 0
+ poxedge = 1
+ acnqsmod = 0
+ wtvoff = 1.1608419e-9
+ wags = 1.3113859e-7
+ weta0 = -1.09928e-7
+ wetab = 2.7482e-8
+ wcit = 5.1909255e-10
+ binunit = 2
+ rbodymod = 0
+ voff = -0.1094379
+ acde = 0.4
+ capmod = 2
+ cgidl = 0.22
+ vsat = 106133.02
+ wint = 0
+ wku0we = 2e-11
+ vth0 = 0.34194059
+ wkt1 = 4.1808867e-8
+ wkt2 = 1.7617127e-8
+ wmax = 9e-7
+ mobmod = 0
+ aigc = 0.011757817
+ wmin = 5.4e-7
+ pbswd = 0.8
+ pbsws = 0.8
+ wua1 = 1.1892901e-15
+ wub1 = -1.0395834e-24
+ wuc1 = -9.5481798e-18
+ wpdiblc2 = -8.647129e-9
+ bigc = 0.001442
+ wute = 6.1765795e-7
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ wwlc = 0
+ pdits = 0
+ cigsd = 0.069865
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ laigsd = -2.4859383e-16
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ wkvth0we = 2e-12
+ tnoia = 0
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ trnqsmod = 0
+ peta0 = 0
+ njtsswg = 9
+ wketa = -4.7550208e-8
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ tpbsw = 0.0019
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ cjswd = 8.2e-11
+ cjsws = 8.2e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.028116857
+ k2we = 5e-5
+ pdiblcb = -0.3
+ dsub = 0.75
+ dtox = 2.7e-10
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ rgatemod = 0
+ tnjtsswg = 1
+ toxref = 3e-9
+ eta0 = 0.42133333
+ etab = -0.29033333
+ bigbacc = 0.002588
+ scref = 1e-6
+ pigcd = 2.621
+ aigsd = 0.010772862
+ kvth0we = 0.00018
+ tvfbsdoff = 0.022
+ lvoff = -1.9291251e-8
+ lintnoi = -1.5e-8
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ ltvoff = 2.6402481e-9
+ lvsat = 0
+ lvth0 = 5.2042566e-8
+ delta = 0.007595625
+ laigc = -1.5827875e-10
+ rnoia = 0
+ rnoib = 0
+ lku0we = 2.5e-11
+ pketa = 8.6084224e-14
+ epsrox = 3.9
+ ngate = 8e+20
+ ngcon = 1
+ wvfbsdoff = 0
+ wpclm = 5.7423639e-7
+ lvfbsdoff = 0
+ rdsmod = 0
+ gbmin = 1e-12
+ igbmod = 1
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ pbswgd = 0.95
+ pbswgs = 0.95
+ nfactor = 1
+ ijthsfwd = 0.01
+ igcmod = 1
+ keta = 0.029943688
+ lags = 4.0983681e-7
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 1.6247277e-9
+ ijthsrev = 0.01
+ )

.model nch_tt_19 nmos (
+ level = 54
+ rgatemod = 0
+ tnom = 25
+ tnjtsswg = 1
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ pdits = 0
+ cigsd = 0.069865
+ voffcv = -0.16942
+ wpemod = 1
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ njtsswg = 9
+ wtvfbsdoff = 0
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ ltvfbsdoff = 0
+ ckappad = 0.6
+ ckappas = 0.6
+ wags = -7.83542e-7
+ pdiblc1 = 0
+ pdiblc2 = -0.019237439
+ pdiblcb = -0.3
+ wcit = -4.5548514e-10
+ tnoia = 0
+ voff = -0.12566406
+ acde = 0.4
+ peta0 = 0
+ vsat = 106133.02
+ wketa = 9.2259042e-8
+ wint = 0
+ tpbswg = 0.0009
+ vth0 = 0.40014179
+ tpbsw = 0.0019
+ wkt1 = -6.9953249e-8
+ wkt2 = 3.7202325e-9
+ wmax = 9e-7
+ bigbacc = 0.002588
+ cjswd = 8.2e-11
+ aigc = 0.01160027
+ cjsws = 8.2e-11
+ wmin = 5.4e-7
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ ptvfbsdoff = 0
+ kvth0we = 0.00018
+ ptvoff = 9.96032e-16
+ wua1 = 1.1798319e-17
+ wub1 = 1.8760115e-25
+ wuc1 = -8.2926019e-17
+ lintnoi = -1.5e-8
+ waigsd = 3.0878745e-12
+ bigbinv = 0.004953
+ bigc = 0.001442
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ wwlc = 0
+ diomod = 1
+ cdsc = 0
+ cgbo = 0
+ pditsd = 0
+ pditsl = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ cjswgd = 2.82e-10
+ ijthsfwd = 0.01
+ scref = 1e-6
+ pku0we = -1.5e-18
+ cjswgs = 2.82e-10
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ pigcd = 2.621
+ tvfbsdoff = 0.022
+ aigsd = 0.010772861
+ lvoff = -4.8499703e-9
+ mjswgd = 0.85
+ mjswgs = 0.85
+ lvsat = 0
+ lvth0 = 2.434924e-10
+ ijthsrev = 0.01
+ tcjswg = 0.001
+ delta = 0.007595625
+ laigc = -1.8062176e-11
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ rnoia = 0
+ rnoib = 0
+ nfactor = 1
+ pketa = -3.8346008e-14
+ ngate = 8e+20
+ k2we = 5e-5
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ ngcon = 1
+ dsub = 0.75
+ wpclm = 5.7423639e-7
+ dtox = 2.7e-10
+ ppdiblc2 = -1.3176269e-14
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ fprout = 300
+ eta0 = 0.42133333
+ etab = -0.29033333
+ xrcrg1 = 12
+ xrcrg2 = 1
+ nigbacc = 10
+ a0 = 1.6362276
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 209176.65
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.014938798
+ k3 = -1.8419
+ em = 1000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.015247274
+ w0 = 0
+ ua = -1.7708735e-9
+ ub = 1.8600147e-18
+ uc = 2.580063e-11
+ ud = 0
+ wtvoff = -2.2391826e-9
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 6e-9
+ pkvth0we = -1.3e-19
+ nigbinv = 10
+ capmod = 2
+ wku0we = 2e-11
+ tvoff = 0.004406442
+ vfbsdoff = 0.02
+ mobmod = 0
+ ags = 2.477561
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ cjd = 0.001357
+ cit = 0.0020125208
+ cjs = 0.001357
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 9.8024918e-9
+ k3b = 1.9326
+ fnoimod = 1
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ eigbinv = 1.1
+ paramchk = 1
+ ku0we = -0.0007
+ beta0 = 13
+ la0 = -5.2381924e-7
+ leta0 = 0
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.04519122
+ kt1 = -0.12585017
+ lk2 = -1.0614987e-8
+ kt2 = -0.061139846
+ llc = 0
+ lln = 1
+ lu0 = -1.5360873e-9
+ mjd = 0.26
+ lua = -1.4843753e-16
+ mjs = 0.26
+ lub = 5.1224193e-26
+ luc = -8.8907704e-19
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 9.5948774e-14
+ nsd = 1e+20
+ pbd = 0.52
+ pat = -4.974413e-9
+ pbs = 0.52
+ laigsd = 2.1900591e-16
+ pk2 = -1.0578878e-15
+ pu0 = 1.1957724e-17
+ dlcig = 2.5e-9
+ prt = 0
+ pua = 5.0063903e-23
+ pub = -8.0709098e-32
+ puc = -9.2074471e-24
+ pud = 0
+ bgidl = 2320000000.0
+ ijthdfwd = 0.01
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 7.2552224e-10
+ ub1 = -4.8701436e-19
+ uc1 = 1.8003493e-10
+ tpb = 0.0014
+ wa0 = 8.4566389e-8
+ ute = -1
+ wat = 0.0055892281
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 3.2733514e-9
+ keta = -0.17327473
+ cigbacc = 0.32875
+ wlc = 0
+ wln = 1
+ wu0 = -1.2336364e-10
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -1.6393515e-16
+ wub = 2.3014917e-25
+ wuc = 3.0819536e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ dmcgt = 0
+ tcjsw = 0.000357
+ lags = -1.250857e-6
+ tnoimod = 0
+ jswd = 1.28e-13
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ jsws = 1.28e-13
+ lcit = -2.712838e-10
+ ijthdrev = 0.01
+ kt1l = 0
+ cigbinv = 0.006
+ lpdiblc2 = 2.0025765e-8
+ bigsd = 0.00125
+ lint = 6.5375218e-9
+ lkt1 = -6.2283496e-8
+ lkt2 = -7.1579117e-9
+ lmax = 8.9908e-7
+ lmin = 4.4908e-7
+ wvoff = 5.2999378e-9
+ lpe0 = 9.2e-8
+ version = 4.5
+ lpeb = 2.5e-7
+ tempmod = 0
+ wvsat = -0.0045771271
+ wvth0 = -7.5199227e-9
+ minv = -0.3
+ lua1 = -9.9922063e-18
+ lub1 = 1.2052288e-26
+ luc1 = -2.3596511e-17
+ toxref = 3e-9
+ waigc = 6.3350032e-11
+ ndep = 1e+18
+ aigbacc = 0.02
+ lwlc = 0
+ lkvth0we = -2e-12
+ moin = 5.1
+ lketa = 4.735968e-8
+ nigc = 3.083
+ xpart = 1
+ acnqsmod = 0
+ aigbinv = 0.0163
+ egidl = 0.29734
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ ltvoff = -1.4980468e-9
+ rbodymod = 0
+ pags = 6.6837277e-13
+ ntox = 1
+ pvfbsdoff = 0
+ pcit = 2.3789891e-16
+ pclm = 0.629885
+ phin = 0.15
+ lku0we = 2.5e-11
+ epsrox = 3.9
+ pkt1 = 2.9945144e-14
+ pkt2 = -2.7112972e-15
+ poxedge = 1
+ rdsmod = 0
+ igbmod = 1
+ wpdiblc2 = 2.8360352e-8
+ pvoff = -2.2228894e-15
+ binunit = 2
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ rbdb = 50
+ pua1 = 3.8966634e-24
+ prwb = 0
+ prwg = 0
+ pub1 = -1.0420346e-31
+ cdscb = 0
+ cdscd = 0
+ puc1 = 2.1559776e-23
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ pvsat = 0
+ rbsb = 50
+ pvag = 1.2
+ pbswgd = 0.95
+ pbswgs = 0.95
+ wk2we = 5e-12
+ pvth0 = 1.3421337e-15
+ drout = 0.56
+ rdsw = 100
+ igcmod = 1
+ paigc = -1.3106622e-17
+ voffl = 0
+ weta0 = -1.09928e-7
+ wetab = 2.7482e-8
+ wkvth0we = 2e-12
+ trnqsmod = 0
+ cgidl = 0.22
+ rshg = 15.6
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ paigsd = -1.1957726e-22
+ permod = 1
+ pbswd = 0.8
+ pbsws = 0.8
+ )

.model nch_tt_20 nmos (
+ level = 54
+ rgatemod = 0
+ tnom = 25
+ tnjtsswg = 1
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ pdits = 0
+ cigsd = 0.069865
+ voffcv = -0.16942
+ wpemod = 1
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ njtsswg = 9
+ wtvfbsdoff = 0
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ ltvfbsdoff = 0
+ ckappad = 0.6
+ ckappas = 0.6
+ wags = 2.514663e-6
+ pdiblc1 = 0
+ pdiblc2 = 0.041730695
+ pdiblcb = -0.3
+ wcit = 1.5646633e-10
+ tnoia = 0
+ voff = -0.11119538
+ acde = 0.4
+ peta0 = 0
+ vsat = 99029.765
+ wketa = 8.4379468e-9
+ wint = 0
+ tpbswg = 0.0009
+ vth0 = 0.40849989
+ tpbsw = 0.0019
+ wkt1 = 1.0316763e-8
+ wkt2 = -6.4493333e-9
+ wmax = 9e-7
+ bigbacc = 0.002588
+ cjswd = 8.2e-11
+ aigc = 0.011620363
+ cjsws = 8.2e-11
+ wmin = 5.4e-7
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ ptvfbsdoff = 0
+ kvth0we = 0.00018
+ ptvoff = -1.0913215e-16
+ wua1 = 2.6150731e-17
+ wub1 = -7.4432483e-26
+ wuc1 = -3.5091334e-17
+ lintnoi = -1.5e-8
+ waigsd = 3.0877293e-12
+ bigbinv = 0.004953
+ bigc = 0.001442
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ wwlc = 0
+ diomod = 1
+ cdsc = 0
+ cgbo = 0
+ pditsd = 0
+ pditsl = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ cjswgd = 2.82e-10
+ ijthsfwd = 0.01
+ scref = 1e-6
+ pku0we = -1.5e-18
+ cjswgs = 2.82e-10
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ pigcd = 2.621
+ tvfbsdoff = 0.022
+ aigsd = 0.010772861
+ lvoff = -1.121619e-8
+ mjswgd = 0.85
+ mjswgs = 0.85
+ lvsat = 0.0031254309
+ lvth0 = -3.434068e-9
+ ijthsrev = 0.01
+ tcjswg = 0.001
+ delta = 0.007595625
+ laigc = -2.6902885e-11
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ rnoia = 0
+ rnoib = 0
+ nfactor = 1
+ pketa = -1.4647263e-15
+ ngate = 8e+20
+ k2we = 5e-5
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ ngcon = 1
+ dsub = 0.75
+ wpclm = 5.7423639e-7
+ dtox = 2.7e-10
+ ppdiblc2 = 1.3236303e-15
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ fprout = 300
+ eta0 = 0.42133333
+ etab = -0.29033333
+ xrcrg1 = 12
+ xrcrg2 = 1
+ nigbacc = 10
+ a0 = -0.63009793
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 152816.98
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.01390817
+ k3 = -1.8419
+ em = 1000000.0
+ ll = -1.18e-13
+ lw = 0
+ u0 = 0.013170665
+ w0 = 0
+ ua = -2.0345741e-9
+ ub = 2.0265059e-18
+ uc = 2.0750138e-11
+ ud = 0
+ wtvoff = 2.7255415e-10
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 6e-9
+ pkvth0we = -1.3e-19
+ nigbinv = 10
+ capmod = 2
+ wku0we = 2e-11
+ tvoff = 0.001369836
+ vfbsdoff = 0.02
+ mobmod = 0
+ ags = -5.4834702
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ cjd = 0.001357
+ cit = 0.0010906361
+ cjs = 0.001357
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 1.30529375e-8
+ k3b = 1.9326
+ fnoimod = 1
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ eigbinv = 1.1
+ paramchk = 1
+ ku0we = -0.0007
+ beta0 = 13
+ la0 = 4.73364e-7
+ leta0 = 0
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.020392964
+ kt1 = -0.257877
+ lk2 = -1.0161511e-8
+ kt2 = -0.061294719
+ llc = -1.18e-13
+ lln = 0.7
+ lu0 = -6.2237936e-10
+ mjd = 0.26
+ lua = -3.2409276e-17
+ mjs = 0.26
+ lub = -2.2031936e-26
+ luc = 1.3331392e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = -5.6835585e-13
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 5.4880901e-9
+ pbs = 0.52
+ laigsd = 6.148791e-17
+ pk2 = 5.7885716e-16
+ pu0 = 5.5708054e-18
+ dlcig = 2.5e-9
+ prt = 0
+ pua = 1.3198419e-23
+ pub = -1.7542132e-32
+ puc = -4.6237685e-24
+ pud = 0
+ bgidl = 2320000000.0
+ ijthdfwd = 0.01
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 7.2295613e-10
+ ub1 = -3.1143135e-19
+ uc1 = 1.5561971e-10
+ tpb = 0.0014
+ wa0 = 1.5943496e-6
+ ute = -1
+ wat = -0.018189188
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -4.4652352e-10
+ keta = -0.031454297
+ cigbacc = 0.32875
+ wlc = 0
+ wln = 1
+ wu0 = -1.0884792e-10
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -8.0149958e-17
+ wub = 8.6587882e-26
+ wuc = 2.0402085e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ dmcgt = 0
+ tcjsw = 0.000357
+ lags = 2.2519967e-6
+ tnoimod = 0
+ jswd = 1.28e-13
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ jsws = 1.28e-13
+ lcit = 1.3434545e-10
+ ijthdrev = 0.01
+ kt1l = 0
+ cigbinv = 0.006
+ lpdiblc2 = -6.8002141e-9
+ bigsd = 0.00125
+ lint = 9.7879675e-9
+ lkt1 = -4.1916909e-9
+ lkt2 = -7.0897675e-9
+ lmax = 4.4908e-7
+ lmin = 2.1577e-7
+ wvoff = -5.5871857e-9
+ lpe0 = 9.2e-8
+ version = 4.5
+ lpeb = 2.5e-7
+ tempmod = 0
+ wvsat = 0.0018584193
+ wvth0 = -6.4953081e-9
+ minv = -0.3
+ lua1 = -8.8631172e-18
+ lub1 = -6.5204234e-26
+ luc1 = -1.2853813e-17
+ toxref = 3e-9
+ waigc = 3.2137522e-11
+ ndep = 1e+18
+ aigbacc = 0.02
+ lwlc = 0
+ lkvth0we = -2e-12
+ moin = 5.1
+ lketa = -1.5041313e-8
+ nigc = 3.083
+ xpart = 1
+ acnqsmod = 0
+ aigbinv = 0.0163
+ egidl = 0.29734
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ ltvoff = -1.6194017e-10
+ rbodymod = 0
+ pags = -7.8283743e-13
+ ntox = 1
+ pvfbsdoff = 0
+ pcit = -3.1359735e-17
+ pclm = 0.629885
+ phin = 0.15
+ lku0we = 2.5e-11
+ epsrox = 3.9
+ pkt1 = -5.3736613e-15
+ pkt2 = 1.7633117e-15
+ poxedge = 1
+ rdsmod = 0
+ igbmod = 1
+ wpdiblc2 = -4.5939646e-9
+ pvoff = 2.567445e-15
+ binunit = 2
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ rbdb = 50
+ pua1 = -2.4183981e-24
+ prwb = 0
+ prwg = 0
+ pub1 = 1.1091342e-32
+ cdscb = 0
+ cdscd = 0
+ puc1 = 5.125141e-25
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ pvsat = -2.8316404e-9
+ rbsb = 50
+ pvag = 1.2
+ pbswgd = 0.95
+ pbswgs = 0.95
+ wk2we = 5e-12
+ pvth0 = 8.9130324e-16
+ drout = 0.56
+ rdsw = 100
+ igcmod = 1
+ paigc = 6.2688273e-19
+ voffl = 0
+ weta0 = -1.09928e-7
+ wetab = 2.7482e-8
+ wkvth0we = 2e-12
+ trnqsmod = 0
+ cgidl = 0.22
+ rshg = 15.6
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ paigsd = -5.5708045e-23
+ permod = 1
+ pbswd = 0.8
+ pbsws = 0.8
+ )

.model nch_tt_21 nmos (
+ level = 54
+ acnqsmod = 0
+ dmcgt = 0
+ version = 4.5
+ tcjsw = 0.000357
+ ptvfbsdoff = 0
+ tempmod = 0
+ rbodymod = 0
+ tpbswg = 0.0009
+ aigbacc = 0.02
+ bigsd = 0.00125
+ wvoff = 4.2089489999999885e-10
+ ptvoff = 6.7086074e-18
+ wvsat = -0.0116031636
+ waigsd = 3.0872445e-12
+ aigbinv = 0.0163
+ wvth0 = 8.290214590000001e-9
+ wpdiblc2 = 3.4958017e-9
+ waigc = 1.7847398e-12
+ diomod = 1
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 2.82e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.82e-10
+ lketa = -3.6124213e-8
+ xpart = 1
+ keta = 0.068466797
+ egidl = 0.29734
+ mjswgd = 0.85
+ mjswgs = 0.85
+ wkvth0we = 2e-12
+ poxedge = 1
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ tcjswg = 0.001
+ lcit = 6.1521194e-11
+ pvfbsdoff = 0
+ kt1l = 0
+ trnqsmod = 0
+ binunit = 2
+ lint = 9.7879675e-9
+ lkt1 = 7.1588252e-10
+ lkt2 = 9.4878496e-10
+ lmax = 2.1577e-7
+ lmin = 9e-8
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ rgatemod = 0
+ minv = -0.3
+ lua1 = 1.428412e-17
+ pvoff = 1.2997136100000001e-15
+ lub1 = -6.3260104e-26
+ luc1 = -5.9196014e-18
+ tnjtsswg = 1
+ fprout = 300
+ ndep = 1e+18
+ cdscb = 0
+ cdscd = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ pvsat = 8.752865999999776e-12
+ lwlc = 0
+ wk2we = 5e-12
+ pvth0 = -2.22841744e-15
+ moin = 5.1
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ drout = 0.56
+ nigc = 3.083
+ paigc = 7.0313197e-18
+ wtvoff = -2.7645419e-10
+ voffl = 0
+ noff = 2.7195
+ weta0 = -1.09928e-7
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ wetab = 2.7482e-8
+ lpclm = 5.9671804e-8
+ capmod = 2
+ wku0we = 2e-11
+ ntox = 1
+ cgidl = 0.22
+ pcit = -3.3161007e-17
+ pclm = 0.34708024
+ mobmod = 0
+ njtsswg = 9
+ phin = 0.15
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ pkt1 = -1.1050175e-15
+ pkt2 = -1.739649e-15
+ pbswd = 0.8
+ pbsws = 0.8
+ a0 = 1.2892878
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 51380.779
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = -0.033282087
+ k3 = -1.8419
+ em = 1000000.0
+ ckappad = 0.6
+ ckappas = 0.6
+ ll = -1.18e-13
+ lw = 0
+ u0 = 0.011299764
+ w0 = 0
+ ua = -2.2703742e-9
+ ub = 2.053795462e-18
+ uc = 5.2246809e-11
+ ud = 0
+ pdiblc1 = 0
+ pdiblc2 = 0.010471563
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 6e-9
+ pdiblcb = -0.3
+ rbdb = 50
+ pua1 = -9.0422848e-24
+ prwb = 0
+ pdits = 0
+ laigsd = -6.8373623e-17
+ prwg = 0
+ pub1 = 1.3277736e-32
+ puc1 = 4.9546192e-24
+ cigsd = 0.069865
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ rdsw = 100
+ ijthsfwd = 0.01
+ bigbacc = 0.002588
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ kvth0we = 0.00018
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ tnoia = 0
+ ijthsrev = 0.01
+ lintnoi = -1.5e-8
+ bigbinv = 0.004953
+ peta0 = 0
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ rshg = 15.6
+ wketa = -5.2502872e-8
+ tpbsw = 0.0019
+ cjswd = 8.2e-11
+ cjsws = 8.2e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ ppdiblc2 = -3.8331042e-16
+ toxref = 3e-9
+ tnom = 25
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ scref = 1e-6
+ tvfbsdoff = 0.022
+ pigcd = 2.621
+ aigsd = 0.010772862
+ nfactor = 1
+ ltvoff = 9.6416574e-11
+ wags = -1.195467e-6
+ lvoff = -8.878213999999996e-10
+ pkvth0we = -1.3e-19
+ wcit = 1.6500316e-10
+ lvsat = -0.00023817471000000005
+ lvth0 = -6.196310299999999e-9
+ voff = -0.16014500000000004
+ acde = 0.4
+ delta = 0.007595625
+ laigc = -1.4310771e-11
+ vfbsdoff = 0.02
+ vsat = 114971.1026
+ wint = 0
+ vth0 = 0.42159110699999996
+ rnoia = 0
+ rnoib = 0
+ lku0we = 2.5e-11
+ wkt1 = -9.9137768e-9
+ wkt2 = 1.0152376e-8
+ nigbacc = 10
+ wmax = 9e-7
+ epsrox = 3.9
+ aigc = 0.011560684
+ wmin = 5.4e-7
+ wvfbsdoff = 0
+ pketa = 1.139354e-14
+ lvfbsdoff = 0
+ ngate = 8e+20
+ rdsmod = 0
+ ngcon = 1
+ paramchk = 1
+ wpclm = 8.9560432e-7
+ igbmod = 1
+ wua1 = 5.7543559e-17
+ wub1 = -8.4794537e-26
+ wuc1 = -5.6143964e-17
+ gbmin = 1e-12
+ nigbinv = 10
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ bigc = 0.001442
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ wwlc = 0
+ pbswgd = 0.95
+ pbswgs = 0.95
+ cdsc = 0
+ igcmod = 1
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ ijthdfwd = 0.01
+ xtis = 3
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ fnoimod = 1
+ eigbinv = 1.1
+ ags = 5.1895
+ ijthdrev = 0.01
+ cjd = 0.001357
+ cit = 0.0014357747
+ cjs = 0.001357
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 1.30529375e-8
+ paigsd = 4.6587859e-23
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ tvoff = 0.00014539643
+ lpdiblc2 = -2.045371e-10
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ permod = 1
+ la0 = 6.8373618e-8
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = 0.0010100743
+ kt1 = -0.28113564
+ lk2 = -2.0436616e-10
+ kt2 = -0.099392124
+ llc = -1.18e-13
+ lln = 0.7
+ wtvfbsdoff = 0
+ lu0 = -2.2761917e-10
+ mjd = 0.26
+ lua = 1.7344554e-17
+ mjs = 0.26
+ lub = -2.7790142600000004e-26
+ luc = -5.3126584e-18
+ lud = 0
+ k2we = 5e-5
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = -4.6587862e-14
+ nsd = 1e+20
+ dsub = 0.75
+ pbd = 0.52
+ pat = -1.7932973e-9
+ pbs = 0.52
+ pk2 = -1.7344476e-15
+ cigbacc = 0.32875
+ dtox = 2.7e-10
+ ku0we = -0.0007
+ pu0 = 3.028211e-18
+ beta0 = 13
+ prt = 0
+ pua = 1.2335294e-23
+ pub = -1.88032504e-32
+ puc = -1.1996375e-24
+ pud = 0
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ leta0 = 0
+ ltvfbsdoff = 0
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 6.1325358e-10
+ ub1 = -3.2064524e-19
+ uc1 = 1.2275615e-10
+ tnoimod = 0
+ tpb = 0.0014
+ ppclm = -6.7808634e-14
+ wa0 = -8.7848444e-7
+ voffcv = -0.16942
+ wpemod = 1
+ ute = -1
+ wat = 0.016319757
+ eta0 = 0.42133333
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 1.0517006e-8
+ lkvth0we = -2e-12
+ etab = -0.29033333
+ wlc = 0
+ wln = 1
+ wu0 = -9.6797711e-11
+ xgl = -1.09e-8
+ xgw = 0
+ dlcig = 2.5e-9
+ wua = -7.6059319e-17
+ wub = 9.256491399999999e-26
+ wuc = 4.1739756e-18
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ bgidl = 2320000000.0
+ cigbinv = 0.006
+ )

.model nch_tt_22 nmos (
+ level = 54
+ phin = 0.15
+ cjswd = 8.2e-11
+ cjsws = 8.2e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ pkt1 = -2.447551e-15
+ pkt2 = 8.0276583e-16
+ ptvoff = -9.1490879e-17
+ nfactor = 1
+ paramchk = 1
+ waigsd = 3.0879615e-12
+ diomod = 1
+ rbdb = 50
+ pua1 = -1.6477593e-25
+ prwb = 0
+ prwg = 0
+ pub1 = 1.4533022e-32
+ puc1 = 1.092524e-23
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ pditsd = 0
+ pditsl = 0
+ rbsb = 50
+ pvag = 1.2
+ cjswgd = 2.82e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.82e-10
+ rdsw = 100
+ ijthdfwd = 0.01
+ scref = 1e-6
+ tvfbsdoff = 0.022
+ nigbacc = 10
+ pigcd = 2.621
+ aigsd = 0.010772861
+ mjswgd = 0.85
+ mjswgs = 0.85
+ lvoff = -4.968304999999992e-10
+ tcjswg = 0.001
+ lvsat = 0.001475182984
+ ijthdrev = 0.01
+ lvth0 = 2.877403999999998e-10
+ nigbinv = 10
+ delta = 0.007595625
+ rshg = 15.6
+ laigc = -8.7106488e-12
+ lpdiblc2 = -4.1841324e-15
+ rnoia = 0
+ rnoib = 0
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ pketa = -2.7052976e-14
+ ngate = 8e+20
+ ngcon = 1
+ wpclm = 4.0103412e-7
+ fnoimod = 1
+ fprout = 300
+ eigbinv = 1.1
+ gbmin = 1e-12
+ tnom = 25
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ xrcrg1 = 12
+ xrcrg2 = 1
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ lkvth0we = -2e-12
+ wtvoff = 7.682212e-10
+ ags = 5.1895
+ cjd = 0.001357
+ cit = 0.00076911293
+ cjs = 0.001357
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ acnqsmod = 0
+ dlc = 3.26497e-9
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ wags = -1.195467e-6
+ capmod = 2
+ wcit = -2.7211371e-10
+ cigbacc = 0.32875
+ rbodymod = 0
+ wku0we = 2e-11
+ la0 = -1.9182963e-7
+ voff = -0.164304478
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.0016942500800000001
+ acde = 0.4
+ kt1 = -0.33033037
+ lk2 = -1.3785596e-9
+ kt2 = -0.066210327
+ mobmod = 0
+ llc = 0
+ lln = 1
+ lu0 = -6.7155919e-11
+ tnoimod = 0
+ mjd = 0.26
+ tvoff = 0.00053139469
+ lua = 2.7860169e-17
+ mjs = 0.26
+ lub = -2.7395085e-26
+ luc = 1.41139916e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ vsat = 96743.889
+ njs = 1.02
+ pa0 = 2.0809981e-13
+ wint = 0
+ vth0 = 0.352611848
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 2.0789444199999997e-9
+ pbs = 0.52
+ pk2 = 9.5324632e-16
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ wkt1 = 4.3684939e-9
+ wkt2 = -1.689459e-8
+ pu0 = -2.5471417e-18
+ wmax = 9e-7
+ prt = 0
+ pua = -6.3654423e-24
+ pub = 7.034010899999999e-33
+ puc = -7.127418999999999e-24
+ pud = 0
+ cigbinv = 0.006
+ aigc = 0.011501109
+ wmin = 5.4e-7
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 8.1588744e-10
+ ub1 = -6.9089562e-19
+ uc1 = 1.6549472299999998e-10
+ tpb = 0.0014
+ wa0 = -3.5879278e-6
+ ute = -1
+ wat = -0.024874303599999998
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -1.8075483e-8
+ ku0we = -0.0007
+ wlc = 0
+ wln = 1
+ wu0 = -3.7485448e-11
+ xgl = -1.09e-8
+ xgw = 0
+ beta0 = 13
+ wua = 1.2288469e-16
+ wub = -1.8229956900000002e-25
+ wua1 = -3.6898024e-17
+ wuc = 6.7235478e-17
+ wud = 0
+ wub1 = -9.8148649e-26
+ wuc1 = -1.19661208e-16
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ leta0 = -1.0826782e-8
+ wpdiblc2 = -5.8202891e-10
+ letab = -2.2164189e-8
+ version = 4.5
+ bigc = 0.001442
+ laigsd = 3.8113519e-17
+ tempmod = 0
+ wwlc = 0
+ ppclm = -2.1319035e-14
+ dlcig = 2.5e-9
+ cdsc = 0
+ bgidl = 2320000000.0
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ aigbacc = 0.02
+ xtis = 3
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ dmcgt = 0
+ tcjsw = 0.000357
+ wkvth0we = 2e-12
+ aigbinv = 0.0163
+ a0 = 4.0574074
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 80150.18699999999
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = -0.020790667
+ k3 = -1.8419
+ em = 1000000.0
+ ll = 0
+ lw = 0
+ trnqsmod = 0
+ u0 = 0.009592708
+ w0 = 0
+ ua = -2.3822425e-9
+ ub = 2.049592666e-18
+ uc = -1.5441968e-10
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 6e-9
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ bigsd = 0.00125
+ wvoff = 3.044252900000001e-8
+ k2we = 5e-5
+ dsub = 0.75
+ dtox = 2.7e-10
+ wvsat = -0.017460159999999995
+ toxref = 3e-9
+ wvth0 = -3.533284300000001e-8
+ rgatemod = 0
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ tnjtsswg = 1
+ poxedge = 1
+ waigc = 1.9067031e-10
+ eta0 = 0.53651186
+ etab = -0.054544089
+ binunit = 2
+ lketa = 6.7720908e-8
+ xpart = 1
+ ltvoff = 6.0132739e-11
+ egidl = 0.29734
+ pvfbsdoff = 0
+ lku0we = 2.5e-11
+ epsrox = 3.9
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ rdsmod = 0
+ igbmod = 1
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ pvoff = -1.5223199999999999e-15
+ pbswgd = 0.95
+ pbswgs = 0.95
+ cdscb = 0
+ cdscd = 0
+ pvsat = 5.593105999999996e-10
+ wk2we = 5e-12
+ igcmod = 1
+ pvth0 = 1.8721500000000003e-15
+ drout = 0.56
+ paigc = -1.0723924e-17
+ ijthsfwd = 0.01
+ njtsswg = 9
+ voffl = 0
+ keta = -1.0362685
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ weta0 = -2.7932191e-7
+ wetab = 6.5877739e-8
+ wtvfbsdoff = 0
+ lpclm = -1.3225653e-8
+ ckappad = 0.6
+ ckappas = 0.6
+ jswd = 1.28e-13
+ pdiblc1 = 0
+ jsws = 1.28e-13
+ pdiblc2 = 0.0082956805
+ lcit = 1.2418741e-10
+ paigsd = -2.0809977e-23
+ pdiblcb = -0.3
+ ijthsrev = 0.01
+ kt1l = 0
+ cgidl = 0.22
+ ltvfbsdoff = 0
+ permod = 1
+ lint = 0
+ lkt1 = 5.3401869e-9
+ lkt2 = -2.1703039e-9
+ lmax = 9e-8
+ lmin = 5.4e-8
+ pbswd = 0.8
+ pbsws = 0.8
+ bigbacc = 0.002588
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ ppdiblc2 = 5.6582339e-21
+ minv = -0.3
+ kvth0we = 0.00018
+ lua1 = -4.7634626e-18
+ lub1 = -2.8456569e-26
+ luc1 = -9.937027189999999e-18
+ voffcv = -0.16942
+ wpemod = 1
+ pdits = 0
+ ndep = 1e+18
+ lintnoi = -1.5e-8
+ cigsd = 0.069865
+ ptvfbsdoff = 0
+ lwlc = 0
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ moin = 5.1
+ vtsswgs = 4.2
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ nigc = 3.083
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ pkvth0we = -1.3e-19
+ tnoia = 0
+ tpbswg = 0.0009
+ peta0 = 1.5923028e-14
+ ntox = 1
+ pcit = 7.9279785e-18
+ petab = -3.6091995e-15
+ pclm = 1.1225851
+ vfbsdoff = 0.02
+ wketa = 3.5650261e-7
+ tpbsw = 0.0019
+ )

.model nch_tt_23 nmos (
+ level = 54
+ pditsl = 0
+ cjswgd = 2.82e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.82e-10
+ cdsc = 0
+ lketa = -2.0578185e-8
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ ijthsfwd = 0.01
+ xtid = 3
+ xtis = 3
+ xpart = 1
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ mjswgd = 0.85
+ mjswgs = 0.85
+ egidl = 0.29734
+ tcjswg = 0.001
+ pvfbsdoff = 0
+ ijthsrev = 0.01
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ njtsswg = 9
+ k2we = 5e-5
+ dsub = 0.75
+ dtox = 2.7e-10
+ fprout = 300
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ xrcrg1 = 12
+ xrcrg2 = 1
+ pvoff = -3.925098540000001e-15
+ ckappad = 0.6
+ ckappas = 0.6
+ cdscb = 0
+ pdiblc1 = 0
+ pdiblc2 = 0.0082956083
+ cdscd = 0
+ pdiblcb = -0.3
+ pvsat = 4.031319111000001e-9
+ eta0 = 0.49180426
+ etab = -1.1686036
+ wk2we = 5e-12
+ pvth0 = 4.7434049e-15
+ drout = 0.56
+ wtvoff = -4.625476e-9
+ paigc = -1.7630641e-18
+ voffl = 0
+ weta0 = 1.6706711e-7
+ capmod = 2
+ bigbacc = 0.002588
+ wetab = -6.7375536e-8
+ pkvth0we = -1.3e-19
+ lpclm = -4.9784452e-8
+ wku0we = 2e-11
+ mobmod = 0
+ kvth0we = 0.00018
+ cgidl = 0.22
+ vfbsdoff = 0.02
+ lintnoi = -1.5e-8
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ pbswd = 0.8
+ pbsws = 0.8
+ paramchk = 1
+ laigsd = -3.1577826e-17
+ pdits = 0
+ cigsd = 0.069865
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ ijthdfwd = 0.01
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ keta = 0.48612964
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ nfactor = 1
+ tnoia = 0
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ ijthdrev = 0.01
+ lcit = 3.8601345e-10
+ peta0 = -9.9675358e-15
+ kt1l = 0
+ petab = 4.1194905e-15
+ wketa = -1.8474011e-7
+ tpbsw = 0.0019
+ lint = 0
+ cjswd = 8.2e-11
+ cjsws = 8.2e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ lkt1 = -1.4874128e-8
+ lkt2 = -1.4213753e-9
+ lmax = 5.4e-8
+ lmin = 4.5e-8
+ nigbacc = 10
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ toxref = 3e-9
+ minv = -0.3
+ lua1 = 7.7308837e-17
+ lub1 = -1.58914262e-25
+ luc1 = -7.236573999999998e-18
+ ndep = 1e+18
+ lkvth0we = -2e-12
+ nigbinv = 10
+ lwlc = 0
+ moin = 5.1
+ a0 = 11.080765
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 31524.241299999994
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ tvfbsdoff = 0.022
+ k2 = 0.013147898
+ k3 = -1.8419
+ em = 1000000.0
+ ll = 0
+ lw = 0
+ u0 = -0.00068107274
+ scref = 1e-6
+ nigc = 3.083
+ w0 = 0
+ ua = -5.2066121e-9
+ ub = 5.20056154e-18
+ uc = 2.7090556e-10
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 6e-9
+ pigcd = 2.621
+ aigsd = 0.010772862
+ ltvoff = -1.4697355e-10
+ acnqsmod = 0
+ lvoff = 1.6118058999999991e-9
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ fnoimod = 1
+ lvsat = -0.005682873369999999
+ rbodymod = 0
+ lvth0 = -3.5936672999999988e-9
+ eigbinv = 1.1
+ ntox = 1
+ delta = 0.007595625
+ pcit = 2.2096077e-17
+ lku0we = 2.5e-11
+ pclm = 1.7529092
+ laigc = -1.8175152e-11
+ epsrox = 3.9
+ rnoia = 0
+ rnoib = 0
+ wvfbsdoff = 0
+ phin = 0.15
+ lvfbsdoff = 0
+ rdsmod = 0
+ pketa = 4.339103e-15
+ igbmod = 1
+ ngate = 8e+20
+ pkt1 = 1.1940455e-14
+ pkt2 = 3.1759909e-15
+ ngcon = 1
+ wpclm = -7.2697212e-7
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ wpdiblc2 = -5.8193135e-10
+ pbswgd = 0.95
+ gbmin = 1e-12
+ pbswgs = 0.95
+ cigbacc = 0.32875
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ ags = 5.1895
+ rbdb = 50
+ pua1 = -6.2039198e-23
+ prwb = 0
+ prwg = 0
+ pub1 = 1.08440889e-31
+ puc1 = 1.0847755599999997e-23
+ igcmod = 1
+ wtvfbsdoff = 0
+ cjd = 0.001357
+ cit = -0.0037451293
+ cjs = 0.001357
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ dlc = 3.26497e-9
+ k3b = 1.9326
+ tnoimod = 0
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ rdsw = 100
+ ltvfbsdoff = 0
+ cigbinv = 0.006
+ la0 = -5.9918439e-7
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = 0.0011260548200000002
+ kt1 = 0.018192305
+ lk2 = -3.3469964e-9
+ kt2 = -0.079122889
+ llc = 0
+ lln = 1
+ lu0 = 5.2872336e-10
+ mjd = 0.26
+ lua = 1.9167361e-16
+ mjs = 0.26
+ lub = -2.101512744e-25
+ luc = -1.0554871600000002e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 1.4611928e-13
+ wkvth0we = 2e-12
+ nsd = 1e+20
+ pbd = 0.52
+ pat = -1.44553358e-9
+ pbs = 0.52
+ pk2 = 2.1253177e-15
+ paigsd = 1.0451534e-29
+ pu0 = -5.7605924e-17
+ prt = 0
+ pua = -7.1470289e-23
+ pub = 9.665873609999999e-32
+ puc = 4.556057900000002e-24
+ pud = 0
+ version = 4.5
+ rsh = 17.5
+ trnqsmod = 0
+ tcj = 0.00076
+ ua1 = -5.9915221e-10
+ ub1 = 1.5583749700000001e-18
+ uc1 = 1.1893518999999988e-10
+ rshg = 15.6
+ tempmod = 0
+ tvoff = 0.0041021928
+ tpb = 0.0014
+ wa0 = -2.5192978e-6
+ permod = 1
+ ute = -1
+ wat = 0.035892558
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -3.8283609e-8
+ xjbvd = 1
+ xjbvs = 1
+ wlc = 0
+ wln = 1
+ lk2we = -1.5e-12
+ wu0 = 9.118039e-10
+ xgl = -1.09e-8
+ xgw = 0
+ wua = 1.2453821e-15
+ wub = -1.72755342e-24
+ wuc = -1.3420376999999993e-16
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ ptvfbsdoff = 0
+ aigbacc = 0.02
+ ku0we = -0.0007
+ beta0 = 13
+ rgatemod = 0
+ leta0 = -8.2337409e-9
+ letab = 4.245126e-8
+ voffcv = -0.16942
+ wpemod = 1
+ tnom = 25
+ tnjtsswg = 1
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ aigbinv = 0.0163
+ ppclm = 4.4105328e-14
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ wags = -1.195467e-6
+ dmcgt = 0
+ tcjsw = 0.000357
+ wcit = -5.1639126e-10
+ tpbswg = 0.0009
+ voff = -0.20066027000000003
+ acde = 0.4
+ poxedge = 1
+ vsat = 220158.66399999996
+ wint = 0
+ vth0 = 0.41953267
+ bigsd = 0.00125
+ binunit = 2
+ wkt1 = -2.4370058e-7
+ wkt2 = -5.7812263e-8
+ wmax = 9e-7
+ aigc = 0.01166429
+ wmin = 5.4e-7
+ ptvoff = 2.2134356e-16
+ wvoff = 7.186973409999998e-8
+ waigsd = 3.0876027e-12
+ wvsat = -0.07732237247
+ wua1 = 1.0299024e-15
+ wub1 = -1.71724981e-24
+ wuc1 = -1.1832528899999998e-16
+ wvth0 = -8.483723199999998e-8
+ diomod = 1
+ bigc = 0.001442
+ waigc = 3.6172725e-11
+ wwlc = 0
+ pditsd = 0
+ )

.model nch_tt_24 nmos (
+ level = 54
+ lvsat = -0.0030618311999999993
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lvth0 = 3.859772699999999e-9
+ lcit = 1.5105388e-10
+ trnqsmod = 0
+ kt1l = 0
+ cigbacc = 0.32875
+ delta = 0.007595625
+ laigc = -7.4258513e-12
+ rnoia = 0
+ rnoib = 0
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ tnoimod = 0
+ lint = 0
+ lkt1 = 1.0114149e-9
+ lkt2 = 6.4873536e-9
+ lmax = 4.5e-8
+ pketa = 3.05233408e-14
+ ags = 5.1895
+ ngate = 8e+20
+ lmin = 3.6e-8
+ cigbinv = 0.006
+ ngcon = 1
+ lpe0 = 9.2e-8
+ cjd = 0.001357
+ cit = 0.001049964
+ fprout = 300
+ cjs = 0.001357
+ clc = 1e-7
+ wpclm = 9.524622100000001e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ lpeb = 2.5e-7
+ dlc = 3.26497e-9
+ k3b = 1.9326
+ xrcrg1 = 12
+ xrcrg2 = 1
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ rgatemod = 0
+ gbmin = 1e-12
+ minv = -0.3
+ tnjtsswg = 1
+ lua1 = -6.7547343e-17
+ lub1 = 1.29809254e-25
+ luc1 = 1.834266e-17
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ ndep = 1e+18
+ la0 = -5.581062559999999e-7
+ version = 4.5
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.00167504779
+ wtvoff = -5.6534448e-10
+ lwlc = 0
+ kt1 = -0.30600245
+ lk2 = -3.4047834e-9
+ kt2 = -0.24052552
+ llc = 0
+ moin = 5.1
+ lln = 1
+ lu0 = 8.1748395e-10
+ tempmod = 0
+ mjd = 0.26
+ lua = 1.9963428e-16
+ mjs = 0.26
+ lub = -1.86515944e-25
+ luc = -1.3855022100000003e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 1.41312605e-13
+ nigc = 3.083
+ nsd = 1e+20
+ pbd = 0.52
+ pat = -1.7010081000000005e-10
+ pbs = 0.52
+ pk2 = 1.540171e-16
+ pu0 = -4.6401651e-16
+ prt = 0
+ pua = -1.24177601e-22
+ pub = 1.2166737845000001e-31
+ puc = -3.231882900000001e-24
+ pud = 0
+ aigbacc = 0.02
+ capmod = 2
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 2.3570964e-9
+ ub1 = -4.3339417e-18
+ uc1 = -4.0308999999999995e-10
+ tpb = 0.0014
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ wku0we = 2e-11
+ wa0 = -2.4212027299999997e-6
+ ute = -1
+ wat = 0.009863318999999999
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 1.947015e-9
+ wlc = 0
+ wln = 1
+ wu0 = 9.2058975e-9
+ xgl = -1.09e-8
+ mobmod = 0
+ xgw = 0
+ wua = 2.32104147e-15
+ wub = -2.2379339299999998e-24
+ wuc = 2.4733810000000014e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ ntox = 1
+ pcit = 4.8523743e-17
+ pclm = 0.021884800000000038
+ tvoff = 0.0045807103
+ aigbinv = 0.0163
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ phin = 0.15
+ pkt1 = -5.2985624e-15
+ pkt2 = -2.9889728e-15
+ ku0we = -0.0007
+ beta0 = 13
+ laigsd = 2.1777751e-17
+ leta0 = 6.023777099999999e-9
+ letab = 3.2196399e-8
+ ppclm = -3.8186956000000005e-14
+ rbdb = 50
+ pua1 = 5.0551945e-23
+ prwb = 0
+ prwg = 0
+ pub1 = -9.568911599999999e-32
+ puc1 = -1.81613879e-23
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ poxedge = 1
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ rdsw = 100
+ ijthsfwd = 0.01
+ binunit = 2
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ dmcgt = 0
+ tcjsw = 0.000357
+ ijthsrev = 0.01
+ rshg = 15.6
+ bigsd = 0.00125
+ wvoff = -2.5396920999999984e-8
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ toxref = 3e-9
+ wvsat = -0.033609850999999996
+ wvth0 = 4.0967673000000005e-8
+ tnom = 25
+ waigc = -1.3685053e-10
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ lketa = -4.89346675e-8
+ xpart = 1
+ ltvoff = -1.7042091e-10
+ egidl = 0.29734
+ njtsswg = 9
+ wags = -1.195467e-6
+ pkvth0we = -1.3e-19
+ pvfbsdoff = 0
+ wcit = -1.0557314e-9
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ voff = -0.003529144999999956
+ lku0we = 2.5e-11
+ acde = 0.4
+ ckappad = 0.6
+ epsrox = 3.9
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.0082956083
+ vfbsdoff = 0.02
+ pdiblcb = -0.3
+ vsat = 166667.996
+ wint = 0
+ vth0 = 0.267421665
+ wkt1 = 1.0811611e-7
+ wkt2 = 6.8003321e-8
+ rdsmod = 0
+ wtvfbsdoff = 0
+ wmax = 9e-7
+ aigc = 0.011444916
+ wmin = 5.4e-7
+ igbmod = 1
+ a0 = 10.24243689
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 88689.602
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.014327223
+ k3 = -1.8419
+ em = 1000000.0
+ ll = 0
+ lw = 0
+ u0 = -0.0065741458
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ paramchk = 1
+ w0 = 0
+ ua = -5.369074800000001e-9
+ ub = 4.718207719999999e-18
+ uc = 3.3825556e-10
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 6e-9
+ ltvfbsdoff = 0
+ pbswgd = 0.95
+ pbswgs = 0.95
+ wua1 = -1.2678761e-15
+ wub1 = 2.44866871e-24
+ wuc1 = 4.7369808e-16
+ bigbacc = 0.002588
+ pvoff = 8.409683299999991e-16
+ bigc = 0.001442
+ igcmod = 1
+ wwlc = 0
+ cdscb = 0
+ cdscd = 0
+ kvth0we = 0.00018
+ pvsat = 1.88940533e-9
+ wk2we = 5e-12
+ pvth0 = -1.4210356999999999e-15
+ drout = 0.56
+ cdsc = 0
+ lintnoi = -1.5e-8
+ paigc = 6.7150752e-18
+ cgbo = 0
+ ijthdfwd = 0.01
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ voffl = 0
+ cigc = 0.000625
+ ptvfbsdoff = 0
+ weta0 = -1.6294544599999998e-7
+ wetab = 1.0177792e-7
+ paigsd = 4.9710031e-30
+ lpclm = 3.5035747999999996e-8
+ ijthdrev = 0.01
+ cgidl = 0.22
+ permod = 1
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ pbswd = 0.8
+ pbsws = 0.8
+ k2we = 5e-5
+ dsub = 0.75
+ dtox = 2.7e-10
+ voffcv = -0.16942
+ wpemod = 1
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ nfactor = 1
+ pdits = 0
+ cigsd = 0.069865
+ eta0 = 0.20083450200000003
+ lkvth0we = -2e-12
+ etab = -0.95932067
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ acnqsmod = 0
+ nigbacc = 10
+ tpbswg = 0.0009
+ tnoia = 0
+ rbodymod = 0
+ peta0 = 6.20307972e-15
+ petab = -4.1690291e-15
+ wketa = -7.1911233e-7
+ tpbsw = 0.0019
+ nigbinv = 10
+ cjswd = 8.2e-11
+ cjsws = 8.2e-11
+ ptvoff = 2.2397114e-17
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ waigsd = 3.0876027e-12
+ diomod = 1
+ wpdiblc2 = -5.8193135e-10
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 2.82e-10
+ pku0we = -1.5e-18
+ fnoimod = 1
+ cjswgs = 2.82e-10
+ eigbinv = 1.1
+ tvfbsdoff = 0.022
+ scref = 1e-6
+ pigcd = 2.621
+ mjswgd = 0.85
+ aigsd = 0.010772861
+ mjswgs = 0.85
+ keta = 1.06483334
+ tcjswg = 0.001
+ lvoff = -8.047620000000002e-9
+ wkvth0we = 2e-12
+ )

.model nch_tt_25 nmos (
+ level = 54
+ fprout = 300
+ xrcrg1 = 12
+ xrcrg2 = 1
+ pvoff = 0
+ tnom = 25
+ cdscb = 0
+ cdscd = 0
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ wtvoff = 0
+ pvsat = 0
+ lkvth0we = -2e-12
+ wk2we = 5e-12
+ pvth0 = 0
+ drout = 0.56
+ voffl = 0
+ capmod = 2
+ acnqsmod = 0
+ wku0we = 2e-11
+ weta0 = -1.1162667e-8
+ wags = -6.546904e-8
+ wetab = 2.2325333e-8
+ mobmod = 0
+ wcit = 2.963688e-10
+ rbodymod = 0
+ nfactor = 1
+ voff = -0.13478422
+ acde = 0.4
+ cgidl = 0.22
+ vsat = 102889.02
+ wint = 0
+ vth0 = 0.36420512
+ wkt1 = -9.7059387e-11
+ wkt2 = -5.3296152e-9
+ wmax = 5.4e-7
+ aigc = 0.011779434
+ wmin = 2.7e-7
+ pbswd = 0.8
+ pbsws = 0.8
+ wua1 = -1.874362e-16
+ nigbacc = 10
+ wub1 = 1.1464267e-25
+ wuc1 = -2.7527136e-17
+ wpdiblc2 = 4.9914968e-9
+ bigc = 0.001442
+ pdits = 0
+ wwlc = 0
+ cigsd = 0.069865
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ nigbinv = 10
+ xtis = 3
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ wkvth0we = 2e-12
+ tnoia = 0
+ trnqsmod = 0
+ peta0 = 0
+ fnoimod = 1
+ wketa = 1.6322115e-8
+ eigbinv = 1.1
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ tpbsw = 0.0019
+ dmdg = 0
+ cjswd = 8.2e-11
+ cjsws = 8.2e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ toxref = 3e-9
+ k2we = 5e-5
+ dsub = 0.75
+ dtox = 2.7e-10
+ rgatemod = 0
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ tnjtsswg = 1
+ tvfbsdoff = 0.022
+ eta0 = 0.24044444
+ etab = -0.28088889
+ cigbacc = 0.32875
+ ltvoff = 0
+ scref = 1e-6
+ pigcd = 2.621
+ tnoimod = 0
+ aigsd = 0.010772818
+ wtvfbsdoff = 0
+ lvoff = 0
+ cigbinv = 0.006
+ lvsat = 0
+ lku0we = 2.5e-11
+ lvth0 = 0
+ ltvfbsdoff = 0
+ epsrox = 3.9
+ delta = 0.007595625
+ ags = 0.98760667
+ wvfbsdoff = 0
+ cjd = 0.001357
+ cit = 0.000342575
+ version = 4.5
+ cjs = 0.001357
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ lvfbsdoff = 0
+ rnoia = 0
+ rnoib = 0
+ rdsmod = 0
+ dlc = 9.8024918e-9
+ k3b = 1.9326
+ tempmod = 0
+ igbmod = 1
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ ngate = 8e+20
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ ngcon = 1
+ la0 = 0
+ wpclm = 9.3989653e-8
+ pbswgd = 0.95
+ jsd = 6.11e-7
+ pbswgs = 0.95
+ jss = 6.11e-7
+ lat = 0
+ aigbacc = 0.02
+ kt1 = -0.22055704
+ kt2 = -0.0354368
+ llc = 0
+ lln = 1
+ lu0 = 0
+ mjd = 0.26
+ mjs = 0.26
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ gbmin = 1e-12
+ njs = 1.02
+ pa0 = 0
+ igcmod = 1
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 0
+ jswgd = 1.28e-13
+ ptvfbsdoff = 0
+ pbs = 0.52
+ jswgs = 1.28e-13
+ pu0 = 0
+ prt = 0
+ pud = 0
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 1.6212811e-9
+ ub1 = -8.7849211e-19
+ uc1 = 6.9356e-11
+ tpb = 0.0014
+ aigbinv = 0.0163
+ wa0 = -1.17208e-8
+ ijthsfwd = 0.01
+ ute = -1
+ wat = 0.071441067
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 1.8596306e-9
+ wlc = 0
+ wln = 1
+ wu0 = -1.2837067e-9
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -1.3097991e-16
+ wub = 9.54408e-26
+ wuc = -2.4557867e-18
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ keta = -0.084351302
+ a0 = 3.5424667
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = -58844.444
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.020167646
+ k3 = -1.8419
+ em = 1000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.017671111
+ jswd = 1.28e-13
+ w0 = 0
+ jsws = 1.28e-13
+ ijthsrev = 0.01
+ ua = -1.6762565e-9
+ ub = 2.0222e-18
+ uc = 6.1497778e-11
+ ud = 0
+ lcit = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 6e-9
+ permod = 1
+ kt1l = 0
+ tvoff = 0.0017628809
+ xjbvd = 1
+ xjbvs = 1
+ poxedge = 1
+ lk2we = -1.5e-12
+ lint = 6.5375218e-9
+ lkt1 = 0
+ lmax = 2.001e-5
+ binunit = 2
+ lmin = 8.9991e-6
+ lpe0 = 9.2e-8
+ voffcv = -0.16942
+ wpemod = 1
+ lpeb = 2.5e-7
+ ku0we = -0.0007
+ beta0 = 13
+ leta0 = 0
+ minv = -0.3
+ lub1 = 0
+ ndep = 1e+18
+ lwlc = 0
+ dlcig = 2.5e-9
+ moin = 5.1
+ bgidl = 2320000000.0
+ nigc = 3.083
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ noff = 2.7195
+ dmcgt = 0
+ noia = 3.11e+42
+ noib = 1.22e+22
+ pkvth0we = -1.3e-19
+ noic = 45200000.0
+ tpbswg = 0.0009
+ tcjsw = 0.000357
+ ntox = 1
+ pcit = 0
+ pclm = 1.5094578
+ vfbsdoff = 0.02
+ bigsd = 0.00125
+ ptvoff = 0
+ phin = 0.15
+ waigsd = 3.1112026e-12
+ wvoff = 1.3685577e-8
+ pkt1 = 0
+ paramchk = 1
+ diomod = 1
+ wvsat = -0.0028059037
+ wvth0 = -1.7768414e-8
+ njtsswg = 9
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 2.82e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.82e-10
+ waigc = 2.8724444e-11
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ rbdb = 50
+ prwb = 0
+ prwg = 0
+ pub1 = 0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.0047029422
+ rdsw = 100
+ pdiblcb = -0.3
+ ijthdfwd = 0.01
+ mjswgd = 0.85
+ xpart = 1
+ mjswgs = 0.85
+ tcjswg = 0.001
+ egidl = 0.29734
+ pvfbsdoff = 0
+ bigbacc = 0.002588
+ ijthdrev = 0.01
+ rshg = 15.6
+ kvth0we = 0.00018
+ lintnoi = -1.5e-8
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ )

.model nch_tt_26 nmos (
+ level = 54
+ poxedge = 1
+ capmod = 2
+ wku0we = 2e-11
+ binunit = 2
+ mobmod = 0
+ pkvth0we = -1.3e-19
+ tvoff = 0.0019388906
+ vfbsdoff = 0.02
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ laigsd = -2.019482e-16
+ paramchk = 1
+ ku0we = -0.0007
+ beta0 = 13
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ leta0 = 0
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ ijthdfwd = 0.01
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ keta = -0.091670067
+ dmcgt = 0
+ tcjsw = 0.000357
+ lags = -1.7808411e-7
+ njtsswg = 9
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ ijthdrev = 0.01
+ lcit = 6.6778289e-10
+ kt1l = 0
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ lpdiblc2 = 2.6261368e-8
+ bigsd = 0.00125
+ ckappad = 0.6
+ ckappas = 0.6
+ lint = 6.5375218e-9
+ pdiblc1 = 0
+ pdiblc2 = 0.0017817666
+ toxref = 3e-9
+ pdiblcb = -0.3
+ lkt1 = 9.0572759e-9
+ lkt2 = -2.1662043e-8
+ lmax = 8.9991e-6
+ wvoff = 1.395365e-8
+ lmin = 8.9908e-7
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ wvsat = -0.0028059037
+ wvth0 = -1.8116317e-8
+ minv = -0.3
+ wtvfbsdoff = 0
+ lua1 = -8.9279603e-16
+ lub1 = 6.8544226e-25
+ luc1 = -5.9256432e-18
+ waigc = 2.989874e-11
+ bigbacc = 0.002588
+ ndep = 1e+18
+ lkvth0we = -2e-12
+ lwlc = 0
+ moin = 5.1
+ ltvoff = -1.582327e-9
+ ltvfbsdoff = 0
+ lketa = 6.5795695e-8
+ kvth0we = 0.00018
+ nigc = 3.083
+ xpart = 1
+ lintnoi = -1.5e-8
+ acnqsmod = 0
+ pvfbsdoff = 0
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ egidl = 0.29734
+ vtsswgs = 4.2
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ lku0we = 2.5e-11
+ rbodymod = 0
+ epsrox = 3.9
+ pags = 1.7531187e-13
+ ntox = 1
+ pcit = -1.0698337e-16
+ pclm = 1.5094578
+ rdsmod = 0
+ ptvfbsdoff = 0
+ igbmod = 1
+ phin = 0.15
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ pbswgd = 0.95
+ pkt1 = -2.7377875e-14
+ pkt2 = -4.4253241e-16
+ pbswgs = 0.95
+ igcmod = 1
+ wpdiblc2 = 5.7318301e-9
+ pvoff = -2.4099793e-15
+ cdscb = 0
+ cdscd = 0
+ rbdb = 50
+ pua1 = 1.9942546e-22
+ prwb = 0
+ prwg = 0
+ pub1 = -1.9939615e-31
+ puc1 = 1.7835157e-23
+ nfactor = 1
+ pvsat = 0
+ rbpb = 50
+ rbpd = 50
+ wk2we = 5e-12
+ rbps = 50
+ pvth0 = 3.1276502e-15
+ rbsb = 50
+ pvag = 1.2
+ drout = 0.56
+ rdsw = 100
+ paigc = -1.0556924e-17
+ voffl = 0
+ paigsd = 1.1026372e-22
+ weta0 = -1.1162667e-8
+ wetab = 2.2325333e-8
+ wkvth0we = 2e-12
+ nigbacc = 10
+ permod = 1
+ trnqsmod = 0
+ cgidl = 0.22
+ rshg = 15.6
+ nigbinv = 10
+ pbswd = 0.8
+ pbsws = 0.8
+ voffcv = -0.16942
+ wpemod = 1
+ rgatemod = 0
+ tnjtsswg = 1
+ tnom = 25
+ pdits = 0
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ a0 = 3.8452644
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ cigsd = 0.069865
+ b1 = 0
+ at = -81312.781
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.021723392
+ k3 = -1.8419
+ em = 1000000.0
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ ll = 0
+ lw = 0
+ u0 = 0.01792456
+ w0 = 0
+ fnoimod = 1
+ ua = -1.6436128e-9
+ ub = 2.0158412e-18
+ uc = 5.8736458e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 6e-9
+ eigbinv = 1.1
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ tpbswg = 0.0009
+ wags = -8.4969804e-8
+ wcit = 3.0826906e-10
+ tnoia = 0
+ voff = -0.13348839
+ peta0 = 0
+ acde = 0.4
+ wketa = 1.8850903e-8
+ vsat = 102889.02
+ ptvoff = 2.7553621e-16
+ wint = 0
+ tpbsw = 0.0019
+ vth0 = 0.35849778
+ cigbacc = 0.32875
+ waigsd = 3.1111904e-12
+ wkt1 = 2.9483105e-9
+ wkt2 = -5.2803902e-9
+ cjswd = 8.2e-11
+ cjsws = 8.2e-11
+ wmax = 5.4e-7
+ mjswd = 0.11
+ aigc = 0.011795195
+ mjsws = 0.11
+ wmin = 2.7e-7
+ agidl = 9.41e-8
+ diomod = 1
+ tnoimod = 0
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 2.82e-10
+ pku0we = -1.5e-18
+ wua1 = -2.0961923e-16
+ wub1 = 1.3682244e-25
+ cjswgs = 2.82e-10
+ wuc1 = -2.9511024e-17
+ cigbinv = 0.006
+ bigc = 0.001442
+ wwlc = 0
+ tvfbsdoff = 0.022
+ cdsc = 0
+ mjswgd = 0.85
+ mjswgs = 0.85
+ scref = 1e-6
+ version = 4.5
+ ijthsfwd = 0.01
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ pigcd = 2.621
+ cgsl = 3.31989e-12
+ tcjswg = 0.001
+ cgso = 4.90562e-11
+ tempmod = 0
+ aigsd = 0.010772818
+ cigc = 0.000625
+ ags = 1.0074158
+ lvoff = -1.1649525e-8
+ cjd = 0.001357
+ cit = 0.00026829437
+ cjs = 0.001357
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ aigbacc = 0.02
+ dlc = 9.8024918e-9
+ lvsat = 0
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ lvth0 = 5.1308999e-8
+ ijthsrev = 0.01
+ delta = 0.007595625
+ laigc = -1.416882e-10
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ la0 = -2.722152e-6
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ rnoia = 0
+ rnoib = 0
+ dmdg = 0
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = 0.20199035
+ kt1 = -0.22156452
+ lk2 = -1.3986155e-8
+ kt2 = -0.033027229
+ llc = 0
+ lln = 1
+ lu0 = -2.2785026e-9
+ mjd = 0.26
+ aigbinv = 0.0163
+ lua = -2.9346741e-16
+ mjs = 0.26
+ lub = 5.7165214e-26
+ luc = 2.4824263e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 3.4236885e-13
+ fprout = 300
+ nsd = 1e+20
+ pbd = 0.52
+ pat = -6.3688324e-8
+ pbs = 0.52
+ pketa = -2.2733801e-14
+ pk2 = -1.3939214e-15
+ ngate = 8e+20
+ pu0 = 1.6539558e-16
+ xrcrg1 = 12
+ xrcrg2 = 1
+ k2we = 5e-5
+ prt = 0
+ pua = 4.226297e-23
+ pub = -4.4156209e-32
+ puc = -1.0695581e-23
+ pud = 0
+ ngcon = 1
+ wpclm = 9.3989653e-8
+ dsub = 0.75
+ rsh = 17.5
+ tcj = 0.00076
+ dtox = 2.7e-10
+ ua1 = 1.720591e-9
+ ub1 = -9.5473708e-19
+ uc1 = 7.0015137e-11
+ ppdiblc2 = -6.6555967e-15
+ tpb = 0.0014
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ wa0 = -4.9804098e-8
+ gbmin = 1e-12
+ ute = -1
+ wat = 0.078525419
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 2.0146831e-9
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ wtvoff = -3.0649189e-11
+ wlc = 0
+ wln = 1
+ wu0 = -1.3021044e-9
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -1.3568102e-16
+ wub = 1.003525e-25
+ wuc = -1.2660669e-18
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ eta0 = 0.24044444
+ etab = -0.28088889
+ )

.model nch_tt_27 nmos (
+ level = 54
+ ntox = 1
+ pcit = -1.1605802e-16
+ pclm = 1.5094578
+ fnoimod = 1
+ phin = 0.15
+ eigbinv = 1.1
+ pbswd = 0.8
+ pbsws = 0.8
+ pkt1 = 4.8128443e-15
+ pkt2 = 2.2738921e-15
+ pdits = 0
+ rbdb = 50
+ pua1 = -2.6369043e-23
+ prwb = 0
+ prwg = 0
+ pub1 = 4.8759292e-32
+ cigsd = 0.069865
+ puc1 = 6.8677984e-24
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ dvt0w = 0
+ pvag = 1.2
+ dvt1w = 0
+ dvt2w = 0
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ rdsw = 100
+ ijthsfwd = 0.01
+ cigbacc = 0.32875
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ tnoimod = 0
+ tnoia = 0
+ ijthsrev = 0.01
+ cigbinv = 0.006
+ peta0 = 0
+ rshg = 15.6
+ wketa = -2.2122195e-8
+ wtvfbsdoff = 0
+ tpbsw = 0.0019
+ toxref = 3e-9
+ cjswd = 8.2e-11
+ cjsws = 8.2e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ version = 4.5
+ ltvfbsdoff = 0
+ tempmod = 0
+ ppdiblc2 = 1.7501102e-15
+ tnom = 25
+ aigbacc = 0.02
+ tvfbsdoff = 0.022
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ ltvoff = 1.3913801e-9
+ ags = 0.33766657
+ scref = 1e-6
+ cjd = 0.001357
+ cit = 0.00059502911
+ cjs = 0.001357
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 9.8024918e-9
+ pigcd = 2.621
+ k3b = 1.9326
+ aigsd = 0.010772818
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ ptvfbsdoff = 0
+ aigbinv = 0.0163
+ lvoff = -5.0132203e-10
+ wags = 3.8484036e-7
+ lku0we = 2.5e-11
+ pkvth0we = -1.3e-19
+ la0 = 3.6355951e-7
+ epsrox = 3.9
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.052738453
+ kt1 = -0.19312528
+ lk2 = -1.4722356e-8
+ kt2 = -0.039065148
+ wcit = 3.184653e-10
+ lvsat = 0
+ llc = 0
+ lln = 1
+ lu0 = -1.7516993e-9
+ mjd = 0.26
+ lvth0 = -8.2158156e-9
+ lua = -1.1159069e-16
+ mjs = 0.26
+ lub = -2.3732546e-26
+ luc = -2.9405776e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ voff = -0.14601446
+ njs = 1.02
+ pa0 = -3.8856002e-13
+ nsd = 1e+20
+ delta = 0.007595625
+ acde = 0.4
+ pbd = 0.52
+ wvfbsdoff = 0
+ pat = -8.5362363e-10
+ pbs = 0.52
+ rdsmod = 0
+ pk2 = 1.1847359e-15
+ lvfbsdoff = 0
+ laigc = -3.3762752e-11
+ pu0 = 1.2968191e-16
+ vfbsdoff = 0.02
+ igbmod = 1
+ prt = 0
+ pua = 2.9945529e-23
+ pub = -3.9782718e-32
+ puc = 6.3626704e-24
+ pud = 0
+ vsat = 102889.02
+ wint = 0
+ rnoia = 0
+ rnoib = 0
+ vth0 = 0.42537959
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 6.6639379e-10
+ ub1 = 1.1665789e-19
+ uc1 = 5.9635906e-11
+ wkt1 = -3.3221037e-8
+ wkt2 = -8.3325526e-9
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ tpb = 0.0014
+ wmax = 5.4e-7
+ wa0 = 7.714643e-7
+ aigc = 0.01167393
+ wmin = 2.7e-7
+ ute = -1
+ wat = 0.0079246317
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -8.8268726e-10
+ pbswgd = 0.95
+ pketa = 1.3732256e-14
+ poxedge = 1
+ pbswgs = 0.95
+ ngate = 8e+20
+ wlc = 0
+ wln = 1
+ wu0 = -1.2619767e-9
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -1.218412e-16
+ wub = 9.5438468e-26
+ wuc = -2.0432641e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ ngcon = 1
+ paramchk = 1
+ wpclm = 9.3989653e-8
+ igcmod = 1
+ binunit = 2
+ wua1 = 4.4082452e-17
+ wub1 = -1.420039e-25
+ wuc1 = -1.718815e-17
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ bigc = 0.001442
+ wwlc = 0
+ cdsc = 0
+ ijthdfwd = 0.01
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ permod = 1
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ ijthdrev = 0.01
+ tvoff = -0.0014023534
+ lpdiblc2 = -7.3119259e-9
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ voffcv = -0.16942
+ wpemod = 1
+ k2we = 5e-5
+ ku0we = -0.0007
+ dsub = 0.75
+ dtox = 2.7e-10
+ beta0 = 13
+ leta0 = 0
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ njtsswg = 9
+ lkvth0we = -2e-12
+ eta0 = 0.24044444
+ etab = -0.28088889
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.039504569
+ pdiblcb = -0.3
+ tpbswg = 0.0009
+ acnqsmod = 0
+ dmcgt = 0
+ tcjsw = 0.000357
+ rbodymod = 0
+ ptvoff = -5.8159511e-16
+ bigbacc = 0.002588
+ waigsd = 3.1113143e-12
+ bigsd = 0.00125
+ a0 = 0.37817284
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 204899.36
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.02255059
+ k3 = -1.8419
+ em = 1000000.0
+ kvth0we = 0.00018
+ diomod = 1
+ ll = 0
+ lw = 0
+ u0 = 0.017332646
+ w0 = 0
+ wvoff = 1.6411259e-8
+ ua = -1.8479686e-9
+ ub = 2.1067376e-18
+ uc = 1.1966909e-10
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 6e-9
+ lintnoi = -1.5e-8
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 2.82e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.82e-10
+ bigbinv = 0.004953
+ wvsat = -0.0028059037
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ wvth0 = -2.1299761e-8
+ wpdiblc2 = -3.7127843e-9
+ waigc = 2.313153e-11
+ mjswgd = 0.85
+ mjswgs = 0.85
+ lketa = -4.8021757e-8
+ tcjswg = 0.001
+ xpart = 1
+ pvfbsdoff = 0
+ keta = 0.03621471
+ egidl = 0.29734
+ wkvth0we = 2e-12
+ lags = 4.1799271e-7
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 3.7698897e-10
+ trnqsmod = 0
+ kt1l = 0
+ nfactor = 1
+ lint = 6.5375218e-9
+ fprout = 300
+ lkt1 = -1.6253643e-8
+ lkt2 = -1.6288295e-8
+ xrcrg1 = 12
+ xrcrg2 = 1
+ lmax = 8.9908e-7
+ lmin = 4.4908e-7
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ rgatemod = 0
+ wtvoff = 9.3241971e-10
+ pvoff = -4.5972513e-15
+ minv = -0.3
+ tnjtsswg = 1
+ lua1 = 4.5439491e-17
+ lub1 = -2.6809927e-25
+ luc1 = 3.3118724e-18
+ cdscb = 0
+ cdscd = 0
+ nigbacc = 10
+ ndep = 1e+18
+ pvsat = 0
+ wk2we = 5e-12
+ pvth0 = 5.9609158e-15
+ lwlc = 0
+ drout = 0.56
+ moin = 5.1
+ capmod = 2
+ paigc = -4.5341069e-18
+ nigc = 3.083
+ voffl = 0
+ wku0we = 2e-11
+ nigbinv = 10
+ mobmod = 0
+ weta0 = -1.1162667e-8
+ wetab = 2.2325333e-8
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ pags = -2.4281917e-13
+ cgidl = 0.22
+ )

.model nch_tt_28 nmos (
+ level = 54
+ wuc1 = -1.3268706e-17
+ bigc = 0.001442
+ ppclm = -7.9196439e-14
+ wwlc = 0
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ cdsc = 0
+ bigbacc = 0.002588
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ wtvfbsdoff = 0
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ kvth0we = 0.00018
+ dmcgt = 0
+ tcjsw = 0.000357
+ wkvth0we = 2e-12
+ lintnoi = -1.5e-8
+ ltvfbsdoff = 0
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ trnqsmod = 0
+ toxref = 3e-9
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ bigsd = 0.00125
+ wvoff = 5.1767953e-9
+ k2we = 5e-5
+ dsub = 0.75
+ wvsat = -0.0054199005
+ dtox = 2.7e-10
+ ptvfbsdoff = 0
+ wvth0 = -3.6869543e-9
+ rgatemod = 0
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ tnjtsswg = 1
+ waigc = -1.6608588e-12
+ ltvoff = -7.6859018e-11
+ eta0 = 0.24044444
+ etab = -0.28088889
+ lketa = -5.7215427e-9
+ nfactor = 1
+ xpart = 1
+ pvfbsdoff = 0
+ lku0we = 2.5e-11
+ egidl = 0.29734
+ epsrox = 3.9
+ rdsmod = 0
+ igbmod = 1
+ nigbacc = 10
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ pbswgd = 0.95
+ pbswgs = 0.95
+ igcmod = 1
+ nigbinv = 10
+ pvoff = 3.4591262e-16
+ cdscb = 0
+ cdscd = 0
+ pvsat = 1.1501586e-9
+ wk2we = 5e-12
+ pvth0 = -1.7887192e-15
+ drout = 0.56
+ paigc = 6.374544e-18
+ ijthsfwd = 0.01
+ paigsd = 2.2627557e-23
+ voffl = 0
+ fnoimod = 1
+ eigbinv = 1.1
+ keta = -0.05992214
+ weta0 = -1.1162667e-8
+ wetab = 2.2325333e-8
+ permod = 1
+ lpclm = 1.4504842e-7
+ lags = 5.906061e-7
+ jswd = 1.28e-13
+ ijthsrev = 0.01
+ jsws = 1.28e-13
+ lcit = 9.3365571e-11
+ cgidl = 0.22
+ kt1l = 0
+ lint = 9.7879675e-9
+ voffcv = -0.16942
+ wpemod = 1
+ lkt1 = 8.8603069e-9
+ lkt2 = -2.5638367e-9
+ lmax = 4.4908e-7
+ cigbacc = 0.32875
+ pbswd = 0.8
+ pbsws = 0.8
+ lmin = 2.1577e-7
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ ppdiblc2 = -5.242001e-17
+ tnoimod = 0
+ minv = -0.3
+ lua1 = -4.6794128e-17
+ lub1 = -3.2889654e-26
+ luc1 = -2.1335001e-17
+ pdits = 0
+ ndep = 1e+18
+ cigsd = 0.069865
+ cigbinv = 0.006
+ dvt0w = 0
+ lwlc = 0
+ dvt1w = 0
+ dvt2w = 0
+ moin = 5.1
+ nigc = 3.083
+ tpbswg = 0.0009
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ version = 4.5
+ tempmod = 0
+ pkvth0we = -1.3e-19
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ tnoia = 0
+ pags = 1.2428184e-13
+ peta0 = 0
+ ptvoff = -1.5558646e-16
+ aigbacc = 0.02
+ ntox = 1
+ pcit = -8.9847229e-18
+ pclm = 1.1798023
+ waigsd = 3.1112628e-12
+ wketa = 2.3981389e-8
+ vfbsdoff = 0.02
+ tpbsw = 0.0019
+ cjswd = 8.2e-11
+ cjsws = 8.2e-11
+ diomod = 1
+ mjswd = 0.11
+ phin = 0.15
+ mjsws = 0.11
+ agidl = 9.41e-8
+ pditsd = 0
+ pditsl = 0
+ aigbinv = 0.0163
+ pkt1 = -1.2500052e-14
+ pkt2 = -7.0784646e-16
+ cjswgd = 2.82e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.82e-10
+ paramchk = 1
+ ags = -0.054636584
+ cjd = 0.001357
+ tvfbsdoff = 0.022
+ cit = 0.0012396277
+ cjs = 0.001357
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 1.30529375e-8
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ rbdb = 50
+ pua1 = 1.8291934e-23
+ prwb = 0
+ prwg = 0
+ pub1 = -6.5524188e-33
+ puc1 = 5.143243e-24
+ mjswgd = 0.85
+ mjswgs = 0.85
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ tcjswg = 0.001
+ rdsw = 100
+ scref = 1e-6
+ ijthdfwd = 0.01
+ la0 = -6.0902319e-7
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.015036938
+ kt1 = -0.25020244
+ lk2 = -1.0681005e-8
+ kt2 = -0.070257098
+ pigcd = 2.621
+ llc = -1.18e-13
+ lln = 0.7
+ aigsd = 0.010772818
+ lu0 = -7.0583626e-10
+ mjd = 0.26
+ lua = -1.8564943e-17
+ mjs = 0.26
+ lub = -5.2748233e-26
+ luc = -4.2757753e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 2.2627554e-14
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 2.5637001e-9
+ poxedge = 1
+ pbs = 0.52
+ pk2 = 8.6250113e-16
+ lvoff = -7.1474494e-9
+ a0 = 2.5885881
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ pu0 = 5.1138272e-17
+ at = 119214.09
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.013365692
+ k3 = -1.8419
+ em = 1000000.0
+ prt = 0
+ pua = 5.6394132e-24
+ pub = -7.710339e-34
+ puc = -1.5613012e-24
+ pud = 0
+ ll = -1.18e-13
+ lw = 0
+ u0 = 0.014955684
+ w0 = 0
+ ua = -2.0593908e-9
+ ub = 2.1726824e-18
+ uc = 6.2555449e-11
+ ud = 0
+ wl = 0
+ rsh = 17.5
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 6e-9
+ tcj = 0.00076
+ ua1 = 8.7601565e-10
+ lvsat = -0.0041672412
+ ub1 = -4.1790941e-19
+ uc1 = 1.1565153e-10
+ binunit = 2
+ lvth0 = 1.474398e-9
+ ijthdrev = 0.01
+ tpb = 0.0014
+ wvfbsdoff = 0
+ wa0 = -1.6305293e-7
+ lvfbsdoff = 0
+ ute = -1
+ wat = 0.00015798693
+ delta = 0.007595625
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -1.5033038e-10
+ laigc = -3.7429738e-11
+ wlc = 0
+ wln = 1
+ rshg = 15.6
+ wu0 = -1.0834684e-9
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -6.6600022e-17
+ wub = 6.7755498e-27
+ wuc = -2.4236148e-18
+ wud = 0
+ lpdiblc2 = -4.2799755e-9
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ rnoia = 0
+ rnoib = 0
+ fprout = 300
+ xrcrg1 = 12
+ xrcrg2 = 1
+ pketa = -6.5533207e-15
+ ngate = 8e+20
+ ngcon = 1
+ wpclm = 2.7398156e-7
+ wtvoff = -3.5781771e-11
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ tnom = 25
+ jswgs = 1.28e-13
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ lkvth0we = -2e-12
+ capmod = 2
+ wku0we = 2e-11
+ mobmod = 0
+ acnqsmod = 0
+ wags = -4.4948013e-7
+ wcit = 7.5116891e-11
+ rbodymod = 0
+ voff = -0.13090963
+ acde = 0.4
+ tvoff = 0.0019345538
+ njtsswg = 9
+ vsat = 112360.02
+ wint = 0
+ xjbvd = 1
+ xjbvs = 1
+ vth0 = 0.40335638
+ lk2we = -1.5e-12
+ wkt1 = 6.1264548e-9
+ wkt2 = -1.5558741e-9
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ wmax = 5.4e-7
+ laigsd = -8.1983894e-17
+ aigc = 0.011682264
+ wmin = 2.7e-7
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.032613772
+ pdiblcb = -0.3
+ ku0we = -0.0007
+ beta0 = 13
+ leta0 = 0
+ wua1 = -5.7419768e-17
+ wpdiblc2 = 3.8387521e-10
+ wub1 = -1.6295463e-26
+ )

.model nch_tt_29 nmos (
+ level = 54
+ keta = 0.0092481698
+ aigbinv = 0.0163
+ tnoia = 0
+ ijthdrev = 0.01
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = -1.3537106e-11
+ peta0 = 0
+ ptvfbsdoff = 0
+ kt1l = 0
+ wketa = -2.0169501e-8
+ toxref = 3e-9
+ lpdiblc2 = -9.0824285e-10
+ tpbsw = 0.0019
+ ags = 2.7444444
+ cjswd = 8.2e-11
+ cjsws = 8.2e-11
+ lint = 9.7879675e-9
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ cjd = 0.001357
+ cit = 0.0017462755
+ cjs = 0.001357
+ clc = 1e-7
+ cle = 0.6
+ lkt1 = -2.5262126e-9
+ bvd = 8.7
+ lkt2 = -3.9513595e-9
+ bvs = 8.7
+ lmax = 2.1577e-7
+ dlc = 1.30529375e-8
+ lmin = 9e-8
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ poxedge = 1
+ tvfbsdoff = 0.022
+ la0 = -2.075695e-7
+ minv = -0.3
+ jsd = 6.11e-7
+ ltvoff = 5.8839234e-11
+ jss = 6.11e-7
+ lat = -0.0015937311
+ lua1 = -5.8912951e-18
+ lub1 = -2.9377439e-26
+ luc1 = 1.0640856e-17
+ kt1 = -0.1962379
+ lk2 = -3.2022951e-9
+ kt2 = -0.063681161
+ llc = -1.18e-13
+ binunit = 2
+ lln = 0.7
+ lu0 = -2.5551767e-10
+ mjd = 0.26
+ lua = 5.2959027e-17
+ mjs = 0.26
+ lub = -7.97606935e-26
+ luc = -8.8267893e-18
+ lud = 0
+ lwc = 0
+ ndep = 1e+18
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ lkvth0we = -2e-12
+ njs = 1.02
+ pa0 = 1.0407708e-13
+ nsd = 1e+20
+ lwlc = 0
+ pbd = 0.52
+ pat = -3.7161951e-10
+ pbs = 0.52
+ pk2 = -9.7578421e-17
+ moin = 5.1
+ pu0 = 1.8260797e-17
+ prt = 0
+ pua = -7.1102082e-24
+ pub = 9.57267e-33
+ puc = 7.19078e-25
+ pud = 0
+ scref = 1e-6
+ nigc = 3.083
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 6.8216336e-10
+ pigcd = 2.621
+ ub1 = -4.3455498e-19
+ uc1 = -3.5892821e-11
+ aigsd = 0.010772818
+ tpb = 0.0014
+ lku0we = 2.5e-11
+ wa0 = -5.4906963e-7
+ acnqsmod = 0
+ ute = -1
+ wat = 0.014069454
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 4.3998097e-9
+ epsrox = 3.9
+ lvoff = 2.33236653e-9
+ wlc = 0
+ wln = 1
+ wu0 = -9.2765099e-10
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -6.1752756e-18
+ wub = -4.2246744000000004e-26
+ wuc = -1.3231099e-17
+ wud = 0
+ wwc = 0
+ noff = 2.7195
+ wwl = 0
+ wwn = 1
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ lvsat = -0.00045734827
+ rbodymod = 0
+ rdsmod = 0
+ wvfbsdoff = 0
+ lvth0 = -1.2194990599999998e-8
+ lvfbsdoff = 0
+ igbmod = 1
+ delta = 0.007595625
+ laigc = 2.6175146e-12
+ ntox = 1
+ pcit = 7.8208248e-18
+ jtsswgd = 2.3e-7
+ pclm = 2.3689724
+ jtsswgs = 2.3e-7
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ rnoia = 0
+ rnoib = 0
+ pbswgd = 0.95
+ pbswgs = 0.95
+ phin = 0.15
+ pketa = 2.762517e-15
+ ngate = 8e+20
+ igcmod = 1
+ ngcon = 1
+ pkt1 = 6.6516645e-16
+ pkt2 = 9.3582987e-16
+ wpclm = -2.0834879e-7
+ wpdiblc2 = 1.3111248e-10
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ rbdb = 50
+ pua1 = 1.9734917e-24
+ prwb = 0
+ prwg = 0
+ pub1 = -5.2222001e-33
+ puc1 = -4.0873907e-24
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ njtsswg = 9
+ paigsd = -9.4615512e-24
+ rdsw = 100
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ permod = 1
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.016633997
+ pdiblcb = -0.3
+ wkvth0we = 2e-12
+ trnqsmod = 0
+ tvoff = 0.0012914341
+ rshg = 15.6
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ voffcv = -0.16942
+ wpemod = 1
+ bigbacc = 0.002588
+ ku0we = -0.0007
+ kvth0we = 0.00018
+ beta0 = 13
+ leta0 = 0
+ rgatemod = 0
+ lintnoi = -1.5e-8
+ tnjtsswg = 1
+ tnom = 25
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ ppclm = 2.2575265e-14
+ vtsswgs = 4.2
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ tpbswg = 0.0009
+ dmcgt = 0
+ wags = 1.3953333e-7
+ tcjsw = 0.000357
+ wcit = -4.5302538e-12
+ ptvoff = 2.7225835e-17
+ voff = -0.175837897
+ waigsd = 3.1114149e-12
+ acde = 0.4
+ vsat = 94777.65030000001
+ wint = 0
+ bigsd = 0.00125
+ vth0 = 0.468140454
+ diomod = 1
+ wkt1 = -5.6267946e-8
+ wkt2 = -9.3458092e-9
+ wmax = 5.4e-7
+ aigc = 0.011492467
+ wmin = 2.7e-7
+ nfactor = 1
+ pditsd = 0
+ pditsl = 0
+ wvoff = 8.989216699999998e-9
+ cjswgd = 2.82e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.82e-10
+ wvsat = -0.0005775380999999999
+ wvth0 = -1.7125728000000003e-8
+ wua1 = 1.991882e-17
+ wub1 = -2.2599817e-26
+ wuc1 = 3.0478373e-17
+ waigc = 3.9031408e-11
+ bigc = 0.001442
+ mjswgd = 0.85
+ mjswgs = 0.85
+ wwlc = 0
+ tcjswg = 0.001
+ nigbacc = 10
+ lketa = -2.0316478e-8
+ cdsc = 0
+ ijthsfwd = 0.01
+ cgbo = 0
+ xpart = 1
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ pvfbsdoff = 0
+ xtid = 3
+ xtis = 3
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ egidl = 0.29734
+ nigbinv = 10
+ ijthsrev = 0.01
+ fprout = 300
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ fnoimod = 1
+ k2we = 5e-5
+ wtvoff = -9.0219076e-10
+ eigbinv = 1.1
+ dsub = 0.75
+ dtox = 2.7e-10
+ ppdiblc2 = 9.1292629e-19
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ pvoff = -4.585090499999998e-16
+ a0 = 0.68596391
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 55502.213
+ cf = 8.15e-11
+ cdscb = 0
+ cdscd = 0
+ ef = 1.0
+ k1 = 0.274
+ k2 = -0.02207843
+ k3 = -1.8419
+ em = 1000000.0
+ ll = -1.18e-13
+ lw = 0
+ u0 = 0.012821473
+ pvsat = 1.2842156000000008e-10
+ w0 = 0
+ ua = -2.398367e-9
+ ub = 2.300703286e-18
+ uc = 8.4124236e-11
+ ud = 0
+ wk2we = 5e-12
+ capmod = 2
+ wl = 0
+ wr = 1
+ pvth0 = 1.0468620000000002e-15
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ eta0 = 0.24044444
+ xw = 6e-9
+ drout = 0.56
+ etab = -0.28088889
+ wku0we = 2e-11
+ paigc = -2.2115244e-18
+ mobmod = 0
+ voffl = 0
+ cigbacc = 0.32875
+ weta0 = -1.1162667e-8
+ wetab = 2.2325333e-8
+ pkvth0we = -1.3e-19
+ lpclm = -1.0586647e-7
+ tnoimod = 0
+ cgidl = 0.22
+ vfbsdoff = 0.02
+ cigbinv = 0.006
+ laigsd = 3.4280989e-17
+ pbswd = 0.8
+ pbsws = 0.8
+ paramchk = 1
+ version = 4.5
+ wtvfbsdoff = 0
+ tempmod = 0
+ pdits = 0
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ cigsd = 0.069865
+ ltvfbsdoff = 0
+ dvt0w = 0
+ aigbacc = 0.02
+ dvt1w = 0
+ dvt2w = 0
+ ijthdfwd = 0.01
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ )

.model nch_tt_30 nmos (
+ level = 54
+ keta = -0.29566775
+ aigbinv = 0.0163
+ tnoia = 0
+ ijthdrev = 0.01
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 1.7434428e-10
+ peta0 = -9.3037135e-16
+ ptvfbsdoff = 0
+ petab = -1.2138265e-15
+ kt1l = 0
+ wketa = -4.7865407e-8
+ toxref = 3e-9
+ lpdiblc2 = 8.2379047e-15
+ tpbsw = 0.0019
+ ags = 2.7444444
+ cjswd = 8.2e-11
+ cjsws = 8.2e-11
+ lint = 0
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ cjd = 0.001357
+ cit = -0.00025246267
+ cjs = 0.001357
+ clc = 1e-7
+ cle = 0.6
+ lkt1 = -8.4950836e-9
+ bvd = 8.7
+ lkt2 = 3.8424987e-10
+ bvs = 8.7
+ lmax = 9e-8
+ dlc = 3.26497e-9
+ lmin = 5.4e-8
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ poxedge = 1
+ tvfbsdoff = 0.022
+ la0 = 3.9829889e-7
+ minv = -0.3
+ jsd = 6.11e-7
+ ltvoff = -2.7237524e-10
+ jss = 6.11e-7
+ lat = 0.00528560498
+ lua1 = -1.2736334e-17
+ lub1 = 1.6085594e-26
+ luc1 = 1.132730421e-17
+ kt1 = -0.13273927
+ lk2 = 1.0502722e-9
+ kt2 = -0.10980467
+ llc = 0
+ binunit = 2
+ lln = 1
+ lu0 = -2.0475966e-10
+ mjd = 0.26
+ lua = -7.6887484e-18
+ mjs = 0.26
+ lub = 6.3606825e-27
+ luc = -3.2720592999999998e-18
+ lud = 0
+ lwc = 0
+ ndep = 1e+18
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ lkvth0we = -2e-12
+ njs = 1.02
+ pa0 = -1.1411036e-13
+ nsd = 1e+20
+ lwlc = 0
+ pbd = 0.52
+ pat = -1.7320563000000002e-9
+ pbs = 0.52
+ pk2 = -3.7289588e-16
+ moin = 5.1
+ pu0 = 7.2584501e-17
+ prt = 0
+ pua = 1.3044266e-23
+ pub = -1.13966382e-32
+ puc = 2.3653651e-24
+ pud = 0
+ scref = 1e-6
+ nigc = 3.083
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 7.5498293e-10
+ pigcd = 2.621
+ ub1 = -9.1820427e-19
+ uc1 = -4.319545900000001e-11
+ aigsd = 0.010772818
+ tpb = 0.0014
+ lku0we = 2.5e-11
+ wa0 = 1.7720733e-6
+ acnqsmod = 0
+ ute = -1
+ wat = 0.028542186400000003
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 7.3287188e-9
+ epsrox = 3.9
+ lvoff = -3.2511799e-9
+ wlc = 0
+ wln = 1
+ wu0 = -1.5055627e-9
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -2.2058458e-16
+ wub = 1.80830997e-25
+ wuc = -3.0744792e-17
+ wud = 0
+ wwc = 0
+ noff = 2.7195
+ wwl = 0
+ wwn = 1
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ lvsat = 0.0032456743
+ rbodymod = 0
+ rdsmod = 0
+ wvfbsdoff = 0
+ lvth0 = 3.589724300000001e-9
+ lvfbsdoff = 0
+ igbmod = 1
+ delta = 0.007595625
+ laigc = -3.0244582e-11
+ ntox = 1
+ pcit = -1.9457676e-17
+ jtsswgd = 2.3e-7
+ pclm = 1.7776553
+ jtsswgs = 2.3e-7
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ rnoia = 0
+ rnoib = 0
+ pbswgd = 0.95
+ pbswgs = 0.95
+ phin = 0.15
+ pketa = 5.3659323e-15
+ ngate = 8e+20
+ igcmod = 1
+ ngcon = 1
+ pkt1 = 5.1065068e-15
+ pkt2 = -5.9202052e-16
+ wpclm = 4.3365813e-8
+ wpdiblc2 = 1.4083642e-10
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ rbdb = 50
+ pua1 = 4.1884121e-24
+ prwb = 0
+ prwg = 0
+ pub1 = -9.7869988e-33
+ puc1 = -6.8508479999999965e-25
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ njtsswg = 9
+ rdsw = 100
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ permod = 1
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.0069717513
+ pdiblcb = -0.3
+ wkvth0we = 2e-12
+ trnqsmod = 0
+ tvoff = 0.0048149924
+ rshg = 15.6
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ voffcv = -0.16942
+ wpemod = 1
+ bigbacc = 0.002588
+ ku0we = -0.0007
+ kvth0we = 0.00018
+ beta0 = 13
+ leta0 = 2.0040249e-8
+ rgatemod = 0
+ letab = -2.6551319e-8
+ lintnoi = -1.5e-8
+ tnjtsswg = 1
+ tnom = 25
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ ppclm = -1.085908e-15
+ vtsswgs = 4.2
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ tpbswg = 0.0009
+ dmcgt = 0
+ wags = 1.3953333e-7
+ tcjsw = 0.000357
+ wcit = 2.8566656e-10
+ ptvoff = 9.0058483e-17
+ voff = -0.116438471
+ waigsd = 3.1113143e-12
+ acde = 0.4
+ vsat = 55383.79300000001
+ wint = 0
+ bigsd = 0.00125
+ vth0 = 0.300217953
+ diomod = 1
+ wkt1 = -1.0351625e-7
+ wkt2 = 6.9079183e-9
+ wmax = 5.4e-7
+ aigc = 0.011842064
+ wmin = 2.7e-7
+ nfactor = 1
+ pditsd = 0
+ pditsl = 0
+ wvoff = 4.307686799999997e-9
+ cjswgd = 2.82e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.82e-10
+ wvsat = 0.005122454499999998
+ wvth0 = -6.7257771000000035e-9
+ wua1 = -3.6441631e-18
+ wub1 = 2.5961869999999995e-26
+ wuc1 = -5.7163699999999976e-18
+ waigc = 4.5087747e-12
+ bigc = 0.001442
+ mjswgd = 0.85
+ mjswgs = 0.85
+ wwlc = 0
+ tcjswg = 0.001
+ nigbacc = 10
+ lketa = 8.345618e-9
+ cdsc = 0
+ ijthsfwd = 0.01
+ cgbo = 0
+ xpart = 1
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ pvfbsdoff = 0
+ xtid = 3
+ xtis = 3
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ egidl = 0.29734
+ nigbinv = 10
+ ijthsrev = 0.01
+ fprout = 300
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ fnoimod = 1
+ k2we = 5e-5
+ wtvoff = -1.5706231e-9
+ eigbinv = 1.1
+ dsub = 0.75
+ dtox = 2.7e-10
+ ppdiblc2 = -1.1241984e-21
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ pvoff = -1.8445117999999986e-17
+ a0 = -5.7594444
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = -17682.2125
+ cf = 8.15e-11
+ cdscb = 0
+ cdscd = 0
+ ef = 1.0
+ k1 = 0.274
+ k2 = -0.067318509
+ k3 = -1.8419
+ em = 1000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.012281494
+ pvsat = -4.073777999999999e-10
+ w0 = 0
+ ua = -1.7531779e-9
+ ub = 1.3845184050000002e-18
+ uc = 2.5031363e-11
+ ud = 0
+ wk2we = 5e-12
+ capmod = 2
+ wl = 0
+ wr = 1
+ pvth0 = 6.926666000000025e-17
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ eta0 = 0.027250304
+ xw = 6e-9
+ drout = 0.56
+ etab = 0.001571952
+ wku0we = 2e-11
+ paigc = 1.0336032e-18
+ mobmod = 0
+ voffl = 0
+ cigbacc = 0.32875
+ weta0 = -1.2650991e-9
+ wetab = 3.5238381e-8
+ pkvth0we = -1.3e-19
+ lpclm = -5.0282662e-8
+ tnoimod = 0
+ cgidl = 0.22
+ vfbsdoff = 0.02
+ cigbinv = 0.006
+ pbswd = 0.8
+ pbsws = 0.8
+ paramchk = 1
+ version = 4.5
+ wtvfbsdoff = 0
+ tempmod = 0
+ pdits = 0
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ cigsd = 0.069865
+ ltvfbsdoff = 0
+ dvt0w = 0
+ aigbacc = 0.02
+ dvt1w = 0
+ dvt2w = 0
+ ijthdfwd = 0.01
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ )

.model nch_tt_31 nmos (
+ level = 54
+ nigbacc = 10
+ wvoff = 2.6164685300000083e-9
+ wvsat = 0.023374044200000006
+ wvth0 = -3.0287313e-8
+ ltvoff = 2.6647905e-10
+ waigc = 1.8753243e-11
+ tnom = 25
+ nigbinv = 10
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ lketa = -2.3617222e-8
+ pvfbsdoff = 0
+ xpart = 1
+ lku0we = 2.5e-11
+ epsrox = 3.9
+ egidl = 0.29734
+ fnoimod = 1
+ pkvth0we = -1.3e-19
+ wags = 1.3953333e-7
+ rdsmod = 0
+ eigbinv = 1.1
+ wcit = 3.7128934e-10
+ igbmod = 1
+ voff = -0.07382279000000001
+ acde = 0.4
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ vfbsdoff = 0.02
+ vsat = 35732.98
+ pbswgd = 0.95
+ pbswgs = 0.95
+ wint = 0
+ vth0 = 0.31962439000000004
+ wkt1 = -1.6694349e-8
+ wkt2 = -2.0876247e-8
+ wmax = 5.4e-7
+ igcmod = 1
+ aigc = 0.011696193
+ wmin = 2.7e-7
+ paramchk = 1
+ cigbacc = 0.32875
+ wua1 = -1.1132499e-16
+ wub1 = 7.746802000000003e-26
+ wuc1 = 1.6593491000000002e-16
+ pvoff = 7.964544000000045e-17
+ bigc = 0.001442
+ cdscb = 0
+ cdscd = 0
+ tnoimod = 0
+ wwlc = 0
+ pvsat = -1.4659699999999999e-9
+ wk2we = 5e-12
+ pvth0 = 1.4358358e-15
+ drout = 0.56
+ paigsd = 1.7624612e-23
+ cdsc = 0
+ paigc = 2.0742404e-19
+ cigbinv = 0.006
+ ijthdfwd = 0.01
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ voffl = 0
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ permod = 1
+ weta0 = -1.2005104e-7
+ wetab = 5.6750807e-8
+ lpclm = 5.458214e-8
+ version = 4.5
+ tempmod = 0
+ ijthdrev = 0.01
+ cgidl = 0.22
+ voffcv = -0.16942
+ wpemod = 1
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ aigbacc = 0.02
+ pbswd = 0.8
+ pbsws = 0.8
+ k2we = 5e-5
+ dsub = 0.75
+ dtox = 2.7e-10
+ aigbinv = 0.0163
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ pdits = 0
+ cigsd = 0.069865
+ lkvth0we = -2e-12
+ eta0 = 1.0176617
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ etab = -1.3959412
+ tpbswg = 0.0009
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ acnqsmod = 0
+ tnoia = 0
+ ptvoff = -4.401556e-18
+ poxedge = 1
+ rbodymod = 0
+ ags = 2.7444444
+ waigsd = 3.1110104e-12
+ peta0 = 5.9592132e-15
+ cjd = 0.001357
+ cit = -0.0053709179
+ cjs = 0.001357
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ petab = -2.4615472e-15
+ dlc = 3.26497e-9
+ binunit = 2
+ wketa = -5.877032e-8
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ diomod = 1
+ tpbsw = 0.0019
+ cjswd = 8.2e-11
+ cjsws = 8.2e-11
+ mjswd = 0.11
+ pditsd = 0
+ pditsl = 0
+ mjsws = 0.11
+ agidl = 9.41e-8
+ cjswgd = 2.82e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.82e-10
+ la0 = -1.4097724e-8
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.0007194377000000001
+ kt1 = -0.39757001
+ lk2 = 7.4338958e-10
+ kt2 = -0.14677127
+ llc = 0
+ lln = 1
+ lu0 = 5.0770058e-10
+ mjd = 0.26
+ lua = 6.4763643e-17
+ mjs = 0.26
+ lub = -2.3096342000000002e-26
+ luc = -1.0931136000000001e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = -1.7333804e-13
+ nsd = 1e+20
+ pbd = 0.52
+ pat = -4.378947099999998e-10
+ tvfbsdoff = 0.022
+ pbs = 0.52
+ pk2 = -1.0803308e-16
+ wpdiblc2 = 1.4081704e-10
+ pu0 = -4.6127483e-17
+ prt = 0
+ pua = -2.1774501e-24
+ pub = -5.473259300000002e-33
+ puc = 4.761497700000001e-24
+ pud = 0
+ mjswgd = 0.85
+ mjswgs = 0.85
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 1.4910078e-9
+ ub1 = -1.7286540799999999e-18
+ uc1 = -4.0168785999999996e-10
+ tpb = 0.0014
+ tcjswg = 0.001
+ wa0 = 2.7932403e-6
+ ute = -1
+ wat = 0.006229054600000004
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 2.7621189e-9
+ wlc = 0
+ wln = 1
+ wu0 = 5.411956e-10
+ jtsswgd = 2.3e-7
+ xgl = -1.09e-8
+ jtsswgs = 2.3e-7
+ xgw = 0
+ wua = 4.1858808e-17
+ wub = 7.870378029999999e-26
+ wuc = -7.2057435e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ scref = 1e-6
+ pigcd = 2.621
+ aigsd = 0.010772819
+ keta = 0.2554158
+ lvoff = -5.722889800000002e-9
+ wkvth0we = 2e-12
+ wvfbsdoff = 0
+ lvsat = 0.004385421569999999
+ lvfbsdoff = 0
+ lvth0 = 2.4641506e-9
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 4.7121469e-10
+ trnqsmod = 0
+ delta = 0.007595625
+ laigc = -2.1784105e-11
+ kt1l = 0
+ fprout = 300
+ xrcrg1 = 12
+ xrcrg2 = 1
+ rnoia = 0
+ rnoib = 0
+ lint = 0
+ njtsswg = 9
+ lkt1 = 6.8650994e-9
+ lkt2 = 2.528313e-9
+ pketa = 5.998417e-15
+ ngate = 8e+20
+ lmax = 5.4e-8
+ lmin = 4.5e-8
+ wtvoff = 5.799816e-11
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ ngcon = 1
+ wpclm = 2.4669208e-7
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ ckappad = 0.6
+ ckappas = 0.6
+ rgatemod = 0
+ gbmin = 1e-12
+ pdiblc1 = 0
+ pdiblc2 = 0.0069718933
+ pdiblcb = -0.3
+ tnjtsswg = 1
+ minv = -0.3
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ lua1 = -5.5425775e-17
+ lub1 = 6.309168e-26
+ luc1 = 3.2119863e-17
+ capmod = 2
+ ndep = 1e+18
+ wku0we = 2e-11
+ lwlc = 0
+ moin = 5.1
+ mobmod = 0
+ nigc = 3.083
+ bigbacc = 0.002588
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ kvth0we = 0.00018
+ wtvfbsdoff = 0
+ lintnoi = -1.5e-8
+ bigbinv = 0.004953
+ tvoff = -0.0044755986
+ ntox = 1
+ vtsswgd = 4.2
+ pcit = -2.4423797e-17
+ vtsswgs = 4.2
+ pclm = -0.030358553
+ laigsd = -6.385731e-17
+ xjbvd = 1
+ a0 = 1.350842
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ xjbvs = 1
+ lk2we = -1.5e-12
+ at = 85853.00300000001
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = -0.062027428
+ k3 = -1.8419
+ em = 1000000.0
+ ltvfbsdoff = 0
+ ll = 0
+ lw = 0
+ u0 = -2.3029531e-6
+ w0 = 0
+ ua = -3.002357e-9
+ ub = 1.89239813e-18
+ uc = 1.5708441000000004e-10
+ ud = 0
+ phin = 0.15
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 6e-9
+ pkt1 = 7.083666e-17
+ pkt2 = 1.019461e-15
+ ku0we = -0.0007
+ beta0 = 13
+ leta0 = -3.7403611e-8
+ letab = 5.4504443e-8
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ ppclm = -1.2878832e-14
+ rbdb = 50
+ pua1 = 1.04339e-23
+ prwb = 0
+ prwg = 0
+ pub1 = -1.2774356e-32
+ puc1 = -1.0640858600000001e-23
+ rbpb = 50
+ rbpd = 50
+ dlcig = 2.5e-9
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ bgidl = 2320000000.0
+ ptvfbsdoff = 0
+ rdsw = 100
+ ijthsfwd = 0.01
+ nfactor = 1
+ dmcgt = 0
+ tcjsw = 0.000357
+ ijthsrev = 0.01
+ toxref = 3e-9
+ rshg = 15.6
+ bigsd = 0.00125
+ )

.model nch_tt_32 nmos (
+ level = 54
+ eta0 = -0.25440451
+ etab = -0.81370191
+ scref = 1e-6
+ lku0we = 2.5e-11
+ pigcd = 2.621
+ epsrox = 3.9
+ aigsd = 0.010772817
+ njtsswg = 9
+ lvoff = -6.3267068e-9
+ rdsmod = 0
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ igbmod = 1
+ lvsat = -0.0013704545999999999
+ ckappad = 0.6
+ ckappas = 0.6
+ lvth0 = 3.9667989999999906e-10
+ pdiblc1 = 0
+ pdiblc2 = 0.0069718933
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ pdiblcb = -0.3
+ delta = 0.007595625
+ laigc = 9.707156e-12
+ pbswgd = 0.95
+ pbswgs = 0.95
+ rnoia = 0
+ rnoib = 0
+ igcmod = 1
+ pketa = -6.053668000000001e-15
+ ngate = 8e+20
+ ngcon = 1
+ wpclm = 1.6305740000000013e-7
+ bigbacc = 0.002588
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ kvth0we = 0.00018
+ paigsd = -1.2154906e-23
+ lintnoi = -1.5e-8
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ ijthsfwd = 0.01
+ permod = 1
+ keta = -0.59506219
+ ijthsrev = 0.01
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 3.03749e-10
+ tvoff = 0.0034020192
+ kt1l = 0
+ voffcv = -0.16942
+ wpemod = 1
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ lint = 0
+ lkt1 = -1.8529946e-8
+ lkt2 = 1.0897551e-9
+ lmax = 4.5e-8
+ lmin = 3.6e-8
+ ku0we = -0.0007
+ nfactor = 1
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ beta0 = 13
+ leta0 = 2.4927632200000002e-8
+ letab = 2.5974719e-8
+ minv = -0.3
+ lua1 = 7.6118385e-17
+ lub1 = -1.2790425e-25
+ luc1 = -3.7246243e-17
+ ppclm = -8.780734400000002e-15
+ ndep = 1e+18
+ dlcig = 2.5e-9
+ lwlc = 0
+ tpbswg = 0.0009
+ bgidl = 2320000000.0
+ moin = 5.1
+ nigc = 3.083
+ nigbacc = 10
+ dmcgt = 0
+ pkvth0we = -1.3e-19
+ noff = 2.7195
+ tcjsw = 0.000357
+ ptvoff = -5.392468e-18
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ waigsd = 3.1116181e-12
+ nigbinv = 10
+ diomod = 1
+ ntox = 1
+ pcit = -3.4847791e-17
+ vfbsdoff = 0.02
+ pclm = 1.46768105
+ bigsd = 0.00125
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 2.82e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.82e-10
+ phin = 0.15
+ wvoff = 6.255152000000001e-9
+ paramchk = 1
+ pkt1 = 5.3710205e-15
+ pkt2 = -4.1883975e-17
+ wvsat = -0.026256236
+ wvth0 = -1.0572559e-8
+ fnoimod = 1
+ mjswgd = 0.85
+ mjswgs = 0.85
+ eigbinv = 1.1
+ waigc = 7.6854687e-11
+ tcjswg = 0.001
+ rbdb = 50
+ pua1 = -2.7889543e-23
+ prwb = 0
+ prwg = 0
+ pub1 = 4.5022459e-32
+ puc1 = 1.2190153e-23
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ pvfbsdoff = 0
+ lketa = 1.80561909e-8
+ ijthdfwd = 0.01
+ rdsw = 100
+ xpart = 1
+ egidl = 0.29734
+ cigbacc = 0.32875
+ ijthdrev = 0.01
+ fprout = 300
+ rshg = 15.6
+ xrcrg1 = 12
+ xrcrg2 = 1
+ tnoimod = 0
+ cigbinv = 0.006
+ wtvoff = 7.822084e-11
+ pvoff = -9.865003999999993e-17
+ version = 4.5
+ capmod = 2
+ tnom = 25
+ cdscb = 0
+ cdscd = 0
+ tempmod = 0
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ pvsat = 9.6591382e-10
+ wku0we = 2e-11
+ lkvth0we = -2e-12
+ wk2we = 5e-12
+ pvth0 = 4.698127899999999e-16
+ drout = 0.56
+ mobmod = 0
+ wtvfbsdoff = 0
+ paigc = -2.6395467e-18
+ aigbacc = 0.02
+ voffl = 0
+ acnqsmod = 0
+ ltvfbsdoff = 0
+ weta0 = 8.5615058e-8
+ wetab = 2.2270081e-8
+ wags = 1.3953333e-7
+ lpclm = -1.8821805999999992e-8
+ wcit = 5.840239e-10
+ rbodymod = 0
+ aigbinv = 0.0163
+ voff = -0.061499972999999986
+ cgidl = 0.22
+ acde = 0.4
+ laigsd = 4.4039511e-17
+ vsat = 153199.842
+ wint = 0
+ vth0 = 0.36181767099999995
+ wkt1 = -1.2486137e-7
+ wkt2 = 7.8385579e-10
+ wmax = 5.4e-7
+ aigc = 0.011053515
+ wmin = 2.7e-7
+ pbswd = 0.8
+ pbsws = 0.8
+ ptvfbsdoff = 0
+ wpdiblc2 = 1.4081704e-10
+ wua1 = 6.7078609e-16
+ wub1 = -1.1020589000000001e-24
+ wuc1 = -3.0000411e-16
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ poxedge = 1
+ bigc = 0.001442
+ pdits = 0
+ wwlc = 0
+ cigsd = 0.069865
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ binunit = 2
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ ags = 2.7444444
+ cgsl = 3.31989e-12
+ pk2we = -1e-19
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ a0 = 10.55945905
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 101543.357
+ cf = 8.15e-11
+ cjd = 0.001357
+ cit = -0.0019532508
+ cjs = 0.001357
+ clc = 1e-7
+ ef = 1.0
+ k1 = 0.274
+ cle = 0.6
+ k2 = 0.039127322
+ k3 = -1.8419
+ em = 1000000.0
+ bvd = 8.7
+ bvs = 8.7
+ ll = 0
+ lw = 0
+ dlc = 3.26497e-9
+ u0 = 0.0080463574
+ w0 = 0
+ k3b = 1.9326
+ ua = -1.7148580999999998e-9
+ ub = 1.250859149999999e-18
+ uc = 5.4381728e-10
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ dwb = 0
+ ww = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ xw = 6e-9
+ wkvth0we = 2e-12
+ tnoia = 0
+ toxref = 3e-9
+ peta0 = -4.1184253e-15
+ la0 = -4.65319969e-7
+ trnqsmod = 0
+ petab = -7.719916e-16
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.0014882648800000002
+ kt1 = 0.12069622
+ lk2 = -4.2131932e-9
+ kt2 = -0.11741295
+ wketa = 1.87190595e-7
+ llc = 0
+ lln = 1
+ lu0 = 1.1331622e-10
+ mjd = 0.26
+ lua = 1.6761980000000137e-18
+ mjs = 0.26
+ lub = 8.339062399999967e-27
+ luc = -2.98810456e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ tpbsw = 0.0019
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 9.065128000000001e-14
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ nsd = 1e+20
+ pbd = 0.52
+ pat = -2.7208428e-10
+ pbs = 0.52
+ pk2 = 5.9540883e-16
+ cjswd = 8.2e-11
+ cjsws = 8.2e-11
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ pu0 = -7.954093e-17
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ prt = 0
+ pua = -1.6092489999999997e-23
+ pub = 1.5276544400000003e-32
+ puc = 5.518326299999999e-24
+ pud = 0
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = -1.1935669e-9
+ ub1 = 2.1692222300000005e-18
+ uc1 = 1.0139469700000001e-9
+ tpb = 0.0014
+ k2we = 5e-5
+ wa0 = -2.59429679e-6
+ tvfbsdoff = 0.022
+ ute = -1
+ wat = 0.0028451685
+ dsub = 0.75
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -1.1593839e-8
+ ltvoff = -1.1952424e-10
+ dtox = 2.7e-10
+ wlc = 0
+ wln = 1
+ rgatemod = 0
+ wu0 = 1.2231027e-9
+ xgl = -1.09e-8
+ xgw = 0
+ wua = 3.2583921000000013e-16
+ wub = -3.447615700000002e-25
+ wuc = -8.750290400000002e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ tnjtsswg = 1
+ )

.model nch_tt_33 nmos (
+ level = 54
+ rbodymod = 0
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ version = 4.5
+ pbswgd = 0.95
+ pbswgs = 0.95
+ ntox = 1
+ pcit = 0
+ pclm = 1.8851852
+ tempmod = 0
+ igcmod = 1
+ phin = 0.15
+ aigbacc = 0.02
+ pkt1 = 0
+ wpdiblc2 = -2.9834e-10
+ pvoff = 0
+ cdscb = 0
+ cdscd = 0
+ pvsat = 0
+ aigbinv = 0.0163
+ rbdb = 50
+ prwb = 0
+ prwg = 0
+ pub1 = 0
+ wk2we = 5e-12
+ pvth0 = 0
+ drout = 0.56
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ rdsw = 100
+ permod = 1
+ voffl = 0
+ weta0 = 0
+ wkvth0we = 2e-12
+ cgidl = 0.22
+ trnqsmod = 0
+ voffcv = -0.16942
+ wpemod = 1
+ poxedge = 1
+ rshg = 15.6
+ binunit = 2
+ pbswd = 0.8
+ pbsws = 0.8
+ rgatemod = 0
+ tnjtsswg = 1
+ tnom = 25
+ pdits = 0
+ ags = 0.68882593
+ cigsd = 0.069865
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ tpbswg = 0.0009
+ cjd = 0.001357
+ dvt0w = 0
+ cit = 0.002342713
+ dvt1w = 0
+ cjs = 0.001357
+ clc = 1e-7
+ cle = 0.6
+ dvt2w = 0
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 9.8024918e-9
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ jtsswgd = 2.3e-7
+ pk2we = -1e-19
+ jtsswgs = 2.3e-7
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ la0 = 0
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = 0
+ kt1 = -0.21767878
+ kt2 = -0.055117852
+ ptvoff = 0
+ llc = 0
+ lln = 1
+ lu0 = 0
+ wags = 1.6994444e-8
+ mjd = 0.26
+ mjs = 0.26
+ lub = 0
+ lud = 0
+ lwc = 0
+ waigsd = 3.1789128e-12
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 0
+ tnoia = 0
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 0
+ wcit = -2.5566928e-10
+ pbs = 0.52
+ pu0 = 0
+ prt = 0
+ pub = 0
+ pud = 0
+ peta0 = 0
+ diomod = 1
+ voff = -0.095952978
+ acde = 0.4
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 9.5347726e-10
+ wketa = -1.1490089e-9
+ ub1 = -5.3850981e-19
+ uc1 = -6.0041111e-11
+ tpb = 0.0014
+ tpbsw = 0.0019
+ pditsd = 0
+ pditsl = 0
+ vsat = 84306.193
+ wa0 = 0
+ cjswgd = 2.82e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.82e-10
+ wint = 0
+ ute = -1
+ wat = 0
+ vth0 = 0.31269411
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 3.0219344e-9
+ cjswd = 8.2e-11
+ cjsws = 8.2e-11
+ wlc = 0
+ wln = 1
+ wu0 = 2.3306667e-11
+ wkt1 = -8.9145825e-10
+ wkt2 = 1.0235511e-10
+ xgl = -1.09e-8
+ mjswd = 0.11
+ xgw = 0
+ mjsws = 0.11
+ wua = -1.6467997e-17
+ wub = 3.619626e-26
+ wuc = -1.4955111e-18
+ wud = 0
+ agidl = 9.41e-8
+ wmax = 2.7e-7
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ aigc = 0.01181895
+ wmin = 1.08e-7
+ tvfbsdoff = 0.022
+ njtsswg = 9
+ mjswgd = 0.85
+ mjswgs = 0.85
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ wua1 = -3.1223388e-18
+ wub1 = 2.0807554e-26
+ wuc1 = 8.1864667e-18
+ tcjswg = 0.001
+ bigc = 0.001442
+ ckappad = 0.6
+ ckappas = 0.6
+ wwlc = 0
+ pdiblc1 = 0
+ pdiblc2 = 0.023869018
+ pdiblcb = -0.3
+ scref = 1e-6
+ cdsc = 0
+ ijthsfwd = 0.01
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ pigcd = 2.621
+ aigsd = 0.010772573
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ lvoff = 0
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ bigbacc = 0.002588
+ lvsat = 0
+ lvth0 = 0
+ fprout = 300
+ ijthsrev = 0.01
+ delta = 0.007595625
+ xrcrg1 = 12
+ xrcrg2 = 1
+ kvth0we = 0.00018
+ rnoia = 0
+ rnoib = 0
+ lintnoi = -1.5e-8
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ wtvoff = 2.5061202e-10
+ ngate = 8e+20
+ wtvfbsdoff = 0
+ ngcon = 1
+ wpclm = -9.7111111e-9
+ k2we = 5e-5
+ dsub = 0.75
+ dtox = 2.7e-10
+ gbmin = 1e-12
+ capmod = 2
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ ltvfbsdoff = 0
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ wku0we = 2e-11
+ mobmod = 0
+ eta0 = 0.2
+ etab = -0.2
+ pkvth0we = -1.3e-19
+ nfactor = 1
+ ptvfbsdoff = 0
+ tvoff = 0.00085486634
+ vfbsdoff = 0.02
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ paramchk = 1
+ nigbacc = 10
+ ku0we = -0.0007
+ beta0 = 13
+ leta0 = 0
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ dlcig = 2.5e-9
+ nigbinv = 10
+ bgidl = 2320000000.0
+ ijthdfwd = 0.01
+ keta = -0.021050128
+ dmcgt = 0
+ tcjsw = 0.000357
+ toxref = 3e-9
+ ijthdrev = 0.01
+ fnoimod = 1
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 0
+ eigbinv = 1.1
+ kt1l = 0
+ bigsd = 0.00125
+ lint = 6.5375218e-9
+ lkt1 = 0
+ wvoff = 2.9681533e-9
+ lmax = 2.001e-5
+ lmin = 8.9991e-6
+ ltvoff = 0
+ lpe0 = 9.2e-8
+ wvsat = 0.002322956
+ lpeb = 2.5e-7
+ wvth0 = -3.5513739e-9
+ a0 = 3.5
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 200000
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.015956401
+ k3 = -1.8419
+ em = 1000000.0
+ minv = -0.3
+ waigc = 1.7818122e-11
+ ll = 0
+ lw = 0
+ u0 = 0.012935556
+ w0 = 0
+ lub1 = 0
+ ua = -2.0911548e-9
+ ub = 2.2368542e-18
+ uc = 5.8018519e-11
+ ud = 0
+ cigbacc = 0.32875
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 6e-9
+ ndep = 1e+18
+ lkvth0we = -2e-12
+ pvfbsdoff = 0
+ lwlc = 0
+ moin = 5.1
+ lku0we = 2.5e-11
+ tnoimod = 0
+ epsrox = 3.9
+ xpart = 1
+ nigc = 3.083
+ cigbinv = 0.006
+ acnqsmod = 0
+ rdsmod = 0
+ egidl = 0.29734
+ igbmod = 1
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ )

.model nch_tt_34 nmos (
+ level = 54
+ paramchk = 1
+ wpclm = -9.7111111e-9
+ gbmin = 1e-12
+ wua1 = -1.7574281e-19
+ wub1 = 1.7597088e-26
+ wuc1 = 8.3134424e-18
+ jswgd = 1.28e-13
+ nfactor = 1
+ jswgs = 1.28e-13
+ paigsd = -3.8370159e-23
+ bigc = 0.001442
+ wwlc = 0
+ permod = 1
+ cdsc = 0
+ ijthdfwd = 0.01
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ nigbacc = 10
+ ijthdrev = 0.01
+ voffcv = -0.16942
+ wpemod = 1
+ tvoff = 0.00082419905
+ lpdiblc2 = -9.2950492e-9
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ nigbinv = 10
+ k2we = 5e-5
+ ku0we = -0.0007
+ beta0 = 13
+ dsub = 0.75
+ leta0 = 0
+ dtox = 2.7e-10
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ tpbswg = 0.0009
+ fnoimod = 1
+ lkvth0we = -2e-12
+ eigbinv = 1.1
+ dlcig = 2.5e-9
+ eta0 = 0.2
+ bgidl = 2320000000.0
+ etab = -0.2
+ acnqsmod = 0
+ ptvoff = -2.3727895e-16
+ waigsd = 3.1789171e-12
+ dmcgt = 0
+ tcjsw = 0.000357
+ rbodymod = 0
+ diomod = 1
+ cigbacc = 0.32875
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 2.82e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.82e-10
+ bigsd = 0.00125
+ tnoimod = 0
+ wvoff = 3.141381e-9
+ mjswgd = 0.85
+ mjswgs = 0.85
+ cigbinv = 0.006
+ wvsat = 0.002322956
+ wvth0 = -3.7363659e-9
+ wpdiblc2 = -6.4961636e-10
+ tcjswg = 0.001
+ waigc = 1.8291238e-11
+ pvfbsdoff = 0
+ version = 4.5
+ lketa = -2.7750915e-8
+ tempmod = 0
+ xpart = 1
+ egidl = 0.29734
+ aigbacc = 0.02
+ keta = -0.017963263
+ wkvth0we = 2e-12
+ wtvfbsdoff = 0
+ fprout = 300
+ lags = 4.3821463e-7
+ xrcrg1 = 12
+ xrcrg2 = 1
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = -9.2651055e-12
+ trnqsmod = 0
+ kt1l = 0
+ ltvfbsdoff = 0
+ aigbinv = 0.0163
+ wtvoff = 2.7700567e-10
+ lint = 6.5375218e-9
+ lkt1 = -8.8818468e-8
+ lkt2 = -1.6837724e-8
+ lmax = 8.9991e-6
+ lmin = 8.9908e-7
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ capmod = 2
+ rgatemod = 0
+ pvoff = -1.5573172e-15
+ tnjtsswg = 1
+ wku0we = 2e-11
+ minv = -0.3
+ lua1 = -7.4262143e-17
+ lub1 = -1.4158035e-25
+ luc1 = 6.2830403e-17
+ cdscb = 0
+ cdscd = 0
+ mobmod = 0
+ pvsat = 0
+ ndep = 1e+18
+ wk2we = 5e-12
+ pvth0 = 1.6630782e-15
+ ptvfbsdoff = 0
+ drout = 0.56
+ lwlc = 0
+ poxedge = 1
+ moin = 5.1
+ paigc = -4.2533129e-18
+ nigc = 3.083
+ voffl = 0
+ binunit = 2
+ weta0 = 0
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ laigsd = 3.3658034e-16
+ pags = 5.2134206e-15
+ cgidl = 0.22
+ ntox = 1
+ pcit = 7.9881874e-17
+ pclm = 1.8851852
+ phin = 0.15
+ pbswd = 0.8
+ pbsws = 0.8
+ ags = 0.64008125
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ pkt1 = -3.6416964e-16
+ pkt2 = -1.7740443e-15
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ cjd = 0.001357
+ cit = 0.0023437436
+ cjs = 0.001357
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 9.8024918e-9
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ pdits = 0
+ cigsd = 0.069865
+ rbdb = 50
+ pua1 = -2.6489898e-23
+ prwb = 0
+ prwg = 0
+ pub1 = 2.886209e-32
+ puc1 = -1.1415122e-24
+ dvt0w = 0
+ la0 = -1.6207075e-6
+ dvt1w = 0
+ dvt2w = 0
+ rbpb = 50
+ rbpd = 50
+ jsd = 6.11e-7
+ rbps = 50
+ jss = 6.11e-7
+ lat = -0.043222769
+ rbsb = 50
+ pvag = 1.2
+ kt1 = -0.20779908
+ lk2 = -1.5849432e-8
+ kt2 = -0.053244913
+ llc = 0
+ lln = 1
+ lu0 = -1.6792432e-9
+ mjd = 0.26
+ lua = -1.2813977e-16
+ mjs = 0.26
+ lub = -8.5009677e-26
+ luc = -2.2547224e-17
+ lud = 0
+ ijthsfwd = 0.01
+ lwc = 0
+ lwl = 0
+ rdsw = 100
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 3.8370159e-14
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 3.9904965e-9
+ pbs = 0.52
+ pk2 = -8.7965669e-16
+ pk2we = -1e-19
+ pu0 = -1.6281621e-30
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ prt = 0
+ pua = -3.3674591e-24
+ pub = -4.9159389e-33
+ puc = 2.3789498e-24
+ pud = 0
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 9.6173779e-10
+ ub1 = -5.2276116e-19
+ uc1 = -6.7030033e-11
+ njtsswg = 9
+ tpb = 0.0014
+ toxref = 3e-9
+ wa0 = -4.2680933e-9
+ tnoia = 0
+ ute = -1
+ wat = -0.0004438817
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 3.1197827e-9
+ wlc = 0
+ wln = 1
+ wu0 = 2.3306667e-11
+ ijthsrev = 0.01
+ xgl = -1.09e-8
+ xtsswgd = 0.18
+ xgw = 0
+ xtsswgs = 0.18
+ wua = -1.6093419e-17
+ wub = 3.6743083e-26
+ wuc = -1.7601329e-18
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ peta0 = 0
+ wketa = -1.4921751e-9
+ ckappad = 0.6
+ ckappas = 0.6
+ rshg = 15.6
+ pdiblc1 = 0
+ pdiblc2 = 0.02490295
+ tpbsw = 0.0019
+ pdiblcb = -0.3
+ cjswd = 8.2e-11
+ cjsws = 8.2e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ tvfbsdoff = 0.022
+ ltvoff = 2.7569894e-10
+ ppdiblc2 = 3.1579745e-15
+ bigbacc = 0.002588
+ tnom = 25
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ kvth0we = 0.00018
+ lku0we = 2.5e-11
+ epsrox = 3.9
+ scref = 1e-6
+ lintnoi = -1.5e-8
+ pigcd = 2.621
+ bigbinv = 0.004953
+ aigsd = 0.010772573
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ rdsmod = 0
+ wvfbsdoff = 0
+ igbmod = 1
+ lvoff = -1.4738881e-8
+ lvfbsdoff = 0
+ pkvth0we = -1.3e-19
+ wags = 1.6414531e-8
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ lvsat = 0
+ wcit = -2.6455491e-10
+ lvth0 = 5.661542e-8
+ pbswgd = 0.95
+ pbswgs = 0.95
+ voff = -0.094313503
+ delta = 0.007595625
+ laigc = -1.6452737e-10
+ acde = 0.4
+ a0 = 3.6802789
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ vfbsdoff = 0.02
+ igcmod = 1
+ at = 204807.87
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.017719408
+ k3 = -1.8419
+ em = 1000000.0
+ rnoia = 0
+ rnoib = 0
+ ll = 0
+ lw = 0
+ vsat = 84306.193
+ u0 = 0.013122346
+ w0 = 0
+ wint = 0
+ ua = -2.0769012e-9
+ ub = 2.2463102e-18
+ uc = 6.0526552e-11
+ ud = 0
+ vth0 = 0.30639651
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 6e-9
+ wkt1 = -8.5094995e-10
+ wkt2 = 2.996904e-10
+ wmax = 2.7e-7
+ aigc = 0.011837251
+ wmin = 1.08e-7
+ pketa = 3.0850638e-15
+ ngate = 8e+20
+ ngcon = 1
+ )

.model nch_tt_35 nmos (
+ level = 54
+ a0 = 2.7573663
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ voffl = 0
+ at = 225908.74
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.010686581
+ k3 = -1.8419
+ em = 1000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.01271229
+ w0 = 0
+ ua = -2.2251639e-9
+ ub = 2.3450974e-18
+ uc = 3.6825844e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 6e-9
+ weta0 = 0
+ keta = -0.063873893
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ voffcv = -0.16942
+ wpemod = 1
+ lags = -4.2829945e-7
+ ijthsrev = 0.01
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ cgidl = 0.22
+ lcit = -6.1890204e-10
+ kt1l = 0
+ ags = 1.6136926
+ cjd = 0.001357
+ cit = 0.0030287289
+ cjs = 0.001357
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 9.8024918e-9
+ k3b = 1.9326
+ lint = 6.5375218e-9
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ lkt1 = 4.9051427e-8
+ lkt2 = -1.4519819e-8
+ pbswd = 0.8
+ pbsws = 0.8
+ lmax = 8.9908e-7
+ lmin = 4.4908e-7
+ lpe0 = 9.2e-8
+ la0 = -7.9931523e-7
+ lpeb = 2.5e-7
+ jsd = 6.11e-7
+ ppdiblc2 = -1.3141262e-15
+ jss = 6.11e-7
+ lat = -0.062002545
+ kt1 = -0.36270908
+ lk2 = -9.5902228e-9
+ kt2 = -0.0558493
+ llc = 0
+ lln = 1
+ lu0 = -1.3142934e-9
+ njtsswg = 9
+ mjd = 0.26
+ lua = 3.8140531e-18
+ mjs = 0.26
+ lub = -1.7293024e-25
+ luc = -1.4535934e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ tpbswg = 0.0009
+ njd = 1.02
+ minv = -0.3
+ njs = 1.02
+ pa0 = -6.7606598e-14
+ lua1 = -1.6437259e-16
+ lub1 = 2.2818043e-26
+ nsd = 1e+20
+ pdits = 0
+ luc1 = 5.6450349e-17
+ pbd = 0.52
+ pat = 1.7032657e-9
+ pbs = 0.52
+ pk2 = -2.3173279e-16
+ cigsd = 0.069865
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ pu0 = 8.9578742e-18
+ prt = 0
+ ndep = 1e+18
+ pua = -1.9061799e-24
+ pub = 1.3958464e-33
+ puc = -1.352132e-24
+ pud = 0
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ lwlc = 0
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 1.0629855e-9
+ ckappad = 0.6
+ ub1 = -7.0747845e-19
+ moin = 5.1
+ uc1 = -5.9861432e-11
+ ckappas = 0.6
+ tpb = 0.0014
+ pdiblc1 = 0
+ pdiblc2 = 0.01020022
+ pdiblcb = -0.3
+ wa0 = 1.1480691e-7
+ ute = -1
+ nigc = 3.083
+ wat = 0.0021260405
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 2.3917793e-9
+ wlc = 0
+ pk2we = -1e-19
+ ptvoff = -4.8469984e-16
+ wln = 1
+ wu0 = 1.324164e-11
+ xgl = -1.09e-8
+ dvtp0 = 4e-7
+ xgw = 0
+ dvtp1 = 0.01
+ wua = -1.7735306e-17
+ wub = 2.9651178e-26
+ wuc = 2.4320938e-18
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ waigsd = 3.178874e-12
+ pkvth0we = -1.3e-19
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ tnoia = 0
+ diomod = 1
+ bigbacc = 0.002588
+ peta0 = 0
+ pags = -9.2425378e-15
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 2.82e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.82e-10
+ wketa = 5.5022601e-9
+ vfbsdoff = 0.02
+ ntox = 1
+ pcit = 1.588079e-16
+ pclm = 1.8851852
+ tpbsw = 0.0019
+ kvth0we = 0.00018
+ cjswd = 8.2e-11
+ cjsws = 8.2e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ phin = 0.15
+ tvfbsdoff = 0.022
+ lintnoi = -1.5e-8
+ bigbinv = 0.004953
+ mjswgd = 0.85
+ mjswgs = 0.85
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ paramchk = 1
+ pkt1 = -1.3211355e-14
+ pkt2 = 1.7857928e-15
+ tcjswg = 0.001
+ wtvfbsdoff = 0
+ rbdb = 50
+ pua1 = 3.1539092e-23
+ prwb = 0
+ prwg = 0
+ pub1 = -3.1533886e-32
+ puc1 = -7.798421e-24
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ scref = 1e-6
+ ijthdfwd = 0.01
+ rdsw = 100
+ pigcd = 2.621
+ aigsd = 0.010772573
+ ltvfbsdoff = 0
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ lvoff = -2.8456354e-8
+ fprout = 300
+ lvsat = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ lvth0 = 1.8754806e-8
+ ijthdrev = 0.01
+ delta = 0.007595625
+ nfactor = 1
+ laigc = -6.1235169e-11
+ lpdiblc2 = 3.7903799e-9
+ rshg = 15.6
+ rnoia = 0
+ rnoib = 0
+ wtvoff = 5.5500668e-10
+ ptvfbsdoff = 0
+ pketa = -3.1399835e-15
+ ngate = 8e+20
+ ngcon = 1
+ wpclm = -9.7111111e-9
+ capmod = 2
+ wku0we = 2e-11
+ gbmin = 1e-12
+ nigbacc = 10
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ mobmod = 0
+ tnom = 25
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ lkvth0we = -2e-12
+ nigbinv = 10
+ acnqsmod = 0
+ wags = 3.2657181e-8
+ rbodymod = 0
+ wcit = -3.5323584e-10
+ voff = -0.078900611
+ tvoff = -3.4914836e-5
+ acde = 0.4
+ fnoimod = 1
+ xjbvd = 1
+ xjbvs = 1
+ vsat = 84306.193
+ lk2we = -1.5e-12
+ eigbinv = 1.1
+ wint = 0
+ vth0 = 0.34893652
+ wkt1 = 1.358409e-8
+ wkt2 = -3.7001265e-9
+ wmax = 2.7e-7
+ aigc = 0.011721192
+ wmin = 1.08e-7
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ ku0we = -0.0007
+ beta0 = 13
+ leta0 = 0
+ wpdiblc2 = 4.3752159e-9
+ wua1 = -6.5376855e-17
+ wub1 = 8.5457734e-26
+ wuc1 = 1.5793115e-17
+ bigc = 0.001442
+ wwlc = 0
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ cigbacc = 0.32875
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ tnoimod = 0
+ cigc = 0.000625
+ toxref = 3e-9
+ dmcgt = 0
+ tcjsw = 0.000357
+ wkvth0we = 2e-12
+ cigbinv = 0.006
+ trnqsmod = 0
+ bigsd = 0.00125
+ version = 4.5
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ tempmod = 0
+ ltvoff = 1.0403103e-9
+ wvoff = -2.1121636e-9
+ k2we = 5e-5
+ wvsat = 0.002322956
+ aigbacc = 0.02
+ dsub = 0.75
+ wvth0 = -2.014741e-10
+ dtox = 2.7e-10
+ rgatemod = 0
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ tnjtsswg = 1
+ waigc = 1.00872e-11
+ pvfbsdoff = 0
+ lku0we = 2.5e-11
+ epsrox = 3.9
+ eta0 = 0.2
+ etab = -0.2
+ lketa = 1.3109546e-8
+ aigbinv = 0.0163
+ xpart = 1
+ rdsmod = 0
+ igbmod = 1
+ egidl = 0.29734
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ pbswgd = 0.95
+ pbswgs = 0.95
+ igcmod = 1
+ poxedge = 1
+ binunit = 2
+ pvoff = 3.1183375e-15
+ cdscb = 0
+ cdscd = 0
+ pvsat = 0
+ wk2we = 5e-12
+ pvth0 = -1.4829756e-15
+ drout = 0.56
+ permod = 1
+ paigc = 3.0482801e-18
+ ijthsfwd = 0.01
+ )

.model nch_tt_36 nmos (
+ level = 54
+ rshg = 15.6
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ cigbacc = 0.32875
+ tnoimod = 0
+ ku0we = -0.0007
+ a0 = 2.8517872
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ beta0 = 13
+ at = 72186.119
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.0041801551
+ k3 = -1.8419
+ em = 1000000.0
+ leta0 = 0
+ rgatemod = 0
+ ll = -1.18e-13
+ lw = 0
+ u0 = 0.010928434
+ tpbswg = 0.0009
+ w0 = 0
+ ua = -2.2247872e-9
+ ub = 2.0937783e-18
+ uc = 7.1203963e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ tnjtsswg = 1
+ ww = 0
+ xw = 6e-9
+ cigbinv = 0.006
+ tnom = 25
+ ppclm = 2.75592e-14
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ ptvoff = 2.8225911e-16
+ version = 4.5
+ waigsd = 3.178874e-12
+ tempmod = 0
+ dmcgt = 0
+ tcjsw = 0.000357
+ diomod = 1
+ wags = 2.460818e-7
+ aigbacc = 0.02
+ wcit = 1.8683634e-10
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 2.82e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.82e-10
+ voff = -0.13810998
+ acde = 0.4
+ bigsd = 0.00125
+ vsat = 84306.193
+ wint = 0
+ vth0 = 0.41155442
+ wtvfbsdoff = 0
+ wkt1 = -3.8570623e-8
+ wkt2 = -4.3121065e-11
+ aigbinv = 0.0163
+ wmax = 2.7e-7
+ mjswgd = 0.85
+ mjswgs = 0.85
+ aigc = 0.011581706
+ wmin = 1.08e-7
+ wvoff = 7.1640927e-9
+ tcjswg = 0.001
+ wvsat = 0.002322956
+ ltvfbsdoff = 0
+ wvth0 = -5.9496131e-9
+ wua1 = 2.3276683e-17
+ wub1 = 1.5603072e-26
+ wuc1 = -5.1034561e-18
+ waigc = 2.6093343e-11
+ pvfbsdoff = 0
+ bigc = 0.001442
+ wwlc = 0
+ lketa = -3.8407777e-8
+ ijthsfwd = 0.01
+ cdsc = 0
+ xpart = 1
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ poxedge = 1
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ egidl = 0.29734
+ fprout = 300
+ ptvfbsdoff = 0
+ binunit = 2
+ xrcrg1 = 12
+ xrcrg2 = 1
+ ijthsrev = 0.01
+ wtvoff = -1.1880818e-9
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ capmod = 2
+ k2we = 5e-5
+ wku0we = 2e-11
+ ppdiblc2 = 3.3310302e-16
+ dsub = 0.75
+ dtox = 2.7e-10
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ pvoff = -9.6321526e-16
+ mobmod = 0
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ cdscb = 0
+ cdscd = 0
+ pvsat = 0
+ wk2we = 5e-12
+ pvth0 = 1.0462056e-15
+ drout = 0.56
+ eta0 = 0.2
+ etab = -0.2
+ paigc = -3.9944226e-18
+ voffl = 0
+ weta0 = 0
+ pkvth0we = -1.3e-19
+ ags = -2.5747885
+ lpclm = -2.4174737e-7
+ cjd = 0.001357
+ cit = 0.00083484714
+ cjs = 0.001357
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 1.30529375e-8
+ k3b = 1.9326
+ njtsswg = 9
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ cgidl = 0.22
+ vfbsdoff = 0.02
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ la0 = -8.4086042e-7
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = 0.0056354098
+ kt1 = -0.088256509
+ lk2 = -6.7273888e-9
+ kt2 = -0.075738087
+ ckappad = 0.6
+ ckappas = 0.6
+ llc = -1.18e-13
+ lln = 0.7
+ lu0 = -5.2939671e-10
+ mjd = 0.26
+ pdiblc1 = 0
+ pdiblc2 = 0.031716534
+ lua = 3.6483177e-18
+ mjs = 0.26
+ lub = -6.2349821e-26
+ luc = -1.6579966e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ pdiblcb = -0.3
+ njd = 1.02
+ njs = 1.02
+ pa0 = 8.661463e-14
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ pbswd = 0.8
+ pbsws = 0.8
+ nsd = 1e+20
+ pbd = 0.52
+ pat = -3.1418679e-9
+ pbs = 0.52
+ pk2 = -2.2869691e-16
+ paramchk = 1
+ pu0 = 2.4409578e-18
+ prt = 0
+ pua = -4.9144669e-25
+ pub = 1.8790045e-33
+ puc = 1.8346553e-24
+ pud = 0
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 5.8363721e-10
+ ub1 = -5.3348382e-19
+ uc1 = 8.6067289e-11
+ tpb = 0.0014
+ wa0 = -2.3569588e-7
+ ute = -1
+ wat = 0.013137708
+ pdits = 0
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 2.3848778e-9
+ wlc = 0
+ wln = 1
+ cigsd = 0.069865
+ wu0 = 2.8052813e-11
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -2.0950609e-17
+ wub = 2.8553091e-26
+ wuc = -4.8106046e-18
+ wud = 0
+ wwc = 0
+ bigbacc = 0.002588
+ wwl = 0
+ wwn = 1
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ ijthdfwd = 0.01
+ kvth0we = 0.00018
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ toxref = 3e-9
+ lintnoi = -1.5e-8
+ keta = 0.053210932
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ tnoia = 0
+ lags = 1.4146322e-6
+ ijthdrev = 0.01
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ peta0 = 0
+ lcit = 3.4640592e-10
+ wketa = -7.2433388e-9
+ kt1l = 0
+ lpdiblc2 = -5.676798e-9
+ tpbsw = 0.0019
+ cjswd = 8.2e-11
+ cjsws = 8.2e-11
+ mjswd = 0.11
+ tvfbsdoff = 0.022
+ mjsws = 0.11
+ ltvoff = -1.663256e-9
+ agidl = 9.41e-8
+ lint = 9.7879675e-9
+ lkt1 = -7.1707703e-8
+ lkt2 = -5.7687528e-9
+ lmax = 4.4908e-7
+ lmin = 2.1577e-7
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ minv = -0.3
+ lku0we = 2.5e-11
+ lua1 = 4.6540649e-17
+ lub1 = -5.3739597e-26
+ luc1 = -7.7582888e-18
+ epsrox = 3.9
+ lkvth0we = -2e-12
+ ndep = 1e+18
+ nfactor = 1
+ lwlc = 0
+ moin = 5.1
+ scref = 1e-6
+ rdsmod = 0
+ pigcd = 2.621
+ nigc = 3.083
+ igbmod = 1
+ aigsd = 0.010772573
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ acnqsmod = 0
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ lvoff = -2.4042325e-9
+ pbswgd = 0.95
+ noff = 2.7195
+ pbswgs = 0.95
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ lvsat = 0
+ rbodymod = 0
+ lvth0 = -8.7970687e-9
+ igcmod = 1
+ nigbacc = 10
+ delta = 0.007595625
+ pags = -1.0314937e-13
+ laigc = 1.3898222e-13
+ ntox = 1
+ pcit = -7.882386e-17
+ pclm = 2.434611
+ rnoia = 0
+ rnoib = 0
+ phin = 0.15
+ pketa = 2.46808e-15
+ ngate = 8e+20
+ nigbinv = 10
+ ngcon = 1
+ wpclm = -7.2345657e-8
+ pkt1 = 9.7367187e-15
+ pkt2 = 1.7671038e-16
+ wpdiblc2 = 6.3151306e-10
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ permod = 1
+ rbdb = 50
+ pua1 = -7.4684646e-24
+ prwb = 0
+ prwg = 0
+ pub1 = -7.978346e-34
+ puc1 = 1.3960704e-24
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ fnoimod = 1
+ rdsw = 100
+ eigbinv = 1.1
+ wkvth0we = 2e-12
+ voffcv = -0.16942
+ wpemod = 1
+ trnqsmod = 0
+ tvoff = 0.006109554
+ )

.model nch_tt_37 nmos (
+ level = 54
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ pdits = 0
+ cigsd = 0.069865
+ lkvth0we = -2e-12
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ eta0 = 0.2
+ etab = -0.2
+ ptvoff = -1.8615536e-17
+ waigsd = 3.178874e-12
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ acnqsmod = 0
+ diomod = 1
+ wtvfbsdoff = 0
+ tnoia = 0
+ pditsd = 0
+ pditsl = 0
+ rbodymod = 0
+ cjswgd = 2.82e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.82e-10
+ a0 = -2.4455841
+ a1 = 0
+ a2 = 1
+ peta0 = 0
+ b0 = 0
+ b1 = 0
+ ltvfbsdoff = 0
+ at = 121458.51
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = -0.005397302
+ k3 = -1.8419
+ em = 1000000.0
+ ll = -1.18e-13
+ wketa = 1.5290605e-8
+ lw = 0
+ u0 = 0.009324213
+ w0 = 0
+ ua = -2.2679307e-9
+ ub = 1.903479518e-18
+ uc = 2.5998306e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 6e-9
+ tpbsw = 0.0019
+ nfactor = 1
+ tvfbsdoff = 0.022
+ cjswd = 8.2e-11
+ cjsws = 8.2e-11
+ mjswgd = 0.85
+ mjswd = 0.11
+ mjswgs = 0.85
+ mjsws = 0.11
+ agidl = 9.41e-8
+ tcjswg = 0.001
+ wpdiblc2 = 2.0871493e-9
+ ptvfbsdoff = 0
+ nigbacc = 10
+ scref = 1e-6
+ wvfbsdoff = 0
+ pigcd = 2.621
+ lvfbsdoff = 0
+ aigsd = 0.010772573
+ fprout = 300
+ lvoff = 6.451419999999991e-11
+ nigbinv = 10
+ keta = -0.11923047
+ xrcrg1 = 12
+ xrcrg2 = 1
+ wkvth0we = 2e-12
+ lvsat = -0.0003892742950000001
+ lvth0 = -7.861937700000001e-9
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ trnqsmod = 0
+ delta = 0.007595625
+ lcit = -3.9333293e-11
+ wtvoff = 2.3786433e-10
+ laigc = -6.7426314e-12
+ kt1l = 0
+ rnoia = 0
+ rnoib = 0
+ fnoimod = 1
+ lint = 9.7879675e-9
+ pketa = -2.286582e-15
+ ngate = 8e+20
+ capmod = 2
+ eigbinv = 1.1
+ lkt1 = 5.5879381e-10
+ lkt2 = 1.6714521e-10
+ lmax = 2.1577e-7
+ ngcon = 1
+ lmin = 9e-8
+ wpclm = 1.5314007e-7
+ wku0we = 2e-11
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ mobmod = 0
+ rgatemod = 0
+ gbmin = 1e-12
+ tnjtsswg = 1
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ minv = -0.3
+ lua1 = -6.7367772e-18
+ lub1 = -3.8361216e-26
+ luc1 = -1.0970607e-17
+ ndep = 1e+18
+ lwlc = 0
+ moin = 5.1
+ nigc = 3.083
+ cigbacc = 0.32875
+ tnoimod = 0
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ cigbinv = 0.006
+ tvoff = -0.0028392003
+ ntox = 1
+ pcit = 1.4940572e-17
+ pclm = 1.0592301
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ phin = 0.15
+ version = 4.5
+ tempmod = 0
+ pkt1 = -1.8629533e-16
+ pkt2 = -2.0087744e-16
+ ku0we = -0.0007
+ beta0 = 13
+ leta0 = 0
+ ppclm = -2.0018289e-14
+ aigbacc = 0.02
+ rbdb = 50
+ pua1 = 2.2068447e-24
+ prwb = 0
+ prwg = 0
+ pub1 = -2.7426774e-33
+ puc1 = 1.8773731e-24
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ ijthsfwd = 0.01
+ rdsw = 100
+ toxref = 3e-9
+ aigbinv = 0.0163
+ dmcgt = 0
+ tcjsw = 0.000357
+ ijthsrev = 0.01
+ rshg = 15.6
+ bigsd = 0.00125
+ ltvoff = 2.2493116e-10
+ wvoff = 1.8056166e-9
+ poxedge = 1
+ wvsat = 0.00180338308
+ ppdiblc2 = 2.596377e-17
+ wvth0 = -2.8481029999999965e-10
+ binunit = 2
+ pvfbsdoff = 0
+ lku0we = 2.5e-11
+ waigc = 5.3999849e-12
+ tnom = 25
+ epsrox = 3.9
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ rdsmod = 0
+ lketa = -2.0226409e-9
+ igbmod = 1
+ xpart = 1
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ egidl = 0.29734
+ pbswgd = 0.95
+ pbswgs = 0.95
+ pkvth0we = -1.3e-19
+ wags = -2.4277778e-7
+ igcmod = 1
+ wcit = -2.5754486e-10
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ voff = -0.149810363
+ acde = 0.4
+ vfbsdoff = 0.02
+ vsat = 86151.12359999999
+ wint = 0
+ vth0 = 0.407122633
+ wkt1 = 8.4578791e-9
+ wkt2 = 1.7463947e-9
+ wmax = 2.7e-7
+ aigc = 0.01161432
+ wmin = 1.08e-7
+ paramchk = 1
+ pvoff = 1.6741822e-16
+ wua1 = -2.2577864e-17
+ wub1 = 2.4820337e-26
+ wuc1 = -7.3845115e-18
+ cdscb = 0
+ cdscd = 0
+ bigc = 0.001442
+ permod = 1
+ pvsat = 1.0963312e-10
+ wwlc = 0
+ njtsswg = 9
+ wk2we = 5e-12
+ pvth0 = -1.4906061999999999e-16
+ drout = 0.56
+ ags = 4.1296296
+ paigc = 3.7187593e-19
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ ijthdfwd = 0.01
+ cdsc = 0
+ cjd = 0.001357
+ cit = 0.0026629951
+ cgbo = 0
+ cjs = 0.001357
+ clc = 1e-7
+ cle = 0.6
+ voffl = 0
+ cgdl = 3.31989e-12
+ bvd = 8.7
+ cgdo = 4.90562e-11
+ xtid = 3
+ bvs = 8.7
+ xtis = 3
+ dlc = 1.30529375e-8
+ ckappad = 0.6
+ ckappas = 0.6
+ k3b = 1.9326
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ cigc = 0.000625
+ pdiblc1 = 0
+ pdiblc2 = 0.0095469071
+ pdiblcb = -0.3
+ weta0 = 0
+ voffcv = -0.16942
+ wpemod = 1
+ lpclm = 4.8457997e-8
+ la0 = 2.768849e-7
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.0047610641
+ kt1 = -0.43075175
+ lk2 = -4.7065454e-9
+ kt2 = -0.10387031
+ ijthdrev = 0.01
+ llc = -1.18e-13
+ lln = 0.7
+ lu0 = -1.9090617e-10
+ mjd = 0.26
+ mjs = 0.26
+ lua = 1.2751594e-17
+ lub = -2.21968369e-26
+ cgidl = 0.22
+ luc = -7.0415723e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = -2.9632335e-14
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 5.025644e-10
+ pbs = 0.52
+ pk2 = 3.1759465e-16
+ lpdiblc2 = -9.9900678e-10
+ pu0 = 4.2802262e-19
+ bigbacc = 0.002588
+ prt = 0
+ pua = 3.9870432e-24
+ pub = -6.31495433e-33
+ puc = 2.2635812e-25
+ pud = 0
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 8.3613685e-10
+ ub1 = -6.0636714e-19
+ uc1 = 1.0129155e-10
+ tpb = 0.0014
+ wa0 = 3.1523761e-7
+ kvth0we = 0.00018
+ pbswd = 0.8
+ pbsws = 0.8
+ ute = -1
+ wat = -0.0041344832
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -2.0418175e-10
+ wlc = 0
+ wln = 1
+ wu0 = 3.759279e-11
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -4.2175679e-17
+ wub = 6.73870221e-26
+ wuc = 2.8116572e-18
+ wud = 0
+ k2we = 5e-5
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ lintnoi = -1.5e-8
+ tpbswg = 0.0009
+ dsub = 0.75
+ bigbinv = 0.004953
+ dtox = 2.7e-10
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ )

.model nch_tt_38 nmos (
+ level = 54
+ dmcgt = 0
+ poxedge = 1
+ pkvth0we = -1.3e-19
+ tcjsw = 0.000357
+ pditsd = 0
+ pditsl = 0
+ noff = 2.7195
+ cjswgd = 2.82e-10
+ pku0we = -1.5e-18
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ cjswgs = 2.82e-10
+ binunit = 2
+ vfbsdoff = 0.02
+ ntox = 1
+ pcit = -1.2745239e-18
+ pclm = 2.2357699
+ bigsd = 0.00125
+ ptvfbsdoff = 0
+ mjswgd = 0.85
+ mjswgs = 0.85
+ tcjswg = 0.001
+ phin = 0.15
+ wvoff = 4.874463324000002e-9
+ paramchk = 1
+ pkt1 = -2.4505624e-15
+ pkt2 = 3.9546557e-16
+ wvsat = 0.0029164640999999984
+ wvth0 = 2.0191566000000033e-9
+ pvfbsdoff = 0
+ waigc = -1.2918923e-11
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ rbdb = 50
+ pua1 = -4.7371604e-25
+ prwb = 0
+ pub1 = 1.7893787999999998e-33
+ prwg = 0
+ puc1 = -4.218097e-24
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ lketa = 2.9224258e-8
+ a0 = 0.7744856
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ ijthdfwd = 0.01
+ at = 98374.6784
+ cf = 8.15e-11
+ xpart = 1
+ ef = 1.0
+ k1 = 0.274
+ k2 = -0.043338197
+ k3 = -1.8419
+ em = 1000000.0
+ rdsw = 100
+ ll = 0
+ lw = 0
+ u0 = 0.0051212099
+ w0 = 0
+ ua = -2.6695158e-9
+ ub = 2.0926996330000003e-18
+ uc = -9.6044814e-11
+ ud = 0
+ fprout = 300
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 6e-9
+ xrcrg1 = 12
+ xrcrg2 = 1
+ egidl = 0.29734
+ ijthdrev = 0.01
+ wtvoff = 2.7545299e-10
+ lpdiblc2 = 4.9724259e-14
+ rshg = 15.6
+ njtsswg = 9
+ capmod = 2
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ wku0we = 2e-11
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = -0.0010813536
+ mobmod = 0
+ pdiblcb = -0.3
+ ags = 4.1296296
+ pvoff = -1.2105337000000015e-16
+ cjd = 0.001357
+ cit = 0.001090691
+ cjs = 0.001357
+ clc = 1e-7
+ cle = 0.6
+ cdscb = 0
+ cdscd = 0
+ bvd = 8.7
+ tnom = 25
+ bvs = 8.7
+ dlc = 3.26497e-9
+ pvsat = 5.003500000000013e-12
+ k3b = 1.9326
+ lkvth0we = -2e-12
+ wk2we = 5e-12
+ toxe = 2.43e-9
+ dwb = 0
+ dwc = 0
+ toxm = 2.43e-9
+ dwg = 0
+ dwj = 0
+ pvth0 = -3.6563349999999995e-16
+ drout = 0.56
+ paigc = 2.0938533e-18
+ bigbacc = 0.002588
+ la0 = -2.5801646e-8
+ voffl = 0
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.0025911842499999997
+ kt1 = -0.62571779
+ kt2 = -0.068117715
+ lk2 = -1.1401013e-9
+ llc = 0
+ lln = 1
+ lu0 = 2.0417612e-10
+ mjd = 0.26
+ acnqsmod = 0
+ mjs = 0.26
+ lua = 5.0500592e-17
+ lub = -3.9983527e-26
+ luc = 4.4304811e-18
+ lud = 0
+ laigsd = 1.06572e-17
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ kvth0we = 0.00018
+ weta0 = 4.2794074e-8
+ pa0 = 2.9413877e-15
+ wetab = -1.5859302e-8
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 4.4193749e-10
+ pbs = 0.52
+ pk2 = 2.316472e-16
+ lpclm = -6.2136744e-8
+ pu0 = -4.0281775e-17
+ wags = -2.4277778e-7
+ prt = 0
+ pua = -3.0159915e-24
+ pub = 1.3943639e-33
+ puc = 2.394639e-25
+ pud = 0
+ lintnoi = -1.5e-8
+ rbodymod = 0
+ wcit = -8.5043837e-11
+ bigbinv = 0.004953
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 7.2026227e-10
+ vtsswgd = 4.2
+ ub1 = -7.393822000000001e-19
+ vtsswgs = 4.2
+ uc1 = -2.7209866e-10
+ cgidl = 0.22
+ tpb = 0.0014
+ wa0 = -3.1291358e-8
+ voff = -0.11849200800000002
+ ute = -1
+ wat = -0.00348951596
+ acde = 0.4
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 7.1015279e-10
+ wlc = 0
+ wln = 1
+ wu0 = 4.7067574e-10
+ xgl = -1.09e-8
+ xgw = 0
+ wua = 3.2324691e-17
+ wub = -1.4627000299999995e-26
+ wuc = 2.6722336e-18
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ vsat = 63376.513000000006
+ wint = 0
+ vth0 = 0.26853340800000003
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ wkt1 = 3.2545826e-8
+ wkt2 = -4.5976799e-9
+ wmax = 2.7e-7
+ aigc = 0.011905208
+ wmin = 1.08e-7
+ pbswd = 0.8
+ pbsws = 0.8
+ wpdiblc2 = 2.3634934e-9
+ wua1 = 5.9387403e-18
+ wub1 = -2.3393026e-26
+ wuc1 = 5.7460914e-17
+ pdits = 0
+ bigc = 0.001442
+ cigsd = 0.069865
+ wwlc = 0
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ cdsc = 0
+ nfactor = 1
+ toxref = 3e-9
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ wkvth0we = 2e-12
+ tnoia = 0
+ peta0 = -4.0226429e-15
+ trnqsmod = 0
+ petab = 1.4907744e-15
+ wketa = -4.815885e-9
+ tpbsw = 0.0019
+ ltvoff = 1.3417313e-10
+ nigbacc = 10
+ tvfbsdoff = 0.022
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ cjswd = 8.2e-11
+ cjsws = 8.2e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ k2we = 5e-5
+ nigbinv = 10
+ dsub = 0.75
+ rgatemod = 0
+ lku0we = 2.5e-11
+ dtox = 2.7e-10
+ tnjtsswg = 1
+ epsrox = 3.9
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ rdsmod = 0
+ eta0 = -0.13238438
+ etab = 0.18670848
+ igbmod = 1
+ scref = 1e-6
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ pigcd = 2.621
+ aigsd = 0.010772573
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ fnoimod = 1
+ pbswgd = 0.95
+ pbswgs = 0.95
+ eigbinv = 1.1
+ lvoff = -2.8794112000000013e-9
+ igcmod = 1
+ lvsat = 0.0017515391499999995
+ lvth0 = 5.1654495e-9
+ delta = 0.007595625
+ laigc = -3.4086068e-11
+ rnoia = 0
+ rnoib = 0
+ pketa = -3.9657201e-16
+ ngate = 8e+20
+ paigsd = -2.9413875e-24
+ ngcon = 1
+ cigbacc = 0.32875
+ wpclm = -8.3073835e-8
+ gbmin = 1e-12
+ tnoimod = 0
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ permod = 1
+ cigbinv = 0.006
+ ijthsfwd = 0.01
+ voffcv = -0.16942
+ wpemod = 1
+ version = 4.5
+ keta = -0.45164428
+ tempmod = 0
+ ijthsrev = 0.01
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 1.084633e-10
+ tvoff = -0.0018736893
+ aigbacc = 0.02
+ kt1l = 0
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ lint = 0
+ lkt1 = 1.8885602e-8
+ lkt2 = -3.1935983e-9
+ lmax = 9e-8
+ lmin = 5.4e-8
+ tpbswg = 0.0009
+ ku0we = -0.0007
+ aigbinv = 0.0163
+ beta0 = 13
+ lpe0 = 9.2e-8
+ ppdiblc2 = -1.2574432e-20
+ lpeb = 2.5e-7
+ leta0 = 3.1244132e-8
+ letab = -3.6350598e-8
+ wtvfbsdoff = 0
+ minv = -0.3
+ ppclm = 2.1858187e-15
+ lua1 = 4.1554342e-18
+ lub1 = -2.5857803e-26
+ luc1 = 2.4128073e-17
+ ndep = 1e+18
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ ptvoff = -2.2148869e-17
+ lwlc = 0
+ moin = 5.1
+ ltvfbsdoff = 0
+ waigsd = 3.1789053e-12
+ nigc = 3.083
+ diomod = 1
+ )

.model nch_tt_39 nmos (
+ level = 54
+ wkt1 = 5.960945e-9
+ wkt2 = 1.1625249e-8
+ wmax = 2.7e-7
+ aigc = 0.011615807
+ wmin = 1.08e-7
+ fnoimod = 1
+ eigbinv = 1.1
+ wua1 = -1.0774777e-16
+ wub1 = 1.7109629e-25
+ wuc1 = 1.606153e-17
+ bigc = 0.001442
+ wwlc = 0
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ scref = 1e-6
+ ijthsfwd = 0.01
+ cdsc = 0
+ fprout = 300
+ pigcd = 2.621
+ cgbo = 0
+ aigsd = 0.010772573
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ xrcrg1 = 12
+ xrcrg2 = 1
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ lvoff = -6.4884398999999995e-9
+ cigbacc = 0.32875
+ lvsat = -0.0022565101000000002
+ wtvoff = 7.91509e-11
+ lvth0 = 7.910732700000003e-9
+ ijthsrev = 0.01
+ tnoimod = 0
+ delta = 0.007595625
+ laigc = -1.730084e-11
+ rnoia = 0
+ rnoib = 0
+ cigbinv = 0.006
+ dmcg = 3.1e-8
+ capmod = 2
+ dmci = 3.1e-8
+ dmdg = 0
+ wku0we = 2e-11
+ pketa = 1.224516e-15
+ ngate = 8e+20
+ a0 = 19.191807
+ a1 = 0
+ a2 = 1
+ ngcon = 1
+ b0 = 0
+ b1 = 0
+ mobmod = 0
+ wpclm = -5.2664346e-8
+ at = 103079.96199999998
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = -0.057713829
+ k3 = -1.8419
+ em = 1000000.0
+ k2we = 5e-5
+ ll = 0
+ lw = 0
+ u0 = 0.0021507365
+ w0 = 0
+ ua = -2.3710013e-9
+ ub = 1.4550579529999998e-18
+ uc = -1.4785261e-10
+ ud = 0
+ version = 4.5
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 6e-9
+ dsub = 0.75
+ dtox = 2.7e-10
+ gbmin = 1e-12
+ tempmod = 0
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ eta0 = 1.1504337
+ aigbacc = 0.02
+ etab = -1.3364008
+ pkvth0we = -1.3e-19
+ aigbinv = 0.0163
+ tvoff = -0.0045522389
+ vfbsdoff = 0.02
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ paramchk = 1
+ ku0we = -0.0007
+ beta0 = 13
+ leta0 = -4.3159315e-8
+ poxedge = 1
+ letab = 5.198974e-8
+ ppclm = 4.2206835e-16
+ binunit = 2
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ ijthdfwd = 0.01
+ toxref = 3e-9
+ dmcgt = 0
+ keta = 0.16119603
+ tcjsw = 0.000357
+ ijthdrev = 0.01
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 4.6179023e-10
+ ltvoff = 2.8952901e-10
+ kt1l = 0
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ bigsd = 0.00125
+ lint = 0
+ wvoff = -2.2288246e-9
+ lkt1 = 1.0413925e-8
+ lkt2 = 8.1983323e-9
+ lmax = 5.4e-8
+ lmin = 4.5e-8
+ wvsat = -0.0033283578000000017
+ lku0we = 2.5e-11
+ pvfbsdoff = 0
+ lpe0 = 9.2e-8
+ wvth0 = -3.1224421e-9
+ lpeb = 2.5e-7
+ epsrox = 3.9
+ waigc = 4.0939876e-11
+ minv = -0.3
+ lua1 = -3.9796071e-17
+ lub1 = 5.119547099999998e-26
+ luc1 = 1.4911728e-19
+ rdsmod = 0
+ lkvth0we = -2e-12
+ ndep = 1e+18
+ igbmod = 1
+ lwlc = 0
+ lketa = -6.3204807e-9
+ moin = 5.1
+ njtsswg = 9
+ xpart = 1
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ nigc = 3.083
+ pbswgd = 0.95
+ pbswgs = 0.95
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ acnqsmod = 0
+ egidl = 0.29734
+ igcmod = 1
+ ckappad = 0.6
+ ckappas = 0.6
+ noff = 2.7195
+ pdiblc1 = 0
+ pdiblc2 = -0.0010804963
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ pdiblcb = -0.3
+ rbodymod = 0
+ ntox = 1
+ pcit = -2.1822647e-17
+ pclm = 1.0542662
+ ags = 4.1296296
+ bigbacc = 0.002588
+ phin = 0.15
+ cjd = 0.001357
+ cit = -0.0050011527
+ cjs = 0.001357
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 3.26497e-9
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ pkt1 = -9.0863924e-16
+ pkt2 = -5.454643e-16
+ dwg = 0
+ dwj = 0
+ kvth0we = 0.00018
+ wpdiblc2 = 2.3632766e-9
+ permod = 1
+ pvoff = 2.9093734999999984e-16
+ lintnoi = -1.5e-8
+ la0 = -1.0940063e-6
+ cdscb = 0
+ cdscd = 0
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.0028640905800000004
+ bigbinv = 0.004953
+ kt1 = -0.47965441
+ kt2 = -0.26453031
+ lk2 = -3.0631458e-10
+ vtsswgd = 4.2
+ pvsat = 3.6720318000000004e-10
+ vtsswgs = 4.2
+ llc = 0
+ lln = 1
+ lu0 = 3.7646358e-10
+ wk2we = 5e-12
+ pvth0 = -6.7420746e-17
+ mjd = 0.26
+ mjs = 0.26
+ lua = 3.3186753e-17
+ lub = -3.0003129999999985e-27
+ luc = 7.435334e-18
+ lud = 0
+ rbdb = 50
+ pua1 = 6.1201017e-24
+ prwb = 0
+ lwc = 0
+ pub1 = -9.491001900000001e-33
+ prwg = 0
+ drout = 0.56
+ lwl = 0
+ puc1 = -1.8169327e-24
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 1.2471671e-13
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ nsd = 1e+20
+ pvag = 1.2
+ pbd = 0.52
+ pat = 1.5402954e-10
+ pbs = 0.52
+ pk2 = 1.8168527e-16
+ paigc = -1.0299571e-18
+ pu0 = -9.9060704e-18
+ prt = 0
+ pua = 6.5377716e-24
+ pub = -1.101976303e-32
+ rdsw = 100
+ puc = -3.076481e-25
+ pud = 0
+ voffl = 0
+ rsh = 17.5
+ tcj = 0.00076
+ voffcv = -0.16942
+ wpemod = 1
+ ua1 = 1.4780468e-9
+ ub1 = -2.0678869e-18
+ uc1 = 1.4133161e-10
+ tpb = 0.0014
+ wa0 = -2.130866e-6
+ weta0 = -1.5669611e-7
+ ute = -1
+ wetab = 4.0317659e-8
+ wat = 0.001474414299999999
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 1.5715655e-9
+ wlc = 0
+ wln = 1
+ wu0 = -5.3043297e-11
+ lpclm = 6.3904735e-9
+ xgl = -1.09e-8
+ wkvth0we = 2e-12
+ xgw = 0
+ wua = -1.3239536e-16
+ wub = 1.9940967600000001e-25
+ wuc = 1.2105201e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ cgidl = 0.22
+ trnqsmod = 0
+ rshg = 15.6
+ wtvfbsdoff = 0
+ nfactor = 1
+ pbswd = 0.8
+ pbsws = 0.8
+ tpbswg = 0.0009
+ ltvfbsdoff = 0
+ rgatemod = 0
+ tnjtsswg = 1
+ pdits = 0
+ tnom = 25
+ cigsd = 0.069865
+ toxe = 2.43e-9
+ ptvoff = -1.0763348e-17
+ toxm = 2.43e-9
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ waigsd = 3.1788545e-12
+ nigbacc = 10
+ pk2we = -1e-19
+ diomod = 1
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ ptvfbsdoff = 0
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 2.82e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.82e-10
+ wags = -2.4277778e-7
+ tnoia = 0
+ nigbinv = 10
+ wcit = 2.6923414e-10
+ peta0 = 7.5477876e-15
+ petab = -1.7674893e-15
+ voff = -0.056267378999999965
+ wketa = -3.2765679e-8
+ acde = 0.4
+ tvfbsdoff = 0.022
+ tpbsw = 0.0019
+ mjswgd = 0.85
+ mjswgs = 0.85
+ vsat = 132480.81299999997
+ wint = 0
+ cjswd = 8.2e-11
+ cjsws = 8.2e-11
+ vth0 = 0.22120093900000004
+ tcjswg = 0.001
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ )

.model nch_tt_40 nmos (
+ level = 54
+ wkt1 = -2.6238067e-8
+ wkt2 = -1.1473225e-8
+ wmax = 2.7e-7
+ aigc = 0.011144932
+ wmin = 1.08e-7
+ fnoimod = 1
+ eigbinv = 1.1
+ wua1 = 1.9140234e-16
+ wub1 = -2.597066e-25
+ wuc1 = -2.3798265000000004e-17
+ bigc = 0.001442
+ wwlc = 0
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ scref = 1e-6
+ ijthsfwd = 0.01
+ cdsc = 0
+ fprout = 300
+ pigcd = 2.621
+ cgbo = 0
+ aigsd = 0.010772574
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ xrcrg1 = 12
+ xrcrg2 = 1
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ lvoff = -5.5742293e-9
+ cigbacc = 0.32875
+ lvsat = 0.00560742952
+ wtvoff = -7.2128996e-10
+ lvth0 = -7.795251999999998e-10
+ ijthsrev = 0.01
+ tnoimod = 0
+ delta = 0.007595625
+ laigc = 5.7720314e-12
+ rnoia = 0
+ rnoib = 0
+ cigbinv = 0.006
+ dmcg = 3.1e-8
+ capmod = 2
+ dmci = 3.1e-8
+ dmdg = 0
+ wku0we = 2e-11
+ pketa = -8.4677334e-15
+ ngate = 8e+20
+ a0 = -5.925916599999999
+ a1 = 0
+ a2 = 1
+ ngcon = 1
+ b0 = 0
+ b1 = 0
+ mobmod = 0
+ wpclm = -7.2101286e-7
+ at = 66521.242
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.015523130999999996
+ k3 = -1.8419
+ em = 1000000.0
+ k2we = 5e-5
+ ll = 0
+ lw = 0
+ u0 = 0.013709058
+ w0 = 0
+ ua = -5.589164400000002e-10
+ ub = 8.937269600000036e-20
+ uc = 2.381934e-10
+ ud = 0
+ version = 4.5
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 6e-9
+ dsub = 0.75
+ dtox = 2.7e-10
+ gbmin = 1e-12
+ tempmod = 0
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ eta0 = -0.288265897
+ aigbacc = 0.02
+ etab = -0.74723747
+ laigsd = -1.5325105e-17
+ pkvth0we = -1.3e-19
+ aigbinv = 0.0163
+ tvoff = 0.0062987975
+ vfbsdoff = 0.02
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ paramchk = 1
+ ku0we = -0.0007
+ beta0 = 13
+ leta0 = 2.7336964e-8
+ poxedge = 1
+ letab = 2.3120738e-8
+ ppclm = 3.3171145e-14
+ binunit = 2
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ ijthdfwd = 0.01
+ toxref = 3e-9
+ dmcgt = 0
+ keta = -0.51478944
+ tcjsw = 0.000357
+ ijthdrev = 0.01
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 1.370515e-10
+ ltvoff = -2.4217179e-10
+ kt1l = 0
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ bigsd = 0.00125
+ lint = 0
+ wvoff = 9.960383100000001e-9
+ lkt1 = -1.4940467e-9
+ lkt2 = -1.1864945e-9
+ lmax = 4.5e-8
+ lmin = 3.6e-8
+ wvsat = 0.0237570614
+ lku0we = 2.5e-11
+ pvfbsdoff = 0
+ lpe0 = 9.2e-8
+ wvth0 = -2.0711547e-8
+ lpeb = 2.5e-7
+ epsrox = 3.9
+ waigc = 5.1623453e-11
+ minv = -0.3
+ lua1 = 6.0050187e-18
+ lub1 = -6.8748353e-27
+ luc1 = 6.4275095e-18
+ rdsmod = 0
+ lkvth0we = -2e-12
+ ndep = 1e+18
+ igbmod = 1
+ lwlc = 0
+ lketa = 2.6802806000000003e-8
+ moin = 5.1
+ njtsswg = 9
+ xpart = 1
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ nigc = 3.083
+ pbswgd = 0.95
+ pbswgs = 0.95
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ acnqsmod = 0
+ egidl = 0.29734
+ igcmod = 1
+ ckappad = 0.6
+ ckappas = 0.6
+ noff = 2.7195
+ pdiblc1 = 0
+ pdiblc2 = -0.0010804963
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ pdiblcb = -0.3
+ rbodymod = 0
+ ntox = 1
+ pcit = 1.116072e-17
+ pclm = 4.6708343
+ ags = 4.1296296
+ bigbacc = 0.002588
+ phin = 0.15
+ paigsd = 4.2297301e-24
+ cjd = 0.001357
+ cit = 0.0016261683
+ cjs = 0.001357
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 3.26497e-9
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ pkt1 = 6.6911236e-16
+ pkt2 = 5.863609e-16
+ dwg = 0
+ dwj = 0
+ kvth0we = 0.00018
+ wpdiblc2 = 2.3632766e-9
+ permod = 1
+ pvoff = -3.0633384e-16
+ lintnoi = -1.5e-8
+ la0 = 1.3676219000000002e-7
+ cdscb = 0
+ cdscd = 0
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.00107271332
+ bigbinv = 0.004953
+ kt1 = -0.23663458
+ kt2 = -0.073003235
+ lk2 = -3.894925700000001e-9
+ vtsswgd = 4.2
+ pvsat = -9.5998236e-10
+ vtsswgs = 4.2
+ llc = 0
+ lln = 1
+ lu0 = -1.8989416e-10
+ wk2we = 5e-12
+ pvth0 = 7.9444539e-16
+ mjd = 0.26
+ mjs = 0.26
+ lua = -5.56054081e-17
+ lub = 6.391826569999999e-26
+ luc = -1.14809219e-17
+ lud = 0
+ rbdb = 50
+ pua1 = -8.5382538e-24
+ prwb = 0
+ lwc = 0
+ pub1 = 1.1618339e-32
+ prwg = 0
+ drout = 0.56
+ lwl = 0
+ puc1 = 1.361972e-25
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = -7.5523402e-14
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ nsd = 1e+20
+ pvag = 1.2
+ pbd = 0.52
+ pat = -3.8677652e-10
+ pbs = 0.52
+ pk2 = 5.0756697e-16
+ paigc = -1.5534524e-18
+ pu0 = 4.1451338e-18
+ prt = 0
+ pua = -2.8276596999999977e-25
+ pub = -6.331388000000253e-35
+ rdsw = 100
+ puc = 4.398917e-25
+ pud = 0
+ voffl = 0
+ rsh = 17.5
+ tcj = 0.00076
+ voffcv = -0.16942
+ wpemod = 1
+ ua1 = 5.4333072e-10
+ ub1 = -8.8277854e-19
+ uc1 = 1.3201149999999995e-11
+ tpb = 0.0014
+ wa0 = 1.9556670799999998e-6
+ weta0 = 9.4960797e-8
+ ute = -1
+ wetab = 3.9258957e-9
+ wat = 0.0125112725
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -5.0790816e-9
+ wlc = 0
+ wln = 1
+ wu0 = -3.3980257e-10
+ lpclm = -1.70821362e-7
+ xgl = -1.09e-8
+ wkvth0we = 2e-12
+ xgw = 0
+ wua = 6.799270000000015e-18
+ wub = -2.4191335000000008e-26
+ wuc = -3.150715e-18
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ cgidl = 0.22
+ trnqsmod = 0
+ rshg = 15.6
+ wtvfbsdoff = 0
+ nfactor = 1
+ pbswd = 0.8
+ pbsws = 0.8
+ tpbswg = 0.0009
+ ltvfbsdoff = 0
+ rgatemod = 0
+ tnjtsswg = 1
+ pdits = 0
+ tnom = 25
+ cigsd = 0.069865
+ toxe = 2.43e-9
+ ptvoff = 2.8458255e-17
+ toxm = 2.43e-9
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ waigsd = 3.1787682e-12
+ nigbacc = 10
+ pk2we = -1e-19
+ diomod = 1
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ ptvfbsdoff = 0
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 2.82e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.82e-10
+ wags = -2.4277778e-7
+ tnoia = 0
+ nigbinv = 10
+ wcit = -4.0389578e-10
+ peta0 = -4.7834008e-15
+ petab = 1.5707054e-17
+ voff = -0.074924736
+ wketa = 1.65035329e-7
+ acde = 0.4
+ tvfbsdoff = 0.022
+ tpbsw = 0.0019
+ mjswgd = 0.85
+ mjswgs = 0.85
+ vsat = -28007.757999999987
+ wint = 0
+ cjswd = 8.2e-11
+ cjsws = 8.2e-11
+ vth0 = 0.398553147
+ tcjswg = 0.001
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ )

.model nch_ff_1 nmos (
+ level = 54
+ fprout = 300
+ xrcrg1 = 12
+ xrcrg2 = 1
+ ags = 0.7975000000000001
+ wtvoff = 0
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ tvoff = 0.0019109629
+ keta = -0.06
+ cjd = 0.0012620099999999998
+ cit = 0.0001
+ cjs = 0.0012620099999999998
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 9.8024918e-9
+ xjbvd = 1
+ k3b = 1.9326
+ xjbvs = 1
+ lk2we = -1.5e-12
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ tvfbsdoff = 0.022
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = -1e-11
+ capmod = 2
+ la0 = 0
+ kt1l = 0
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.0001
+ kt1 = -0.200226
+ kt2 = -0.05325
+ wku0we = 2e-11
+ wkvth0we = 2e-12
+ llc = 0
+ ku0we = -0.0007
+ lln = 1
+ lu0 = 6e-12
+ mjd = 0.26
+ mjs = 0.26
+ beta0 = 13
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ leta0 = 0
+ njs = 1.02
+ pa0 = 0
+ mobmod = 0
+ nsd = 1e+20
+ pbd = 0.52
+ pat = -2.8e-11
+ pbs = 0.52
+ lint = 6.5375218e-9
+ trnqsmod = 0
+ pu0 = 2e-18
+ prt = 0
+ pud = 0
+ lkt1 = -1.1e-9
+ lmax = 2.001e-5
+ lmin = 9.00077e-6
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 1.2299687e-9
+ ub1 = -7.2455506e-19
+ uc1 = 3.028e-11
+ dlcig = 2.5e-9
+ tpb = 0.0014
+ lpe0 = 9.2e-8
+ njtsswg = 9
+ bgidl = 2320000000.0
+ lpeb = 2.5e-7
+ wa0 = 0
+ ute = -1.007
+ wat = 0
+ web = 6843.8
+ wec = -25529.0
+ wlc = 0
+ wln = 1
+ wu0 = -3.6e-11
+ xgl = -1.09e-8
+ xgw = 0
+ wud = 0
+ wwc = 0
+ minv = -0.3
+ wwl = 0
+ wwn = 1
+ xtsswgd = 0.18
+ wvfbsdoff = 0
+ xtsswgs = 0.18
+ lvfbsdoff = 0
+ lub1 = 0
+ ndep = 1e+18
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.018555248
+ lwlc = 0
+ rgatemod = 0
+ dmcgt = 0
+ pdiblcb = -0.3
+ moin = 5.1
+ tcjsw = 0.000357
+ tnjtsswg = 1
+ nigc = 3.083
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ bigsd = 0.00125
+ bigbacc = 0.002588
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ wvoff = 0
+ ntox = 2.029
+ pcit = -1.5e-17
+ kvth0we = 0.00018
+ pclm = 1.4
+ wvsat = 0
+ wvth0 = -4e-9
+ lintnoi = -1.5e-8
+ bigbinv = 0.004953
+ phin = 0.15
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ pkt1 = -5e-17
+ a0 = 3.25
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 72000
+ cf = 8.720500000000001e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.022601254
+ k3 = -1.8419
+ em = 1000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.01527
+ w0 = 0
+ ua = -1.8237726e-9
+ ub = 2.103696e-18
+ xpart = 1
+ uc = 7.33e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 2.33e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ toxref = 3e-9
+ rbdb = 50
+ prwb = 0
+ prwg = 0
+ pub1 = 0
+ egidl = 0.29734
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ rdsw = 100
+ ijthsfwd = 0.01
+ ltvoff = 0
+ nfactor = 1
+ rshg = 15.6
+ ijthsrev = 0.01
+ pvoff = 0
+ lku0we = 2.5e-11
+ cdscb = 0
+ cdscd = 0
+ epsrox = 3.9
+ pvsat = -1.8e-11
+ wk2we = 5e-12
+ pvth0 = -2.3e-16
+ drout = 0.56
+ nigbacc = 10
+ rdsmod = 0
+ igbmod = 1
+ voffl = 0
+ tnom = 25
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ toxe = 2.3900000000000002e-9
+ toxm = 2.43e-9
+ weta0 = 0
+ pbswgd = 0.95
+ pbswgs = 0.95
+ nigbinv = 10
+ igcmod = 1
+ cgidl = 0.22
+ wags = -1.5e-8
+ wcit = 5e-11
+ voff = -0.1128204
+ fnoimod = 1
+ pbswd = 0.8
+ pbsws = 0.8
+ acde = 0.4
+ pkvth0we = -1.3e-19
+ eigbinv = 1.1
+ vsat = 102860
+ wint = 0
+ vth0 = 0.32111089
+ wkt1 = -2e-9
+ pvfbsdoff = 0
+ wmax = 0.00090001
+ aigc = 0.011769394
+ wmin = 8.9974e-6
+ pdits = 0
+ vfbsdoff = 0.02
+ permod = 1
+ cigsd = 0.069865
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ bigc = 0.001442
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ paramchk = 1
+ wwlc = 0
+ cigbacc = 0.32875
+ voffcv = -0.16942
+ wpemod = 1
+ cdsc = 0
+ tnoia = 0
+ tnoimod = 0
+ cgbo = 0
+ cgdl = 3.5522823e-12
+ cgdo = 5.2490134000000004e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.5522823e-12
+ cgso = 5.2490134000000004e-11
+ cigc = 0.000625
+ peta0 = 0
+ cigbinv = 0.006
+ tpbsw = 0.0019
+ ijthdfwd = 0.01
+ cjswd = 7.625999999999999e-11
+ cjsws = 7.625999999999999e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ version = 4.5
+ tempmod = 0
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ tpbswg = 0.0009
+ ijthdrev = 0.01
+ aigbacc = 0.02
+ k2we = 5e-5
+ dsub = 0.75
+ dtox = 2.7e-10
+ scref = 1e-6
+ ptvoff = 0
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ pigcd = 2.621
+ aigsd = 0.01077322
+ lvoff = -2e-11
+ eta0 = 0.3
+ aigbinv = 0.0163
+ diomod = 1
+ etab = -0.25
+ wtvfbsdoff = 0
+ lvsat = -0.0003
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 2.6226e-10
+ pku0we = -1.5e-18
+ lvth0 = -1e-10
+ cjswgs = 2.6226e-10
+ lkvth0we = -2e-12
+ delta = 0.007595625
+ ltvfbsdoff = 0
+ rnoia = 0
+ rnoib = 0
+ mjswgd = 0.85
+ mjswgs = 0.85
+ acnqsmod = 0
+ ngate = 8e+20
+ tcjswg = 0.001
+ ngcon = 1
+ poxedge = 1
+ rbodymod = 0
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ binunit = 2
+ ptvfbsdoff = 0
+ )

.model nch_ff_2 nmos (
+ level = 54
+ wtvoff = 0
+ cgidl = 0.22
+ ijthdfwd = 0.01
+ capmod = 2
+ pbswd = 0.8
+ pbsws = 0.8
+ wku0we = 2e-11
+ rshg = 15.6
+ cigbacc = 0.32875
+ mobmod = 0
+ pvfbsdoff = 0
+ ijthdrev = 0.01
+ tnoimod = 0
+ pdits = 0
+ lpdiblc2 = -5.8501673e-10
+ cigsd = 0.069865
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ cigbinv = 0.006
+ tnom = 25
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ toxe = 2.3900000000000002e-9
+ toxm = 2.43e-9
+ version = 4.5
+ tnoia = 0
+ tempmod = 0
+ lkvth0we = -2e-12
+ peta0 = 0
+ tpbsw = 0.0019
+ aigbacc = 0.02
+ wags = -1.5e-8
+ cjswd = 7.625999999999999e-11
+ cjsws = 7.625999999999999e-11
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ wcit = 5e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ acnqsmod = 0
+ voff = -0.11120139
+ acde = 0.4
+ vsat = 102860
+ wint = 0
+ rbodymod = 0
+ aigbinv = 0.0163
+ vth0 = 0.31536703
+ wkt1 = -2e-9
+ wmax = 0.00090001
+ aigc = 0.01178613
+ wmin = 8.9974e-6
+ scref = 1e-6
+ pigcd = 2.621
+ toxref = 3e-9
+ aigsd = 0.01077322
+ bigc = 0.001442
+ wwlc = 0
+ lvoff = -1.4574874e-8
+ poxedge = 1
+ cdsc = 0
+ lvsat = -0.0003
+ cgbo = 0
+ cgdl = 3.5522823e-12
+ cgdo = 5.2490134000000004e-11
+ xtid = 3
+ xtis = 3
+ lvth0 = 5.1537332e-8
+ cgsl = 3.5522823e-12
+ cgso = 5.2490134000000004e-11
+ cigc = 0.000625
+ delta = 0.007595625
+ binunit = 2
+ laigc = -1.5044982e-10
+ rnoia = 0
+ rnoib = 0
+ ltvoff = -1.4627394e-10
+ a0 = 3.4752469
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ ngate = 8e+20
+ at = 61592.494
+ cf = 8.720500000000001e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.024088843
+ k3 = -1.8419
+ em = 1000000.0
+ ngcon = 1
+ ll = 0
+ lw = 0
+ u0 = 0.015491951000000002
+ w0 = 0
+ ua = -1.7995884e-9
+ ub = 2.1046515e-18
+ uc = 7.3387901e-11
+ ud = 0
+ wkvth0we = 2e-12
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 2.33e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ lku0we = 2.5e-11
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ trnqsmod = 0
+ epsrox = 3.9
+ k2we = 5e-5
+ rdsmod = 0
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ dsub = 0.75
+ dtox = 2.7e-10
+ igbmod = 1
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ ags = 0.8010490100000001
+ pbswgd = 0.95
+ pbswgs = 0.95
+ eta0 = 0.3
+ cjd = 0.0012620099999999998
+ rgatemod = 0
+ etab = -0.25
+ cit = -2.3830864e-5
+ cjs = 0.0012620099999999998
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 9.8024918e-9
+ tnjtsswg = 1
+ k3b = 1.9326
+ igcmod = 1
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ tvoff = 0.0019272336
+ la0 = -2.0249698e-6
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = 0.093463481
+ kt1 = -0.19577666
+ lk2 = -1.337342e-8
+ kt2 = -0.051823539
+ xjbvd = 1
+ llc = 0
+ xjbvs = 1
+ lln = 1
+ tvfbsdoff = 0.022
+ lk2we = -1.5e-12
+ lu0 = -1.9893360999999997e-9
+ mjd = 0.26
+ lua = -2.1741579e-16
+ mjs = 0.26
+ lub = -8.5898229e-27
+ luc = -7.902321e-19
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njtsswg = 9
+ njd = 1.02
+ njs = 1.02
+ pa0 = 0
+ nsd = 1e+20
+ pbd = 0.52
+ pat = -2.8e-11
+ pbs = 0.52
+ pu0 = 2e-18
+ xtsswgd = 0.18
+ prt = 0
+ pud = 0
+ xtsswgs = 0.18
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 1.2713861e-9
+ ub1 = -7.4616446e-19
+ ku0we = -0.0007
+ uc1 = 2.5703642e-11
+ ckappad = 0.6
+ ckappas = 0.6
+ beta0 = 13
+ tpb = 0.0014
+ wa0 = 0
+ leta0 = 0
+ pdiblc1 = 0
+ pdiblc2 = 0.018620322
+ pdiblcb = -0.3
+ ute = -1.0077691
+ wat = 0
+ web = 6843.8
+ wec = -25529.0
+ wlc = 0
+ wln = 1
+ wu0 = -3.6e-11
+ xgl = -1.09e-8
+ xgw = 0
+ permod = 1
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ bigbacc = 0.002588
+ voffcv = -0.16942
+ wpemod = 1
+ dmcgt = 0
+ tcjsw = 0.000357
+ kvth0we = 0.00018
+ lintnoi = -1.5e-8
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ keta = -0.059896633
+ ijthsfwd = 0.01
+ bigsd = 0.00125
+ lags = -3.1905621e-8
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 1.1032395e-9
+ wvoff = 0
+ kt1l = 0
+ tpbswg = 0.0009
+ wvsat = 0
+ wvth0 = -4e-9
+ ijthsrev = 0.01
+ lint = 6.5375218e-9
+ lkt1 = -4.1099573000000004e-8
+ lkt2 = -1.2823887e-8
+ wtvfbsdoff = 0
+ lmax = 9.00077e-6
+ lmin = 9.0075e-7
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ ptvoff = 0
+ lketa = -9.2926692e-10
+ xpart = 1
+ ltvfbsdoff = 0
+ minv = -0.3
+ lua1 = -3.7234224e-16
+ lub1 = 1.9426851e-25
+ luc1 = 4.1141459e-17
+ nfactor = 1
+ diomod = 1
+ ndep = 1e+18
+ lute = 6.9145309e-9
+ egidl = 0.29734
+ lwlc = 0
+ moin = 5.1
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 2.6226e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.6226e-10
+ nigc = 3.083
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ mjswgd = 0.85
+ mjswgs = 0.85
+ nigbacc = 10
+ ptvfbsdoff = 0
+ tcjswg = 0.001
+ ntox = 2.029
+ pkvth0we = -1.3e-19
+ pcit = -1.5e-17
+ pclm = 1.4
+ pvoff = 0
+ nigbinv = 10
+ phin = 0.15
+ cdscb = 0
+ cdscd = 0
+ vfbsdoff = 0.02
+ pvsat = -1.8e-11
+ wk2we = 5e-12
+ pkt1 = -5e-17
+ pvth0 = -2.3e-16
+ drout = 0.56
+ voffl = 0
+ fprout = 300
+ paramchk = 1
+ rbdb = 50
+ prwb = 0
+ prwg = 0
+ pub1 = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ fnoimod = 1
+ weta0 = 0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ eigbinv = 1.1
+ rdsw = 100
+ )

.model nch_ff_3 nmos (
+ level = 54
+ ku0we = -0.0007
+ beta0 = 13
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ leta0 = 0
+ ijthsrev = 0.01
+ kvth0we = 0.00018
+ lintnoi = -1.5e-8
+ k2we = 5e-5
+ bigbinv = 0.004953
+ dlcig = 2.5e-9
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ bgidl = 2320000000.0
+ dsub = 0.75
+ wvfbsdoff = 0
+ dtox = 2.7e-10
+ lvfbsdoff = 0
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ eta0 = 0.3
+ dmcgt = 0
+ etab = -0.25
+ tcjsw = 0.000357
+ bigsd = 0.00125
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ wvoff = 0
+ pkvth0we = -1.3e-19
+ nfactor = 1
+ wvsat = 0
+ wvth0 = -4e-9
+ vfbsdoff = 0.02
+ lketa = -2.6515603e-8
+ toxref = 3e-9
+ xpart = 1
+ nigbacc = 10
+ paramchk = 1
+ egidl = 0.29734
+ nigbinv = 10
+ keta = -0.031147941
+ ltvoff = -6.4393769e-10
+ ijthdfwd = 0.01
+ lags = 4.0889306e-7
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = -1.2051822e-10
+ kt1l = 0
+ lku0we = 2.5e-11
+ fnoimod = 1
+ ijthdrev = 0.01
+ epsrox = 3.9
+ eigbinv = 1.1
+ pvoff = 0
+ lint = 6.5375218e-9
+ cdscb = 0
+ cdscd = 0
+ lkt1 = -1.8864368e-8
+ lkt2 = -1.1493547e-8
+ lmax = 9.0075e-7
+ lpdiblc2 = 3.0380287e-9
+ pvsat = -1.8e-11
+ lmin = 4.5075e-7
+ rdsmod = 0
+ wk2we = 5e-12
+ pvth0 = -2.3e-16
+ drout = 0.56
+ igbmod = 1
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ minv = -0.3
+ voffl = 0
+ lua1 = -1.0281867e-16
+ lub1 = 1.8552992e-26
+ luc1 = 3.7680622e-18
+ pbswgd = 0.95
+ pbswgs = 0.95
+ ndep = 1e+18
+ weta0 = 0
+ lwlc = 0
+ igcmod = 1
+ moin = 5.1
+ a0 = 1.288
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ cigbacc = 0.32875
+ at = 219598.22
+ cf = 8.720500000000001e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.023010322
+ k3 = -1.8419
+ em = 1000000.0
+ ll = 0
+ nigc = 3.083
+ lw = 0
+ u0 = 0.014990444
+ w0 = 0
+ ua = -1.9429424e-9
+ ub = 2.1566e-18
+ uc = 9.3717778e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 2.33e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ lkvth0we = -2e-12
+ cgidl = 0.22
+ tnoimod = 0
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ cigbinv = 0.006
+ acnqsmod = 0
+ pbswd = 0.8
+ pbsws = 0.8
+ ntox = 2.029
+ pcit = -1.5e-17
+ pclm = 1.4
+ pvfbsdoff = 0
+ rbodymod = 0
+ version = 4.5
+ permod = 1
+ phin = 0.15
+ tempmod = 0
+ pdits = 0
+ cigsd = 0.069865
+ pkt1 = -5e-17
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ aigbacc = 0.02
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ voffcv = -0.16942
+ wpemod = 1
+ rbdb = 50
+ prwb = 0
+ pub1 = 0
+ prwg = 0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ tnoia = 0
+ rdsw = 100
+ aigbinv = 0.0163
+ peta0 = 0
+ tpbsw = 0.0019
+ wtvfbsdoff = 0
+ cjswd = 7.625999999999999e-11
+ cjsws = 7.625999999999999e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ tpbswg = 0.0009
+ rshg = 15.6
+ ltvfbsdoff = 0
+ wkvth0we = 2e-12
+ poxedge = 1
+ trnqsmod = 0
+ ptvoff = 0
+ binunit = 2
+ scref = 1e-6
+ pigcd = 2.621
+ aigsd = 0.01077322
+ tnom = 25
+ diomod = 1
+ toxe = 2.3900000000000002e-9
+ toxm = 2.43e-9
+ ptvfbsdoff = 0
+ lvoff = -1.3788912e-8
+ pditsd = 0
+ rgatemod = 0
+ pditsl = 0
+ cjswgd = 2.6226e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.6226e-10
+ tnjtsswg = 1
+ lvsat = -0.0003
+ lvth0 = 7.3115504e-9
+ delta = 0.007595625
+ laigc = -5.5724245e-11
+ rnoia = 0
+ rnoib = 0
+ mjswgd = 0.85
+ mjswgs = 0.85
+ wags = -1.5e-8
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ wcit = 5e-11
+ tcjswg = 0.001
+ ngate = 8e+20
+ voff = -0.1120845
+ acde = 0.4
+ ngcon = 1
+ vsat = 102860
+ wint = 0
+ vth0 = 0.36505891999999995
+ gbmin = 1e-12
+ wkt1 = -2e-9
+ jswgd = 1.28e-13
+ wmax = 0.00090001
+ jswgs = 1.28e-13
+ aigc = 0.011679696
+ wmin = 8.9974e-6
+ ags = 0.3057696
+ cjd = 0.0012620099999999998
+ cit = 0.0013511778
+ cjs = 0.0012620099999999998
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 9.8024918e-9
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ fprout = 300
+ dwg = 0
+ dwj = 0
+ njtsswg = 9
+ bigc = 0.001442
+ xrcrg1 = 12
+ xrcrg2 = 1
+ wwlc = 0
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ la0 = -7.832e-8
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.047161618
+ kt1 = -0.22076004
+ kt2 = -0.053318302
+ lk2 = -1.2413537e-8
+ llc = 0
+ cdsc = 0
+ lln = 1
+ lu0 = -1.5429956e-9
+ ckappad = 0.6
+ ckappas = 0.6
+ mjd = 0.26
+ mjs = 0.26
+ lua = -8.9830708e-17
+ lub = -5.4824e-26
+ luc = -1.8883822e-17
+ lud = 0
+ lwc = 0
+ cgbo = 0
+ wtvoff = 0
+ lwl = 0
+ lwn = 1
+ cgdl = 3.5522823e-12
+ cgdo = 5.2490134000000004e-11
+ xtid = 3
+ pdiblc1 = 0
+ pdiblc2 = 0.014549485
+ njd = 1.02
+ xtis = 3
+ njs = 1.02
+ pa0 = 0
+ pdiblcb = -0.3
+ nsd = 1e+20
+ pbd = 0.52
+ pat = -2.8e-11
+ pbs = 0.52
+ cgsl = 3.5522823e-12
+ cgso = 5.2490134000000004e-11
+ cigc = 0.000625
+ pu0 = 2e-18
+ tvoff = 0.0024864064
+ prt = 0
+ pud = 0
+ tvfbsdoff = 0.022
+ rsh = 17.5
+ tcj = 0.00076
+ ijthsfwd = 0.01
+ xjbvd = 1
+ ua1 = 9.685506e-10
+ ub1 = -5.4873129e-19
+ xjbvs = 1
+ uc1 = 6.7696222e-11
+ lk2we = -1.5e-12
+ tpb = 0.0014
+ capmod = 2
+ wa0 = 0
+ ute = -1
+ wat = 0
+ web = 6843.8
+ wec = -25529.0
+ wlc = 0
+ wln = 1
+ wku0we = 2e-11
+ wu0 = -3.6e-11
+ xgl = -1.09e-8
+ xgw = 0
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ bigbacc = 0.002588
+ mobmod = 0
+ )

.model nch_ff_4 nmos (
+ level = 54
+ minv = -0.3
+ lua1 = -3.0475764e-17
+ pk2we = -1e-19
+ lub1 = -2.9971927e-26
+ luc1 = -4.3987511e-18
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ ndep = 1e+18
+ rgatemod = 0
+ lwlc = 0
+ moin = 5.1
+ tnjtsswg = 1
+ tnoia = 0
+ nigc = 3.083
+ peta0 = 0
+ poxedge = 1
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ tpbsw = 0.0019
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ binunit = 2
+ cjswd = 7.625999999999999e-11
+ cjsws = 7.625999999999999e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ ntox = 2.029
+ pcit = -1.5e-17
+ pclm = 1.5439223
+ phin = 0.15
+ pkt1 = -5e-17
+ toxref = 3e-9
+ scref = 1e-6
+ jtsswgd = 2.3e-7
+ pigcd = 2.621
+ jtsswgs = 2.3e-7
+ aigsd = 0.01077322
+ rbdb = 50
+ prwb = 0
+ pub1 = 0
+ prwg = 0
+ lvoff = -6.341613400000001e-9
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ rdsw = 100
+ lvsat = -0.0003
+ lvth0 = -4.790878e-9
+ delta = 0.007595625
+ ltvoff = -1.206053e-10
+ laigc = -1.9935708e-11
+ rnoia = 0
+ rnoib = 0
+ ijthsfwd = 0.01
+ ngate = 8e+20
+ njtsswg = 9
+ ngcon = 1
+ rshg = 15.6
+ lku0we = 2.5e-11
+ ags = -0.015684402000000007
+ epsrox = 3.9
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ cjd = 0.0012620099999999998
+ cit = 0.00073144105
+ ijthsrev = 0.01
+ cjs = 0.0012620099999999998
+ clc = 1e-7
+ cle = 0.6
+ gbmin = 1e-12
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 1.30529375e-8
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ k3b = 1.9326
+ ckappad = 0.6
+ ckappas = 0.6
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ rdsmod = 0
+ pdiblc1 = 0
+ pdiblc2 = 0.027331777
+ pdiblcb = -0.3
+ igbmod = 1
+ la0 = -2.4730306e-7
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.016965258
+ kt1 = -0.23920434
+ kt2 = -0.070668297
+ lk2 = -9.6174482e-9
+ llc = -1.18e-13
+ lln = 0.7
+ lu0 = -6.1833887e-10
+ mjd = 0.26
+ mjs = 0.26
+ lua = -1.0757894e-17
+ lub = -4.7838952e-26
+ luc = -6.6488035e-18
+ lud = 0
+ pbswgd = 0.95
+ pbswgs = 0.95
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ tnom = 25
+ njd = 1.02
+ njs = 1.02
+ pa0 = 0
+ nsd = 1e+20
+ pbd = 0.52
+ pat = -2.8e-11
+ pbs = 0.52
+ toxe = 2.3900000000000002e-9
+ toxm = 2.43e-9
+ pu0 = 2e-18
+ igcmod = 1
+ prt = 0
+ pud = 0
+ bigbacc = 0.002588
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 8.041349e-10
+ ub1 = -4.3844738e-19
+ uc1 = 8.6257162e-11
+ tpb = 0.0014
+ wa0 = 0
+ ute = -1
+ wat = 0
+ web = 6843.8
+ wec = -25529.0
+ kvth0we = 0.00018
+ wlc = 0
+ wln = 1
+ wu0 = -3.6e-11
+ xgl = -1.09e-8
+ xgw = 0
+ tvoff = 0.0012970146
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ tvfbsdoff = 0.022
+ lintnoi = -1.5e-8
+ xjbvd = 1
+ xjbvs = 1
+ wags = -1.5e-8
+ lk2we = -1.5e-12
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ wcit = 5e-11
+ voff = -0.12901018
+ acde = 0.4
+ pkvth0we = -1.3e-19
+ ku0we = -0.0007
+ beta0 = 13
+ vsat = 102860
+ wint = 0
+ permod = 1
+ leta0 = 0
+ vth0 = 0.39256442999999996
+ wkt1 = -2e-9
+ wmax = 0.00090001
+ aigc = 0.011598359
+ wmin = 8.9974e-6
+ vfbsdoff = 0.02
+ a0 = 1.6720524
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 150970.13
+ cf = 8.720500000000001e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.016655575
+ k3 = -1.8419
+ em = 1000000.0
+ dlcig = 2.5e-9
+ ll = -1.18e-13
+ wvfbsdoff = 0
+ lw = 0
+ u0 = 0.012888952
+ bgidl = 2320000000.0
+ w0 = 0
+ lvfbsdoff = 0
+ ua = -2.1226533e-9
+ ub = 2.1407249e-18
+ uc = 6.5910917e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 2.33e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ voffcv = -0.16942
+ wpemod = 1
+ bigc = 0.001442
+ paramchk = 1
+ wwlc = 0
+ wtvfbsdoff = 0
+ dmcgt = 0
+ tcjsw = 0.000357
+ nfactor = 1
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.5522823e-12
+ cgdo = 5.2490134000000004e-11
+ xtid = 3
+ xtis = 3
+ ltvfbsdoff = 0
+ cgsl = 3.5522823e-12
+ cgso = 5.2490134000000004e-11
+ cigc = 0.000625
+ ijthdfwd = 0.01
+ bigsd = 0.00125
+ tpbswg = 0.0009
+ wvoff = 0
+ nigbacc = 10
+ wvsat = 0
+ wvth0 = -4e-9
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ ijthdrev = 0.01
+ ptvfbsdoff = 0
+ lpdiblc2 = -2.58618e-9
+ ptvoff = 0
+ nigbinv = 10
+ k2we = 5e-5
+ dsub = 0.75
+ lketa = -2.2644187e-8
+ dtox = 2.7e-10
+ xpart = 1
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ diomod = 1
+ pditsd = 0
+ pditsl = 0
+ egidl = 0.29734
+ cjswgd = 2.6226e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.6226e-10
+ eta0 = 0.3
+ etab = -0.25
+ fnoimod = 1
+ eigbinv = 1.1
+ lkvth0we = -2e-12
+ mjswgd = 0.85
+ mjswgs = 0.85
+ tcjswg = 0.001
+ acnqsmod = 0
+ rbodymod = 0
+ pvoff = 0
+ cigbacc = 0.32875
+ cdscb = 0
+ cdscd = 0
+ pvsat = -1.8e-11
+ wk2we = 5e-12
+ pvth0 = -2.3e-16
+ drout = 0.56
+ tnoimod = 0
+ fprout = 300
+ voffl = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ cigbinv = 0.006
+ weta0 = 0
+ lpclm = -6.3325799e-8
+ wtvoff = 0
+ version = 4.5
+ cgidl = 0.22
+ tempmod = 0
+ keta = -0.039946614
+ capmod = 2
+ lags = 5.5033282e-7
+ wku0we = 2e-11
+ aigbacc = 0.02
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 1.5216594e-10
+ pbswd = 0.8
+ mobmod = 0
+ pbsws = 0.8
+ kt1l = 0
+ wkvth0we = 2e-12
+ pvfbsdoff = 0
+ lint = 9.7879675e-9
+ trnqsmod = 0
+ pdits = 0
+ lkt1 = -1.07488734e-8
+ lkt2 = -3.8595493e-9
+ aigbinv = 0.0163
+ lmax = 4.5075e-7
+ cigsd = 0.069865
+ lmin = 2.1744e-7
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ laigsd = -8.1082969e-17
+ )

.model nch_ff_5 nmos (
+ level = 54
+ nigbinv = 10
+ bigsd = 0.00125
+ wags = -1.5e-8
+ wcit = 5e-11
+ acnqsmod = 0
+ wvoff = 0
+ voff = -0.15746310460000001
+ acde = 0.4
+ wvsat = 0
+ vsat = 102521.2852
+ wvth0 = -4e-9
+ rbodymod = 0
+ wint = 0
+ vth0 = 0.4085613742
+ wkt1 = -2e-9
+ wmax = 0.00090001
+ aigc = 0.011526753
+ wmin = 8.9974e-6
+ fnoimod = 1
+ eigbinv = 1.1
+ toxref = 3e-9
+ lketa = -1.1430034e-8
+ xpart = 1
+ bigc = 0.001442
+ wwlc = 0
+ egidl = 0.29734
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.5522823e-12
+ cgdo = 5.2490134000000004e-11
+ xtid = 3
+ xtis = 3
+ ltvoff = 1.4850105e-11
+ cgsl = 3.5522823e-12
+ cgso = 5.2490134000000004e-11
+ cigc = 0.000625
+ cigbacc = 0.32875
+ tnoimod = 0
+ lku0we = 2.5e-11
+ cigbinv = 0.006
+ epsrox = 3.9
+ wkvth0we = 2e-12
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ pvoff = 0
+ rdsmod = 0
+ trnqsmod = 0
+ cdscb = 0
+ cdscd = 0
+ igbmod = 1
+ pvsat = -1.8e-11
+ version = 4.5
+ wk2we = 5e-12
+ pvth0 = -2.3e-16
+ k2we = 5e-5
+ drout = 0.56
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ tempmod = 0
+ dsub = 0.75
+ dtox = 2.7e-10
+ pbswgd = 0.95
+ pbswgs = 0.95
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ voffl = 0
+ igcmod = 1
+ aigbacc = 0.02
+ weta0 = 0
+ eta0 = 0.3
+ rgatemod = 0
+ etab = -0.25
+ lpclm = -2.4377173e-8
+ tnjtsswg = 1
+ cgidl = 0.22
+ aigbinv = 0.0163
+ pbswd = 0.8
+ pbsws = 0.8
+ pvfbsdoff = 0
+ permod = 1
+ wtvfbsdoff = 0
+ pdits = 0
+ cigsd = 0.069865
+ dvt0w = 0
+ dvt1w = 0
+ poxedge = 1
+ dvt2w = 0
+ ltvfbsdoff = 0
+ voffcv = -0.16942
+ wpemod = 1
+ binunit = 2
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ tnoia = 0
+ peta0 = 0
+ wketa = 0
+ keta = -0.093093889
+ ptvfbsdoff = 0
+ tpbsw = 0.0019
+ ijthsfwd = 0.01
+ cjswd = 7.625999999999999e-11
+ cjsws = 7.625999999999999e-11
+ a0 = 0.66068814
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ mjswd = 0.11
+ lags = 3.3904274e-13
+ mjsws = 0.11
+ agidl = 9.41e-8
+ tpbswg = 0.0009
+ at = 79499.116
+ cf = 8.720500000000001e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = -0.018112077999999997
+ k3 = -1.8419
+ em = 1000000.0
+ jswd = 1.28e-13
+ ll = -1.18e-13
+ jsws = 1.28e-13
+ lw = 0
+ u0 = 0.010886872
+ w0 = 0
+ lcit = 7.4591162e-11
+ ua = -2.2893587e-9
+ ub = 2.089788886e-18
+ uc = 4.5969231e-11
+ ud = 0
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 2.33e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ kt1l = 0
+ ijthsrev = 0.01
+ lint = 9.7879675e-9
+ ptvoff = 0
+ lkt1 = -4.4075226000000005e-9
+ lkt2 = -6.0180086e-10
+ lmax = 2.1744e-7
+ lmin = 9.167e-8
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ scref = 1e-6
+ diomod = 1
+ pigcd = 2.621
+ minv = -0.3
+ aigsd = 0.01077322
+ lua1 = 7.6861327e-18
+ lub1 = -5.2342256e-26
+ luc1 = -4.2210821e-18
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 2.6226e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.6226e-10
+ ndep = 1e+18
+ lvoff = -3.3806259999999997e-10
+ njtsswg = 9
+ lwlc = 0
+ moin = 5.1
+ lvsat = -0.0002285156999999999
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ lvth0 = -8.1662159e-9
+ nigc = 3.083
+ delta = 0.007595625
+ mjswgd = 0.85
+ mjswgs = 0.85
+ laigc = -4.8268328e-12
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.02163037
+ pdiblcb = -0.3
+ tcjswg = 0.001
+ rnoia = 0
+ rnoib = 0
+ ags = 2.5925264
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ cjd = 0.0012620099999999998
+ cit = 0.001099094
+ cjs = 0.0012620099999999998
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 1.30529375e-8
+ pketa = 0
+ ngate = 8e+20
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ ngcon = 1
+ pkvth0we = -1.3e-19
+ ntox = 2.029
+ pcit = -1.5e-17
+ pclm = 1.3593316
+ bigbacc = 0.002588
+ la0 = -3.3904685e-8
+ gbmin = 1e-12
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.0018848735
+ kt1 = -0.26925814
+ kt2 = -0.086107863
+ lk2 = -2.2814734e-9
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ llc = -1.18e-13
+ lln = 0.7
+ phin = 0.15
+ lu0 = -1.9589995e-10
+ mjd = 0.26
+ mjs = 0.26
+ lua = 2.4416942e-17
+ lub = -3.7091512499999996e-26
+ luc = -2.4411077e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ vfbsdoff = 0.02
+ njd = 1.02
+ njs = 1.02
+ pa0 = 0
+ nsd = 1e+20
+ kvth0we = 0.00018
+ pbd = 0.52
+ pat = -2.8e-11
+ pbs = 0.52
+ pkt1 = -5e-17
+ pu0 = 2e-18
+ prt = 0
+ fprout = 300
+ pub = 0
+ pud = 0
+ lintnoi = -1.5e-8
+ rsh = 17.5
+ xrcrg1 = 12
+ xrcrg2 = 1
+ tcj = 0.00076
+ ua1 = 6.2327283e-10
+ ub1 = -3.3242687e-19
+ uc1 = 8.5415128e-11
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ tpb = 0.0014
+ wa0 = 0
+ ute = -1
+ paramchk = 1
+ wat = 0
+ web = 6843.8
+ wec = -25529.0
+ wlc = 0
+ wln = 1
+ wu0 = -3.6e-11
+ rbdb = 50
+ xgl = -1.09e-8
+ prwb = 0
+ pub1 = 0
+ prwg = 0
+ xgw = 0
+ wub = 0
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ rbpb = 50
+ rbpd = 50
+ wtvoff = 0
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ rdsw = 100
+ tvfbsdoff = 0.022
+ tvoff = 0.00065504585
+ capmod = 2
+ ijthdfwd = 0.01
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ wku0we = 2e-11
+ mobmod = 0
+ rshg = 15.6
+ ku0we = -0.0007
+ beta0 = 13
+ leta0 = 0
+ ijthdrev = 0.01
+ nfactor = 1
+ lpdiblc2 = -1.3831831e-9
+ wvfbsdoff = 0
+ dlcig = 2.5e-9
+ lvfbsdoff = 0
+ bgidl = 2320000000.0
+ laigsd = 3.3904273e-17
+ tnom = 25
+ toxe = 2.3900000000000002e-9
+ toxm = 2.43e-9
+ nigbacc = 10
+ dmcgt = 0
+ tcjsw = 0.000357
+ lkvth0we = -2e-12
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ )

.model nch_ff_6 nmos (
+ level = 54
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ vfbsdoff = 0.02
+ toxref = 3e-9
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.0069155858
+ scref = 1e-6
+ pdiblcb = -0.3
+ pigcd = 2.621
+ aigsd = 0.01077322
+ paramchk = 1
+ lvoff = -2.0844108900000003e-9
+ ags = 2.59253
+ lvsat = 0.00114527187
+ ltvoff = 1.0839662e-10
+ lvth0 = 2.7550711699999997e-9
+ bigbacc = 0.002588
+ cjd = 0.0012620099999999998
+ cit = 0.00080194411
+ cjs = 0.0012620099999999998
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ delta = 0.007595625
+ dlc = 3.26497e-9
+ k3b = 1.9326
+ laigc = -2.2427226e-11
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ keta = -0.52835722
+ rnoia = 0
+ rnoib = 0
+ ijthdfwd = 0.01
+ kvth0we = 0.00018
+ la0 = 3.0288889e-8
+ jsd = 6.11e-7
+ lintnoi = -1.5e-8
+ jss = 6.11e-7
+ lat = -0.00048029214
+ kt1 = -0.40872879
+ kt2 = -0.10088778
+ lk2 = -4.8654938e-10
+ lku0we = 2.5e-11
+ pketa = 0
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ ngate = 8e+20
+ bigbinv = 0.004953
+ llc = 0
+ lln = 1
+ lu0 = 1.1337411000000001e-10
+ lcit = 1.0252326e-10
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ mjd = 0.26
+ mjs = 0.26
+ lua = 3.5218789e-17
+ lub = -1.9869262700000004e-26
+ luc = 2.2716666e-18
+ lud = 0
+ epsrox = 3.9
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ ngcon = 1
+ njd = 1.02
+ njs = 1.02
+ kt1l = 0
+ pa0 = 0
+ nsd = 1e+20
+ pbd = 0.52
+ pat = -2.8e-11
+ pbs = 0.52
+ pu0 = 2e-18
+ prt = 0
+ pub = 0
+ puc = 0
+ pud = 0
+ rdsmod = 0
+ ijthdrev = 0.01
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ rsh = 17.5
+ jswgs = 1.28e-13
+ lint = 0
+ tcj = 0.00076
+ igbmod = 1
+ ua1 = 8.897383e-10
+ ub1 = -8.0235504e-19
+ uc1 = -6.3390556e-11
+ tpb = 0.0014
+ lkt1 = 8.7027184e-9
+ lkt2 = 7.8751111e-10
+ wa0 = 0
+ lpdiblc2 = 6.6256944e-15
+ lmax = 9.167e-8
+ ute = -1
+ wat = 0
+ web = 6843.8
+ pscbe1 = 1000000000.0
+ wec = -25529.0
+ pscbe2 = 1e-20
+ lmin = 5.567e-8
+ wlc = 0
+ wln = 1
+ wu0 = -3.6e-11
+ xgl = -1.09e-8
+ xgw = 0
+ wub = 0
+ wuc = 0
+ wud = 0
+ lpe0 = 9.2e-8
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ pbswgd = 0.95
+ lpeb = 2.5e-7
+ pbswgs = 0.95
+ minv = -0.3
+ igcmod = 1
+ lua1 = -1.7361621e-17
+ lub1 = -8.1690078e-27
+ luc1 = 9.7666522e-18
+ ndep = 1e+18
+ lwlc = 0
+ moin = 5.1
+ nigc = 3.083
+ tvfbsdoff = 0.022
+ nfactor = 1
+ lkvth0we = -2e-12
+ tvoff = -0.00034012981
+ wtvfbsdoff = 0
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ acnqsmod = 0
+ ltvfbsdoff = 0
+ permod = 1
+ ntox = 2.029
+ pcit = -1.5e-17
+ ku0we = -0.0007
+ pclm = 1.2209944
+ beta0 = 13
+ rbodymod = 0
+ leta0 = 3.0288889e-9
+ nigbacc = 10
+ letab = -2.2684433e-8
+ phin = 0.15
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ pkt1 = -5e-17
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ voffcv = -0.16942
+ wpemod = 1
+ nigbinv = 10
+ ptvfbsdoff = 0
+ rbdb = 50
+ prwb = 0
+ pub1 = 0
+ prwg = 0
+ dmcgt = 0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ tcjsw = 0.000357
+ rdsw = 100
+ fnoimod = 1
+ eigbinv = 1.1
+ bigsd = 0.00125
+ tpbswg = 0.0009
+ wvoff = 0
+ rshg = 15.6
+ wkvth0we = 2e-12
+ wvsat = 0.0
+ wvth0 = -4e-9
+ ptvoff = 0
+ trnqsmod = 0
+ cigbacc = 0.32875
+ diomod = 1
+ lketa = 2.9484719e-8
+ xpart = 1
+ pditsd = 0
+ pditsl = 0
+ tnoimod = 0
+ cjswgd = 2.6226e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.6226e-10
+ tnom = 25
+ toxe = 2.3900000000000002e-9
+ toxm = 2.43e-9
+ egidl = 0.29734
+ a0 = -0.02222221999999996
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ rgatemod = 0
+ at = 64556.761
+ cf = 8.720500000000001e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = -0.037207015
+ k3 = -1.8419
+ em = 1000000.0
+ cigbinv = 0.006
+ ll = 0
+ lw = 0
+ u0 = 0.0075967223
+ tnjtsswg = 1
+ w0 = 0
+ ua = -2.404272e-9
+ ub = 1.906573466e-18
+ uc = -4.166667e-12
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 2.33e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ mjswgd = 0.85
+ mjswgs = 0.85
+ tcjswg = 0.001
+ version = 4.5
+ wags = -1.5e-8
+ tempmod = 0
+ wcit = 5e-11
+ voff = -0.138884931
+ acde = 0.4
+ aigbacc = 0.02
+ vsat = 87906.53
+ wint = 0
+ vth0 = 0.29237747599999997
+ pvoff = 0
+ wkt1 = -2e-9
+ wmax = 0.00090001
+ aigc = 0.011713991
+ wmin = 8.9974e-6
+ cdscb = 0
+ cdscd = 0
+ pvsat = -1.8e-11
+ wk2we = 5e-12
+ pvth0 = -2.3e-16
+ fprout = 300
+ drout = 0.56
+ xrcrg1 = 12
+ xrcrg2 = 1
+ aigbinv = 0.0163
+ voffl = 0
+ bigc = 0.001442
+ wwlc = 0
+ wtvoff = 0
+ weta0 = 0
+ lpclm = -1.1373478e-8
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.5522823e-12
+ cgdo = 5.2490134000000004e-11
+ xtid = 3
+ xtis = 3
+ cgidl = 0.22
+ cgsl = 3.5522823e-12
+ cgso = 5.2490134000000004e-11
+ cigc = 0.000625
+ capmod = 2
+ wku0we = 2e-11
+ ijthsfwd = 0.01
+ poxedge = 1
+ mobmod = 0
+ pbswd = 0.8
+ pvfbsdoff = 0
+ pbsws = 0.8
+ binunit = 2
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ ijthsrev = 0.01
+ pdits = 0
+ cigsd = 0.069865
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ k2we = 5e-5
+ dsub = 0.75
+ dtox = 2.7e-10
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ eta0 = 0.26777778
+ etab = -0.0086762422
+ tnoia = 0
+ peta0 = 0
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ wketa = 0
+ tpbsw = 0.0019
+ cjswd = 7.625999999999999e-11
+ cjsws = 7.625999999999999e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ pkvth0we = -1.3e-19
+ njtsswg = 9
+ )

.model nch_ff_7 nmos (
+ level = 54
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ ltvoff = -2.4740506e-10
+ aigbacc = 0.02
+ rdsw = 100
+ ijthsfwd = 0.01
+ lku0we = 2.5e-11
+ aigbinv = 0.0163
+ epsrox = 3.9
+ rshg = 15.6
+ rdsmod = 0
+ igbmod = 1
+ ijthsrev = 0.01
+ pvoff = 0
+ cdscb = 0
+ cdscd = 0
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ pvsat = -1.8e-11
+ wk2we = 5e-12
+ pvth0 = -2.3e-16
+ drout = 0.56
+ pbswgd = 0.95
+ pbswgs = 0.95
+ igcmod = 1
+ poxedge = 1
+ wtvfbsdoff = 0
+ voffl = 0
+ tnom = 25
+ toxe = 2.3900000000000002e-9
+ toxm = 2.43e-9
+ weta0 = 0
+ binunit = 2
+ lpclm = -7.2871722e-8
+ ltvfbsdoff = 0
+ cgidl = 0.22
+ wags = -1.5e-8
+ wcit = 5e-11
+ pvfbsdoff = 0
+ permod = 1
+ pbswd = 0.8
+ pbsws = 0.8
+ voff = -0.112415764
+ pkvth0we = -1.3e-19
+ acde = 0.4
+ ptvfbsdoff = 0
+ vsat = 97937.182
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ wint = 0
+ vth0 = 0.295273177
+ wkt1 = -2e-9
+ wmax = 0.00090001
+ aigc = 0.011692671
+ pdits = 0
+ wmin = 8.9974e-6
+ vfbsdoff = 0.02
+ cigsd = 0.069865
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ voffcv = -0.16942
+ wpemod = 1
+ wub1 = 0.0
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ bigc = 0.001442
+ paramchk = 1
+ wwlc = 0
+ tnoia = 0
+ cdsc = 0
+ cgbo = 0
+ njtsswg = 9
+ cgdl = 3.5522823e-12
+ cgdo = 5.2490134000000004e-11
+ xtid = 3
+ xtis = 3
+ peta0 = 0
+ cgsl = 3.5522823e-12
+ cgso = 5.2490134000000004e-11
+ cigc = 0.000625
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ tpbsw = 0.0019
+ ijthdfwd = 0.01
+ tpbswg = 0.0009
+ ckappad = 0.6
+ cjswd = 7.625999999999999e-11
+ ckappas = 0.6
+ cjsws = 7.625999999999999e-11
+ mjswd = 0.11
+ pdiblc1 = 0
+ pdiblc2 = 0.0069157
+ mjsws = 0.11
+ agidl = 9.41e-8
+ pdiblcb = -0.3
+ ptvoff = 0
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ ijthdrev = 0.01
+ bigbacc = 0.002588
+ diomod = 1
+ k2we = 5e-5
+ dsub = 0.75
+ scref = 1e-6
+ dtox = 2.7e-10
+ pditsd = 0
+ pditsl = 0
+ kvth0we = 0.00018
+ cjswgd = 2.6226e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.6226e-10
+ ags = 2.59253
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ pigcd = 2.621
+ aigsd = 0.01077322
+ cjd = 0.0012620099999999998
+ cit = -0.0014090447
+ cjs = 0.0012620099999999998
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ lintnoi = -1.5e-8
+ dlc = 3.26497e-9
+ bigbinv = 0.004953
+ k3b = 1.9326
+ lvoff = -3.6196222000000007e-9
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ eta0 = 0.35179556
+ etab = -1.0973583
+ lvsat = 0.0005634890999999995
+ mjswgd = 0.85
+ mjswgs = 0.85
+ lvth0 = 2.5871222999999995e-9
+ la0 = -3.1577778e-7
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = 0.0065313337
+ lkvth0we = -2e-12
+ kt1 = 0.010917511
+ kt2 = -0.10990444
+ lk2 = -1.5787889e-9
+ delta = 0.007595625
+ tcjswg = 0.001
+ llc = 0
+ laigc = -2.1190647e-11
+ lln = 1
+ lu0 = 5.1187601e-10
+ mjd = 0.26
+ mjs = 0.26
+ lua = 7.8730998e-17
+ lub = -4.3148946000000005e-26
+ luc = 1.578889e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 0
+ rnoia = 0
+ rnoib = 0
+ nsd = 1e+20
+ pbd = 0.52
+ pat = -2.8e-11
+ pbs = 0.52
+ pu0 = 2e-18
+ prt = 0
+ pub = 0
+ puc = 0
+ pud = 0
+ acnqsmod = 0
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 3.744227e-10
+ ngate = 8e+20
+ ub1 = -1.2872892e-18
+ uc1 = -1.6722222e-10
+ tpb = 0.0014
+ ngcon = 1
+ wa0 = 0
+ ute = -1
+ wat = 0.0
+ web = 6843.8
+ wec = -25529.0
+ wlc = 0
+ wln = 1
+ wu0 = -3.6e-11
+ xgl = -1.09e-8
+ xgw = 0
+ wub = 0
+ wuc = 0
+ wud = 0
+ rbodymod = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ a0 = 5.9444444
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = -56333.367
+ cf = 8.720500000000001e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = -0.018375298999999998
+ k3 = -1.8419
+ em = 1000000.0
+ fprout = 300
+ ll = 0
+ lw = 0
+ u0 = 0.00072599922
+ nfactor = 1
+ w0 = 0
+ ua = -3.1544825e-9
+ ub = 2.30794738e-18
+ uc = 7.77778e-12
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 2.33e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ xrcrg1 = 12
+ xrcrg2 = 1
+ wtvoff = 0
+ tvfbsdoff = 0.022
+ nigbacc = 10
+ capmod = 2
+ tvoff = 0.0057943818
+ wku0we = 2e-11
+ keta = 0.088888889
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ mobmod = 0
+ nigbinv = 10
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 2.3076061000000002e-10
+ kt1l = 0
+ ku0we = -0.0007
+ wkvth0we = 2e-12
+ beta0 = 13
+ leta0 = -1.8441422e-9
+ letab = 4.0459126e-8
+ lint = 0
+ trnqsmod = 0
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ lkt1 = -1.5636766999999998e-8
+ lkt2 = 1.3104778e-9
+ lmax = 5.567e-8
+ lmin = 4.667e-8
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ lpe0 = 9.2e-8
+ fnoimod = 1
+ lpeb = 2.5e-7
+ eigbinv = 1.1
+ minv = -0.3
+ lua1 = 1.2526683e-17
+ lub1 = 1.9957158999999998e-26
+ luc1 = 1.5788889e-17
+ ndep = 1e+18
+ dmcgt = 0
+ rgatemod = 0
+ lwlc = 0
+ tcjsw = 0.000357
+ moin = 5.1
+ tnjtsswg = 1
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ nigc = 3.083
+ bigsd = 0.00125
+ noff = 2.7195
+ cigbacc = 0.32875
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ wvoff = 0
+ tnoimod = 0
+ ntox = 2.029
+ pcit = -1.5e-17
+ pclm = 2.281309
+ wvsat = 0.0
+ wvth0 = -4e-9
+ cigbinv = 0.006
+ phin = 0.15
+ toxref = 3e-9
+ pkt1 = -5e-17
+ lketa = -6.3155556e-9
+ version = 4.5
+ xpart = 1
+ tempmod = 0
+ egidl = 0.29734
+ rbdb = 50
+ prwb = 0
+ pub1 = 0.0
+ prwg = 0
+ )

.model nch_ff_8 nmos (
+ level = 54
+ ngate = 8e+20
+ ngcon = 1
+ wpclm = 0
+ rdsmod = 0
+ wkvth0we = 2e-12
+ wtvfbsdoff = 0
+ igbmod = 1
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ trnqsmod = 0
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ nigbacc = 10
+ ltvfbsdoff = 0
+ pbswgd = 0.95
+ pbswgs = 0.95
+ k2we = 5e-5
+ igcmod = 1
+ dsub = 0.75
+ dtox = 2.7e-10
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ nigbinv = 10
+ rgatemod = 0
+ eta0 = -0.001232
+ etab = -0.88502038
+ tnjtsswg = 1
+ tvfbsdoff = 0.022
+ ptvfbsdoff = 0
+ tvoff = 0.0030235155
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ fnoimod = 1
+ permod = 1
+ eigbinv = 1.1
+ ku0we = -0.0007
+ beta0 = 13
+ leta0 = 1.5454208e-8
+ letab = 3.0054568e-8
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ ppclm = 0
+ voffcv = -0.16942
+ wpemod = 1
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ cigbacc = 0.32875
+ dmcgt = 0
+ tnoimod = 0
+ tcjsw = 0.000357
+ cigbinv = 0.006
+ tpbswg = 0.0009
+ keta = 0.44888889
+ ijthsfwd = 0.01
+ bigsd = 0.00125
+ version = 4.5
+ wvoff = 0
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 5.7703339e-10
+ tempmod = 0
+ kt1l = 0
+ ptvoff = 0
+ wvsat = 0.0
+ wvth0 = -4e-9
+ ijthsrev = 0.01
+ lint = 0
+ aigbacc = 0.02
+ lkt1 = -5.0088498e-9
+ lkt2 = 1.6072e-9
+ diomod = 1
+ lmax = 4.667e-8
+ lmin = 3.6e-8
+ lpe0 = 9.2e-8
+ pditsd = 0
+ pditsl = 0
+ lketa = -2.3955556e-8
+ lpeb = 2.5e-7
+ cjswgd = 2.6226e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.6226e-10
+ xpart = 1
+ minv = -0.3
+ aigbinv = 0.0163
+ lua1 = 7.1708778e-18
+ lub1 = -2.1652990000000025e-27
+ luc1 = -1.63268e-17
+ egidl = 0.29734
+ ndep = 1e+18
+ lwlc = 0
+ mjswgd = 0.85
+ mjswgs = 0.85
+ moin = 5.1
+ nigc = 3.083
+ tcjswg = 0.001
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ poxedge = 1
+ pkvth0we = -1.3e-19
+ ntox = 2.029
+ pcit = -1.5e-17
+ pclm = 2.10165423
+ binunit = 2
+ pvoff = 0
+ fprout = 300
+ phin = 0.15
+ cdscb = 0
+ cdscd = 0
+ vfbsdoff = 0.02
+ pvsat = -1.8e-11
+ xrcrg1 = 12
+ xrcrg2 = 1
+ wk2we = 5e-12
+ pvth0 = -2.3e-16
+ drout = 0.56
+ pkt1 = -5e-17
+ voffl = 0
+ wtvoff = 0
+ paramchk = 1
+ weta0 = 0
+ rbdb = 50
+ prwb = 0
+ pub1 = 0.0
+ prwg = 0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ lpclm = -6.406864000000001e-8
+ rdsw = 100
+ capmod = 2
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ cgidl = 0.22
+ wku0we = 2e-11
+ mobmod = 0
+ ijthdfwd = 0.01
+ a0 = 3.6555556
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 98015.53
+ cf = 8.720500000000001e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.022156861
+ k3 = -1.8419
+ em = 1000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.0035388892999999996
+ pvfbsdoff = 0
+ w0 = 0
+ ua = -2.2580401200000003e-9
+ ub = 1.5627388499999998e-18
+ uc = 2.4e-10
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 2.33e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ pbswd = 0.8
+ pbsws = 0.8
+ rshg = 15.6
+ ijthdrev = 0.01
+ pdits = 0
+ njtsswg = 9
+ cigsd = 0.069865
+ laigsd = -2.1777778e-17
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ ckappad = 0.6
+ ckappas = 0.6
+ pk2we = -1e-19
+ tnom = 25
+ pdiblc1 = 0
+ pdiblc2 = 0.0069157
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ pdiblcb = -0.3
+ toxe = 2.3900000000000002e-9
+ toxm = 2.43e-9
+ tnoia = 0
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ peta0 = 0
+ lkvth0we = -2e-12
+ bigbacc = 0.002588
+ tpbsw = 0.0019
+ wags = -1.5e-8
+ cjswd = 7.625999999999999e-11
+ cjsws = 7.625999999999999e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ wcit = 5e-11
+ kvth0we = 0.00018
+ acnqsmod = 0
+ voff = -0.039834349000000005
+ acde = 0.4
+ lintnoi = -1.5e-8
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ vsat = 69148.62200000002
+ rbodymod = 0
+ vtsswgs = 4.2
+ wint = 0
+ vth0 = 0.372205703
+ toxref = 3e-9
+ wkt1 = -2e-9
+ ags = 2.59253
+ wmax = 0.00090001
+ aigc = 0.011387162
+ wmin = 8.9974e-6
+ cjd = 0.0012620099999999998
+ cit = -0.008475839800000001
+ cjs = 0.0012620099999999998
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 3.26497e-9
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ scref = 1e-6
+ wub1 = 0.0
+ pigcd = 2.621
+ aigsd = 0.010773221
+ la0 = -2.0362223e-7
+ bigc = 0.001442
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.0010317588
+ kt1 = -0.20597876
+ kt2 = -0.11596
+ lk2 = -3.5648647e-9
+ wwlc = 0
+ llc = 0
+ lvoff = -7.176111900000002e-9
+ lln = 1
+ lu0 = 3.7404447e-10
+ mjd = 0.26
+ mjs = 0.26
+ lua = 3.4805321000000004e-17
+ lub = -6.633731000000002e-27
+ luc = -9.7999999e-18
+ lud = 0
+ ltvoff = -1.1163261e-10
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 0
+ nsd = 1e+20
+ pbd = 0.52
+ pat = -2.8e-11
+ pbs = 0.52
+ pk2 = 0
+ lvsat = 0.00197413339
+ cdsc = 0
+ pu0 = 2e-18
+ lvth0 = -1.1825781199999998e-9
+ prt = 0
+ cgbo = 0
+ pua = 0
+ pub = 0
+ puc = 0
+ pud = 0
+ cgdl = 3.5522823e-12
+ cgdo = 5.2490134000000004e-11
+ xtid = 3
+ xtis = 3
+ delta = 0.007595625
+ cgsl = 3.5522823e-12
+ cgso = 5.2490134000000004e-11
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 4.8372486e-10
+ ub1 = -8.3581138e-19
+ cigc = 0.000625
+ laigc = -6.2207351e-12
+ uc1 = 4.882e-10
+ tpb = 0.0014
+ wa0 = 0
+ rnoia = 0
+ rnoib = 0
+ nfactor = 1
+ ute = -1
+ wat = 0.0
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 0
+ wlc = 0
+ lku0we = 2.5e-11
+ wln = 1
+ wu0 = -3.6e-11
+ xgl = -1.09e-8
+ xgw = 0
+ wua = 0
+ wub = 0
+ wuc = 0
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ epsrox = 3.9
+ )

.model nch_ff_9 nmos (
+ level = 54
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ ptvfbsdoff = 0
+ voffl = 0
+ minv = -0.3
+ lub1 = 0
+ weta0 = 0
+ ndep = 1e+18
+ wetab = -1.0073378e-8
+ lwlc = 0
+ moin = 5.1
+ nigc = 3.083
+ cgidl = 0.22
+ lkvth0we = -2e-12
+ njtsswg = 9
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ pvfbsdoff = 0
+ noic = 45200000.0
+ permod = 1
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ acnqsmod = 0
+ pbswd = 0.8
+ pbsws = 0.8
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.018557155
+ pdiblcb = -0.3
+ ntox = 2.029
+ pcit = -1.5e-17
+ pclm = 1.4152454
+ rbodymod = 0
+ phin = 0.15
+ voffcv = -0.16942
+ wpemod = 1
+ pdits = 0
+ cigsd = 0.069865
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ pkt1 = -5e-17
+ bigbacc = 0.002588
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ kvth0we = 0.00018
+ rbdb = 50
+ prwb = 0
+ pub1 = 0
+ prwg = 0
+ wpdiblc2 = -1.7177628e-11
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ lintnoi = -1.5e-8
+ tnoia = 0
+ bigbinv = 0.004953
+ rdsw = 100
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ peta0 = 0
+ tpbswg = 0.0009
+ wketa = 3.3422159e-8
+ tpbsw = 0.0019
+ cjswd = 7.625999999999999e-11
+ cjsws = 7.625999999999999e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ ags = 0.80683314
+ ptvoff = 0
+ cjd = 0.0012620099999999998
+ cit = 4.8708935e-5
+ cjs = 0.0012620099999999998
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ wkvth0we = 2e-12
+ bvs = 8.7
+ rshg = 15.6
+ waigsd = 3.0716751e-12
+ dlc = 9.8024918e-9
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ trnqsmod = 0
+ diomod = 1
+ la0 = 0
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.0001
+ kt1 = -0.19515831
+ kt2 = -0.052853133
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 2.6226e-10
+ llc = 0
+ pku0we = -1.5e-18
+ lln = 1
+ cjswgs = 2.6226e-10
+ lu0 = 6e-12
+ mjd = 0.26
+ mjs = 0.26
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ scref = 1e-6
+ njd = 1.02
+ njs = 1.02
+ pa0 = 0
+ nfactor = 1
+ nsd = 1e+20
+ pbd = 0.52
+ pat = -2.8e-11
+ pbs = 0.52
+ pigcd = 2.621
+ aigsd = 0.010772879
+ pu0 = 2e-18
+ prt = 0
+ pud = 0
+ tnom = 25
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 1.311952e-9
+ toxe = 2.3900000000000002e-9
+ ub1 = -8.0649865e-19
+ toxm = 2.43e-9
+ lvoff = -2e-11
+ uc1 = 3.0375074e-11
+ mjswgd = 0.85
+ mjswgs = 0.85
+ tpb = 0.0014
+ rgatemod = 0
+ wa0 = -2.5183444e-7
+ ute = -0.96248296
+ wat = 0
+ tnjtsswg = 1
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -3.7920026e-9
+ lvsat = -0.0003
+ wlc = 0
+ tcjswg = 0.001
+ wln = 1
+ wu0 = -2.9790781999999996e-10
+ xgl = -1.09e-8
+ xgw = 0
+ lvth0 = -1e-10
+ wua = -4.0765791e-17
+ wub = 4.0599742e-26
+ wuc = -7.8572347e-18
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ delta = 0.007595625
+ nigbacc = 10
+ rnoia = 0
+ rnoib = 0
+ wags = -9.9054279e-8
+ wcit = 5.1192733e-10
+ ngate = 8e+20
+ voff = -0.11308442
+ ngcon = 1
+ wpclm = -1.3730014e-7
+ acde = 0.4
+ nigbinv = 10
+ vsat = 103058.98
+ wint = 0
+ gbmin = 1e-12
+ vth0 = 0.32234844999999995
+ fprout = 300
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ wkt1 = -4.7639654e-8
+ wkt2 = -3.5741805e-9
+ wmax = 8.9974e-6
+ xrcrg1 = 12
+ xrcrg2 = 1
+ aigc = 0.011766468
+ wmin = 8.974e-7
+ wtvoff = -8.3463378e-10
+ wua1 = -7.3834184e-16
+ wub1 = 7.3798399e-25
+ wuc1 = -8.5623711e-19
+ fnoimod = 1
+ bigc = 0.001442
+ wute = -4.0092044e-7
+ eigbinv = 1.1
+ wwlc = 0
+ tvfbsdoff = 0.022
+ capmod = 2
+ cdsc = 0
+ cgbo = 0
+ wku0we = 2e-11
+ cgdl = 3.5522823e-12
+ cgdo = 5.2490134000000004e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.5522823e-12
+ cgso = 5.2490134000000004e-11
+ tvoff = 0.0020036382
+ cigc = 0.000625
+ mobmod = 0
+ xjbvd = 1
+ ijthsfwd = 0.01
+ xjbvs = 1
+ lk2we = -1.5e-12
+ cigbacc = 0.32875
+ ku0we = -0.0007
+ beta0 = 13
+ leta0 = 0
+ tnoimod = 0
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ ijthsrev = 0.01
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ cigbinv = 0.006
+ dlcig = 2.5e-9
+ k2we = 5e-5
+ bgidl = 2320000000.0
+ dsub = 0.75
+ dtox = 2.7e-10
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ a0 = 3.277963
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ version = 4.5
+ at = 72000
+ cf = 8.720500000000001e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.023022307
+ k3 = -1.8419
+ em = 1000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.015299082
+ dmcgt = 0
+ w0 = 0
+ tempmod = 0
+ ua = -1.8192461e-9
+ ub = 2.0991879e-18
+ uc = 7.4172444e-11
+ ud = 0
+ eta0 = 0.3
+ tcjsw = 0.000357
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 2.33e-9
+ alpha0 = 2e-10
+ ww = 0
+ alpha1 = 3.6
+ xw = 8.600000000000001e-9
+ etab = -0.24888148
+ aigbacc = 0.02
+ bigsd = 0.00125
+ wvoff = 2.3777201e-9
+ pkvth0we = -1.3e-19
+ aigbinv = 0.0163
+ wvsat = -0.0017920539
+ wvth0 = -1.5145485e-8
+ toxref = 3e-9
+ waigc = 2.6350949e-11
+ vfbsdoff = 0.02
+ xpart = 1
+ paramchk = 1
+ ltvoff = 0
+ egidl = 0.29734
+ poxedge = 1
+ binunit = 2
+ wtvfbsdoff = 0
+ keta = -0.063711099
+ lku0we = 2.5e-11
+ ijthdfwd = 0.01
+ epsrox = 3.9
+ ltvfbsdoff = 0
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = -1e-11
+ rdsmod = 0
+ kt1l = 0
+ igbmod = 1
+ ijthdrev = 0.01
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ pvoff = 0
+ lint = 6.5375218e-9
+ pbswgd = 0.95
+ cdscb = 0
+ cdscd = 0
+ pbswgs = 0.95
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ lkt1 = -1.1e-9
+ pvsat = -1.8e-11
+ lmax = 2.001e-5
+ wk2we = 5e-12
+ pvth0 = -2.3e-16
+ lmin = 9.00077e-6
+ drout = 0.56
+ igcmod = 1
+ )

.model nch_ff_10 nmos (
+ level = 54
+ xrcrg1 = 12
+ xrcrg2 = 1
+ cgidl = 0.22
+ vfbsdoff = 0.02
+ wtvoff = -8.9580408e-10
+ nfactor = 1
+ pbswd = 0.8
+ pbsws = 0.8
+ paramchk = 1
+ capmod = 2
+ wku0we = 2e-11
+ mobmod = 0
+ pdits = 0
+ cigsd = 0.069865
+ nigbacc = 10
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ ijthdfwd = 0.01
+ keta = -0.064075044
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ nigbinv = 10
+ lags = -6.3328546e-8
+ wtvfbsdoff = 0
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 1.1237416e-9
+ tnoia = 0
+ laigsd = 1.1048614e-17
+ ijthdrev = 0.01
+ kt1l = 0
+ peta0 = 0
+ ltvfbsdoff = 0
+ lpdiblc2 = -6.1589259e-10
+ wketa = 3.7630763e-8
+ lint = 6.5375218e-9
+ tpbsw = 0.0019
+ lkt1 = -4.6637316000000004e-8
+ lkt2 = -1.2972142e-8
+ cjswd = 7.625999999999999e-11
+ lmax = 9.00077e-6
+ cjsws = 7.625999999999999e-11
+ lmin = 9.0075e-7
+ fnoimod = 1
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ lpe0 = 9.2e-8
+ eigbinv = 1.1
+ lpeb = 2.5e-7
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ minv = -0.3
+ lua1 = -4.3996966e-16
+ lub1 = 2.6060002e-25
+ luc1 = 3.9191378e-17
+ ndep = 1e+18
+ lute = -3.7058959e-8
+ lwlc = 0
+ ptvfbsdoff = 0
+ moin = 5.1
+ lkvth0we = -2e-12
+ nigc = 3.083
+ scref = 1e-6
+ pigcd = 2.621
+ aigsd = 0.010772879
+ cigbacc = 0.32875
+ acnqsmod = 0
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ lvoff = -1.4262682e-8
+ toxref = 3e-9
+ tnoimod = 0
+ pags = 2.8299487e-13
+ rbodymod = 0
+ lvsat = -0.0003
+ lvth0 = 5.1155324e-8
+ ntox = 2.029
+ pcit = -1.996418e-16
+ pclm = 1.4152454
+ cigbinv = 0.006
+ delta = 0.007595625
+ laigc = -1.4938914e-10
+ tvfbsdoff = 0.022
+ rnoia = 0
+ rnoib = 0
+ phin = 0.15
+ pkt1 = 4.9822912e-14
+ pkt2 = 1.3351872e-15
+ pketa = -3.7835355e-14
+ version = 4.5
+ ngate = 8e+20
+ ltvoff = -2.0733557e-10
+ ngcon = 1
+ tempmod = 0
+ wpclm = -1.3730014e-7
+ wpdiblc2 = -4.8108443e-11
+ gbmin = 1e-12
+ rbdb = 50
+ pua1 = 6.0905252e-22
+ prwb = 0
+ prwg = 0
+ pub1 = -5.9738158e-31
+ jswgd = 1.28e-13
+ puc1 = 1.7562426e-23
+ jswgs = 1.28e-13
+ rbpb = 50
+ rbpd = 50
+ aigbacc = 0.02
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ pute = 3.9602525e-13
+ lku0we = 2.5e-11
+ rdsw = 100
+ wvfbsdoff = 0
+ epsrox = 3.9
+ lvfbsdoff = 0
+ rdsmod = 0
+ aigbinv = 0.0163
+ igbmod = 1
+ wkvth0we = 2e-12
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ pbswgd = 0.95
+ pbswgs = 0.95
+ rshg = 15.6
+ trnqsmod = 0
+ tvoff = 0.0020267011
+ igcmod = 1
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ poxedge = 1
+ ku0we = -0.0007
+ beta0 = 13
+ tnom = 25
+ rgatemod = 0
+ leta0 = 0
+ binunit = 2
+ tnjtsswg = 1
+ toxe = 2.3900000000000002e-9
+ paigsd = -9.9503825e-23
+ toxm = 2.43e-9
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ permod = 1
+ wags = -1.3053313e-7
+ wcit = 5.3246591e-10
+ dmcgt = 0
+ tcjsw = 0.000357
+ voff = -0.11150014
+ acde = 0.4
+ voffcv = -0.16942
+ wpemod = 1
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ vsat = 103058.98
+ wint = 0
+ vth0 = 0.31664707999999997
+ wkt1 = -5.3187252999999996e-8
+ wkt2 = -3.7226997e-9
+ wmax = 8.9974e-6
+ aigc = 0.011783086
+ bigsd = 0.00125
+ wmin = 8.974e-7
+ wvoff = 2.6904676e-9
+ wua1 = -8.0608962e-16
+ wub1 = 8.0443355e-25
+ wuc1 = -2.8097884e-18
+ wvsat = -0.0017920539
+ wvth0 = -1.5528173e-8
+ bigc = 0.001442
+ wute = -4.4497219e-7
+ wwlc = 0
+ waigc = 2.7413515e-11
+ tpbswg = 0.0009
+ njtsswg = 9
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.5522823e-12
+ cgdo = 5.2490134000000004e-11
+ xtid = 3
+ xtis = 3
+ lketa = 3.2718606e-9
+ xtsswgd = 0.18
+ cgsl = 3.5522823e-12
+ ijthsfwd = 0.01
+ cgso = 5.2490134000000004e-11
+ xtsswgs = 0.18
+ cigc = 0.000625
+ xpart = 1
+ ckappad = 0.6
+ ckappas = 0.6
+ ptvoff = 5.4992103e-16
+ pdiblc1 = 0
+ pdiblc2 = 0.018625664
+ pdiblcb = -0.3
+ waigsd = 3.0716862e-12
+ egidl = 0.29734
+ diomod = 1
+ ijthsrev = 0.01
+ pditsd = 0
+ pditsl = 0
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ cjswgd = 2.6226e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.6226e-10
+ ags = 0.81387747
+ bigbacc = 0.002588
+ cjd = 0.0012620099999999998
+ cit = -7.7402473e-5
+ cjs = 0.0012620099999999998
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 9.8024918e-9
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ k2we = 5e-5
+ kvth0we = 0.00018
+ dsub = 0.75
+ dtox = 2.7e-10
+ mjswgd = 0.85
+ mjswgs = 0.85
+ pvfbsdoff = 0
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ la0 = -2.0592205e-6
+ lintnoi = -1.5e-8
+ ppdiblc2 = 2.7806803e-16
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = 0.094382725
+ tcjswg = 0.001
+ kt1 = -0.19009298
+ lk2 = -1.3154073e-8
+ kt2 = -0.051410181
+ bigbinv = 0.004953
+ llc = 0
+ vtsswgd = 4.2
+ lln = 1
+ vtsswgs = 4.2
+ lu0 = -1.9904409e-9
+ mjd = 0.26
+ lua = -2.2049077e-16
+ mjs = 0.26
+ lub = -1.5408759e-27
+ luc = 1.1211784e-18
+ lud = 0
+ pvoff = -2.8116001e-15
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 3.0846188e-13
+ eta0 = 0.3
+ nsd = 1e+20
+ pbd = 0.52
+ pat = -8.306718700000001e-9
+ pbs = 0.52
+ pk2 = -1.9754424e-15
+ cdscb = 0
+ cdscd = 0
+ etab = -0.24888148
+ pu0 = 1.19503831e-17
+ pvsat = -1.8e-11
+ prt = 0
+ pua = 2.7693259e-23
+ pub = -6.3482817e-32
+ puc = -1.7214163e-23
+ pud = 0
+ wk2we = 5e-12
+ pvth0 = 3.2103638999999997e-15
+ drout = 0.56
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 1.3608919e-9
+ ub1 = -8.3548641e-19
+ uc1 = 2.6015633e-11
+ paigc = -9.5524673e-18
+ tpb = 0.0014
+ wa0 = -2.8614611e-7
+ ute = -0.95836072
+ wat = 0.00092088084
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -3.5722648e-9
+ voffl = 0
+ wlc = 0
+ wln = 1
+ wu0 = -2.9901464999999997e-10
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -4.3846243e-17
+ wub = 4.7661234e-26
+ wuc = -5.9424224e-18
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ a0 = 3.5070197
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ weta0 = 0
+ pkvth0we = -1.3e-19
+ at = 61490.242
+ cf = 8.720500000000001e-11
+ wetab = -1.0073378e-8
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.024485497000000002
+ k3 = -1.8419
+ em = 1000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.015521155
+ fprout = 300
+ w0 = 0
+ ua = -1.7947198e-9
+ ub = 2.0993593e-18
+ uc = 7.4047731e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 2.33e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ )

.model nch_ff_11 nmos (
+ level = 54
+ ku0we = -0.0007
+ beta0 = 13
+ wku0we = 2e-11
+ leta0 = 0
+ rbdb = 50
+ mobmod = 0
+ pua1 = 9.7840116e-23
+ prwb = 0
+ prwg = 0
+ pub1 = -1.2240721e-31
+ puc1 = -3.5940917e-24
+ a0 = 1.2386098
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ wtvfbsdoff = 0
+ at = 220073.87
+ cf = 8.720500000000001e-11
+ rbpb = 50
+ rbpd = 50
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.023732722999999997
+ k3 = -1.8419
+ rbps = 50
+ em = 1000000.0
+ rbsb = 50
+ pvag = 1.2
+ ll = 0
+ lw = 0
+ u0 = 0.015021688
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ w0 = 0
+ ua = -1.9419497e-9
+ ub = 2.1613601e-18
+ uc = 9.7509556e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 2.33e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ rdsw = 100
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ ijthsfwd = 0.01
+ ltvfbsdoff = 0
+ dmcgt = 0
+ tcjsw = 0.000357
+ laigsd = -9.7335958e-18
+ ijthsrev = 0.01
+ rshg = 15.6
+ njtsswg = 9
+ bigsd = 0.00125
+ ptvfbsdoff = 0
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ wvoff = -7.7864574e-9
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.014827337
+ pdiblcb = -0.3
+ wvsat = -0.0017920539
+ ppdiblc2 = 2.4623293e-15
+ tnom = 25
+ wvth0 = -5.226189400000001e-9
+ toxe = 2.3900000000000002e-9
+ toxm = 2.43e-9
+ waigc = -9.5733062e-12
+ lketa = -3.0044615e-8
+ bigbacc = 0.002588
+ xpart = 1
+ wags = 1.2310313e-6
+ kvth0we = 0.00018
+ toxref = 3e-9
+ egidl = 0.29734
+ pkvth0we = -1.3e-19
+ wcit = 2.0976377e-10
+ ags = 0.16741392
+ cjd = 0.0012620099999999998
+ cit = 0.0013334381
+ voff = -0.11121991
+ lintnoi = -1.5e-8
+ cjs = 0.0012620099999999998
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ acde = 0.4
+ dlc = 9.8024918e-9
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ k3b = 1.9326
+ vtsswgs = 4.2
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ vsat = 103058.98
+ wint = 0
+ vfbsdoff = 0.02
+ vth0 = 0.36519506999999996
+ wkt1 = 1.5828642999999998e-8
+ wkt2 = -3.7425887e-9
+ wmax = 8.9974e-6
+ la0 = -4.0335612e-8
+ aigc = 0.011680759
+ wmin = 8.974e-7
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.046756700000000005
+ kt1 = -0.22273968
+ lk2 = -1.2484105e-8
+ kt2 = -0.052902736
+ llc = 0
+ lln = 1
+ lu0 = -1.5459156e-9
+ mjd = 0.26
+ ltvoff = -6.7137092e-10
+ lua = -8.9456155e-17
+ mjs = 0.26
+ lub = -5.6721601e-26
+ luc = -1.9759846e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = -3.420874e-13
+ nsd = 1e+20
+ pbd = 0.52
+ pat = -3.6746881e-9
+ pbs = 0.52
+ pk2 = 6.3553328e-16
+ pvfbsdoff = 0
+ paramchk = 1
+ pu0 = 2.8298232e-17
+ wua1 = -2.3169366e-16
+ wub1 = 2.7075449e-25
+ prt = 0
+ wuc1 = 2.096158e-17
+ pua = -3.3732216e-24
+ pub = 1.7089792e-32
+ puc = 7.8894695e-24
+ pud = 0
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 9.9427719e-10
+ bigc = 0.001442
+ ub1 = -5.7879508e-19
+ uc1 = 6.536871e-11
+ pvoff = 6.5128631e-15
+ tpb = 0.0014
+ wwlc = 0
+ wa0 = 4.4480813e-7
+ ute = -1
+ wat = -0.0042836479
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -6.5059453e-9
+ cdscb = 0
+ cdscd = 0
+ lku0we = 2.5e-11
+ wlc = 0
+ wln = 1
+ wu0 = -3.1738301999999995e-10
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -8.9400845e-18
+ wub = -4.2869787e-26
+ pvsat = -1.8e-11
+ wuc = -3.4148751e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ epsrox = 3.9
+ cdsc = 0
+ wk2we = 5e-12
+ pvth0 = -5.9584018000000004e-15
+ drout = 0.56
+ cgbo = 0
+ cgdl = 3.5522823e-12
+ cgdo = 5.2490134000000004e-11
+ xtid = 3
+ xtis = 3
+ ijthdfwd = 0.01
+ cgsl = 3.5522823e-12
+ paigc = 2.3365803e-17
+ cgso = 5.2490134000000004e-11
+ cigc = 0.000625
+ rdsmod = 0
+ nfactor = 1
+ voffl = 0
+ igbmod = 1
+ weta0 = 0
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ wetab = -1.0073378e-8
+ pbswgd = 0.95
+ pbswgs = 0.95
+ ijthdrev = 0.01
+ igcmod = 1
+ cgidl = 0.22
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ lpdiblc2 = 2.7646188e-9
+ nigbacc = 10
+ k2we = 5e-5
+ pbswd = 0.8
+ pbsws = 0.8
+ dsub = 0.75
+ dtox = 2.7e-10
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ nigbinv = 10
+ paigsd = 8.7660773e-23
+ eta0 = 0.3
+ pdits = 0
+ etab = -0.24888148
+ cigsd = 0.069865
+ lkvth0we = -2e-12
+ permod = 1
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ pk2we = -1e-19
+ fnoimod = 1
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ acnqsmod = 0
+ eigbinv = 1.1
+ voffcv = -0.16942
+ wpemod = 1
+ tnoia = 0
+ rbodymod = 0
+ peta0 = 0
+ wketa = -4.0591301e-8
+ tpbsw = 0.0019
+ cjswd = 7.625999999999999e-11
+ cjsws = 7.625999999999999e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ cigbacc = 0.32875
+ wpdiblc2 = -2.5023346e-9
+ tnoimod = 0
+ tpbswg = 0.0009
+ cigbinv = 0.006
+ scref = 1e-6
+ ptvoff = 2.4706364e-16
+ pigcd = 2.621
+ keta = -0.026640801
+ aigsd = 0.010772879
+ waigsd = 3.0714759e-12
+ version = 4.5
+ lvoff = -1.4512080999999999e-8
+ lags = 5.1202402e-7
+ wkvth0we = 2e-12
+ tempmod = 0
+ jswd = 1.28e-13
+ diomod = 1
+ jsws = 1.28e-13
+ lcit = -1.3190653e-10
+ lvsat = -0.0003
+ kt1l = 0
+ lvth0 = 7.947615400000001e-9
+ pditsd = 0
+ pditsl = 0
+ trnqsmod = 0
+ cjswgd = 2.6226e-10
+ tvfbsdoff = 0.022
+ pku0we = -1.5e-18
+ cjswgs = 2.6226e-10
+ delta = 0.007595625
+ laigc = -5.8318716e-11
+ aigbacc = 0.02
+ lint = 6.5375218e-9
+ rnoia = 0
+ rnoib = 0
+ lkt1 = -1.7581753e-8
+ lkt2 = -1.1643768e-8
+ lmax = 9.0075e-7
+ lmin = 4.5075e-7
+ pketa = 3.1782283e-14
+ mjswgd = 0.85
+ lpe0 = 9.2e-8
+ ngate = 8e+20
+ mjswgs = 0.85
+ lpeb = 2.5e-7
+ ngcon = 1
+ wpclm = -1.3730014e-7
+ aigbinv = 0.0163
+ tcjswg = 0.001
+ minv = -0.3
+ rgatemod = 0
+ lua1 = -1.1368255e-16
+ lub1 = 3.2144732e-26
+ luc1 = 4.1671397e-18
+ gbmin = 1e-12
+ tnjtsswg = 1
+ ndep = 1e+18
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ lwlc = 0
+ moin = 5.1
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ nigc = 3.083
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ poxedge = 1
+ fprout = 300
+ xrcrg1 = 12
+ xrcrg2 = 1
+ pags = -9.2879744e-13
+ ntox = 2.029
+ pcit = 8.756310000000001e-17
+ binunit = 2
+ pclm = 1.4152454
+ tvoff = 0.0025480892
+ wtvoff = -5.5551488e-10
+ xjbvd = 1
+ phin = 0.15
+ xjbvs = 1
+ lk2we = -1.5e-12
+ pkt1 = -1.1601235000000001e-14
+ pkt2 = 1.3528884e-15
+ capmod = 2
+ )

.model nch_ff_12 nmos (
+ level = 54
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ ptvfbsdoff = 0
+ cigbacc = 0.32875
+ laigsd = -9.015225e-17
+ wkvth0we = 2e-12
+ tnoia = 0
+ tnoimod = 0
+ trnqsmod = 0
+ peta0 = 0
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ wketa = 1.7936379e-8
+ tpbsw = 0.0019
+ a0 = 1.7327189
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ cigbinv = 0.006
+ at = 153009.14
+ cf = 8.720500000000001e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.017241707000000002
+ k3 = -1.8419
+ em = 1000000.0
+ cjswd = 7.625999999999999e-11
+ ll = -1.18e-13
+ cjsws = 7.625999999999999e-11
+ lw = 0
+ u0 = 0.012915621
+ w0 = 0
+ mjswd = 0.11
+ ua = -2.1226101e-9
+ ub = 2.1428106e-18
+ uc = 6.8443458e-11
+ ud = 0
+ mjsws = 0.11
+ agidl = 9.41e-8
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 2.33e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ k2we = 5e-5
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ dsub = 0.75
+ dtox = 2.7e-10
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ version = 4.5
+ rgatemod = 0
+ tnjtsswg = 1
+ tempmod = 0
+ eta0 = 0.3
+ etab = -0.24888148
+ aigbacc = 0.02
+ scref = 1e-6
+ pigcd = 2.621
+ aigsd = 0.010772879
+ toxref = 3e-9
+ lvoff = -6.1111145e-9
+ aigbinv = 0.0163
+ lvsat = -0.0003
+ lvth0 = -5.041492e-9
+ tvfbsdoff = 0.022
+ delta = 0.007595625
+ laigc = -1.9233809e-11
+ rnoia = 0
+ rnoib = 0
+ ltvoff = -1.0250882e-10
+ pketa = 6.0301037e-15
+ ngate = 8e+20
+ ngcon = 1
+ wpclm = -2.8227848e-7
+ poxedge = 1
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ lku0we = 2.5e-11
+ wvfbsdoff = 0
+ epsrox = 3.9
+ lvfbsdoff = 0
+ binunit = 2
+ rdsmod = 0
+ ijthsfwd = 0.01
+ igbmod = 1
+ keta = -0.041938217
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ lags = 4.5664516e-7
+ pbswgd = 0.95
+ pbswgs = 0.95
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 1.5914929e-10
+ ijthsrev = 0.01
+ igcmod = 1
+ kt1l = 0
+ tvoff = 0.0012552207
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ lint = 9.7879675e-9
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ lkt1 = -1.06958544e-8
+ lkt2 = -3.7159363e-9
+ lmax = 4.5075e-7
+ lmin = 2.1744e-7
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ ku0we = -0.0007
+ paigsd = 8.167794e-23
+ ppdiblc2 = -2.773275e-15
+ beta0 = 13
+ minv = -0.3
+ lua1 = -3.2594611e-17
+ lub1 = -2.740043e-26
+ leta0 = 0
+ luc1 = -3.5163101e-18
+ ndep = 1e+18
+ ppclm = 6.379047e-14
+ lwlc = 0
+ permod = 1
+ moin = 5.1
+ dlcig = 2.5e-9
+ nigc = 3.083
+ bgidl = 2320000000.0
+ njtsswg = 9
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ pkvth0we = -1.3e-19
+ dmcgt = 0
+ voffcv = -0.16942
+ ckappad = 0.6
+ wpemod = 1
+ ckappas = 0.6
+ tcjsw = 0.000357
+ pdiblc1 = 0
+ pdiblc2 = 0.026288388
+ pags = 8.4375107e-13
+ pdiblcb = -0.3
+ ntox = 2.029
+ pcit = -7.789201199999999e-17
+ pclm = 1.5752657
+ vfbsdoff = 0.02
+ phin = 0.15
+ bigsd = 0.00125
+ pkt1 = -5.274892300000001e-16
+ pkt2 = -1.2933793e-15
+ bigbacc = 0.002588
+ wvoff = 1.1733398e-8
+ paramchk = 1
+ wvsat = -0.0017920539
+ kvth0we = 0.00018
+ wvth0 = -2.3374896e-8
+ tpbswg = 0.0009
+ rbdb = 50
+ pua1 = 1.9082335e-23
+ prwb = 0
+ prwg = 0
+ pub1 = -2.3158905e-32
+ puc1 = -7.9472634e-24
+ waigc = 5.7897385e-11
+ lintnoi = -1.5e-8
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ rdsw = 100
+ ags = 0.29327496999999997
+ lketa = -2.3313752e-8
+ ijthdfwd = 0.01
+ ptvoff = -1.6297696e-16
+ xpart = 1
+ cjd = 0.0012620099999999998
+ cit = 0.00067194759
+ cjs = 0.0012620099999999998
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ waigsd = 3.0714895e-12
+ dlc = 1.30529375e-8
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ egidl = 0.29734
+ diomod = 1
+ la0 = -2.5774361e-7
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.017248219
+ pditsd = 0
+ pditsl = 0
+ kt1 = -0.23838945
+ ijthdrev = 0.01
+ lk2 = -9.6280577e-9
+ kt2 = -0.070920535
+ cjswgd = 2.6226e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.6226e-10
+ llc = -1.18e-13
+ lln = 0.7
+ rshg = 15.6
+ lu0 = -6.192457900000001e-10
+ mjd = 0.26
+ lua = -9.9655811e-18
+ mjs = 0.26
+ lub = -4.8559819e-26
+ luc = -6.9707629e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 9.4027643e-14
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 2.5203517e-9
+ lpdiblc2 = -2.2782436e-9
+ pbs = 0.52
+ pk2 = 9.5548939e-17
+ pu0 = 1.01677938e-17
+ prt = 0
+ pua = -7.1355685e-24
+ pub = 6.4921301e-33
+ puc = 2.8995668e-24
+ pud = 0
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 8.0998641e-10
+ ub1 = -4.4346517e-19
+ uc1 = 8.2831095e-11
+ mjswgd = 0.85
+ mjswgs = 0.85
+ tpb = 0.0014
+ wa0 = -5.4636242e-7
+ nfactor = 1
+ pvfbsdoff = 0
+ ute = -1
+ wat = -0.018363284
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -5.2787082e-9
+ tcjswg = 0.001
+ wlc = 0
+ wln = 1
+ wu0 = -2.7617747999999996e-10
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -3.8929611e-19
+ wub = -1.8784192e-26
+ wuc = -2.2808063e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ tnom = 25
+ pvoff = -2.0758734e-15
+ toxe = 2.3900000000000002e-9
+ toxm = 2.43e-9
+ cdscb = 0
+ cdscd = 0
+ lkvth0we = -2e-12
+ pvsat = -1.8e-11
+ wk2we = 5e-12
+ pvth0 = 2.0270293000000002e-15
+ drout = 0.56
+ paigc = -6.3213007e-18
+ nigbacc = 10
+ voffl = 0
+ acnqsmod = 0
+ wags = -2.7974881e-6
+ fprout = 300
+ weta0 = 0
+ wetab = -1.0073378e-8
+ wcit = 5.8579813e-10
+ xrcrg1 = 12
+ xrcrg2 = 1
+ lpclm = -7.0408907e-8
+ voff = -0.13031302
+ rbodymod = 0
+ nigbinv = 10
+ acde = 0.4
+ cgidl = 0.22
+ vsat = 103058.98
+ wtvoff = 3.7639557e-10
+ wint = 0
+ vth0 = 0.39471576999999997
+ wkt1 = -9.3389616e-9
+ wkt2 = 2.2716562e-9
+ wmax = 8.9974e-6
+ wtvfbsdoff = 0
+ aigc = 0.01159193
+ wmin = 8.974e-7
+ capmod = 2
+ pbswd = 0.8
+ pbsws = 0.8
+ ltvfbsdoff = 0
+ fnoimod = 1
+ wua1 = -5.2698704e-17
+ wub1 = 4.5190152e-26
+ wku0we = 2e-11
+ wuc1 = 3.0855152e-17
+ eigbinv = 1.1
+ wpdiblc2 = 9.3967661e-9
+ bigc = 0.001442
+ mobmod = 0
+ wwlc = 0
+ pdits = 0
+ cigsd = 0.069865
+ cdsc = 0
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ cgbo = 0
+ cgdl = 3.5522823e-12
+ cgdo = 5.2490134000000004e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.5522823e-12
+ cgso = 5.2490134000000004e-11
+ cigc = 0.000625
+ )

.model nch_ff_13 nmos (
+ level = 54
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ lint = 9.7879675e-9
+ bigsd = 0.00125
+ lkt1 = -4.721126e-9
+ lkt2 = -5.6046527e-10
+ lmax = 2.1744e-7
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ lmin = 9.167e-8
+ wvoff = -2.233608000000001e-9
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ wvsat = -0.00035982647999999954
+ minv = -0.3
+ wvth0 = -9.862616999999999e-9
+ lua1 = 8.0644671e-18
+ lub1 = -5.2760301e-26
+ luc1 = -4.6427809e-18
+ ags = 2.4574682
+ ndep = 1e+18
+ waigc = 3.6164887e-11
+ cjd = 0.0012620099999999998
+ cit = 0.0010410649
+ cjs = 0.0012620099999999998
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ lwlc = 0
+ dlc = 1.30529375e-8
+ k3b = 1.9326
+ moin = 5.1
+ lkvth0we = -2e-12
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ nigc = 3.083
+ lketa = -1.0074554e-8
+ xpart = 1
+ la0 = -3.95931149e-8
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.0019760989
+ toxref = 3e-9
+ kt1 = -0.26670569
+ lk2 = -2.2996724e-9
+ kt2 = -0.085875374
+ llc = -1.18e-13
+ lln = 0.7
+ a0 = 0.69883298
+ a1 = 0
+ a2 = 1
+ lu0 = -1.9339705999999998e-10
+ b0 = 0
+ b1 = 0
+ acnqsmod = 0
+ mjd = 0.26
+ lua = 2.3685126e-17
+ mjs = 0.26
+ lub = -3.581049857e-26
+ luc = -1.971816e-18
+ lud = 0
+ at = 80629.42
+ cf = 8.720500000000001e-11
+ lwc = 0
+ noff = 2.7195
+ lwl = 0
+ lwn = 1
+ ef = 1.0
+ k1 = 0.274
+ k2 = -0.017489977
+ k3 = -1.8419
+ em = 1000000.0
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ njd = 1.02
+ njs = 1.02
+ nfactor = 1
+ pa0 = 5.1229998e-14
+ egidl = 0.29734
+ ll = -1.18e-13
+ lw = 0
+ u0 = 0.01089738
+ w0 = 0
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 7.9357566e-10
+ pbs = 0.52
+ ua = -2.2820921e-9
+ ub = 2.0823870489000003e-18
+ uc = 4.4751766e-11
+ ud = 0
+ pk2 = 1.6389978e-16
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 2.33e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ pu0 = -2.0541017e-17
+ prt = 0
+ pua = 6.5907354e-24
+ pub = -1.1536808500000001e-32
+ puc = -4.2264406e-24
+ pud = 0
+ pags = -3.4153056e-19
+ rbodymod = 0
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 6.1728936e-10
+ ub1 = -3.2327621e-19
+ uc1 = 8.8169819e-11
+ ntox = 2.029
+ pcit = -7.5109378e-17
+ pclm = 1.3619854
+ tpb = 0.0014
+ wa0 = -3.4353242e-7
+ ute = -1
+ wat = -0.010179511
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -5.6026458e-9
+ wlc = 0
+ wln = 1
+ wu0 = -1.30638093e-10
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -6.5442869e-17
+ wub = 6.6660889e-26
+ wuc = 1.0964484e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ ltvoff = 4.8985213e-12
+ phin = 0.15
+ pvfbsdoff = 0
+ nigbacc = 10
+ pkt1 = 2.7743122e-15
+ pkt2 = -3.7226831e-16
+ wpdiblc2 = -7.3538749e-9
+ lku0we = 2.5e-11
+ pvoff = 8.711494700000001e-16
+ rbdb = 50
+ pua1 = -3.4072796e-24
+ prwb = 0
+ prwg = 0
+ pub1 = 3.7649133e-33
+ epsrox = 3.9
+ puc1 = 3.7978198e-24
+ cdscb = 0
+ cdscd = 0
+ rbpb = 50
+ rbpd = 50
+ nigbinv = 10
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ pvsat = -3.2019949e-10
+ wk2we = 5e-12
+ pvth0 = -8.240435999999998e-16
+ rdsw = 100
+ drout = 0.56
+ rdsmod = 0
+ igbmod = 1
+ paigc = -1.7357437e-18
+ voffl = 0
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ pbswgd = 0.95
+ pbswgs = 0.95
+ weta0 = 0
+ wetab = -1.0073378e-8
+ wkvth0we = 2e-12
+ fnoimod = 1
+ lpclm = -2.540677e-8
+ igcmod = 1
+ eigbinv = 1.1
+ rshg = 15.6
+ trnqsmod = 0
+ cgidl = 0.22
+ pbswd = 0.8
+ pbsws = 0.8
+ paigsd = -5.1229584e-23
+ rgatemod = 0
+ tnom = 25
+ cigbacc = 0.32875
+ tnjtsswg = 1
+ toxe = 2.3900000000000002e-9
+ toxm = 2.43e-9
+ permod = 1
+ pdits = 0
+ cigsd = 0.069865
+ tnoimod = 0
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ cigbinv = 0.006
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ wags = 1.2013337999999998e-6
+ voffcv = -0.16942
+ wpemod = 1
+ wcit = 5.726102800000001e-10
+ tnoia = 0
+ voff = -0.1572150866
+ version = 4.5
+ acde = 0.4
+ tempmod = 0
+ peta0 = 0
+ vsat = 102561.23895
+ wint = 0
+ vth0 = 0.4092123399
+ wketa = 1.0437078e-7
+ wkt1 = -2.498731e-8
+ wkt2 = -2.0937989e-9
+ tpbsw = 0.0019
+ wmax = 8.9974e-6
+ aigc = 0.011522737
+ wmin = 8.974e-7
+ cjswd = 7.625999999999999e-11
+ aigbacc = 0.02
+ cjsws = 7.625999999999999e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ wua1 = 5.3887147e-17
+ wub1 = -8.2410881e-26
+ wuc1 = -2.4808749e-17
+ tpbswg = 0.0009
+ bigc = 0.001442
+ wwlc = 0
+ aigbinv = 0.0163
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.5522823e-12
+ cgdo = 5.2490134000000004e-11
+ xtid = 3
+ xtis = 3
+ ptvoff = 8.9623963e-17
+ ijthsfwd = 0.01
+ scref = 1e-6
+ cgsl = 3.5522823e-12
+ cgso = 5.2490134000000004e-11
+ cigc = 0.000625
+ waigsd = 3.0721194e-12
+ pigcd = 2.621
+ aigsd = 0.010772879
+ diomod = 1
+ lvoff = -4.3479245999999995e-10
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 2.6226e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.6226e-10
+ lvsat = -0.00019496033999999988
+ tvfbsdoff = 0.022
+ ijthsrev = 0.01
+ lvth0 = -8.10025498e-9
+ poxedge = 1
+ delta = 0.007595625
+ laigc = -4.6341008e-12
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ binunit = 2
+ rnoia = 0
+ rnoib = 0
+ mjswgd = 0.85
+ mjswgs = 0.85
+ k2we = 5e-5
+ pketa = -1.2207451e-14
+ tcjswg = 0.001
+ ngate = 8e+20
+ dsub = 0.75
+ ngcon = 1
+ dtox = 2.7e-10
+ wpclm = -2.3899735e-8
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ ppdiblc2 = 7.6111026e-16
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ eta0 = 0.3
+ etab = -0.24888148
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ fprout = 300
+ wtvfbsdoff = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ pkvth0we = -1.3e-19
+ ltvfbsdoff = 0
+ wtvoff = -8.2076521e-10
+ tvoff = 0.00074618122
+ vfbsdoff = 0.02
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ capmod = 2
+ njtsswg = 9
+ wku0we = 2e-11
+ paramchk = 1
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ ku0we = -0.0007
+ mobmod = 0
+ beta0 = 13
+ leta0 = 0
+ ckappad = 0.6
+ ptvfbsdoff = 0
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.022446923
+ pdiblcb = -0.3
+ ppclm = 9.2725546e-15
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ ijthdfwd = 0.01
+ keta = -0.10468292
+ bigbacc = 0.002588
+ laigsd = 3.9592657e-17
+ lags = 3.7696529e-13
+ dmcgt = 0
+ tcjsw = 0.000357
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 8.1265533e-11
+ kvth0we = 0.00018
+ ijthdrev = 0.01
+ kt1l = 0
+ lintnoi = -1.5e-8
+ lpdiblc2 = -1.4676946e-9
+ bigbinv = 0.004953
+ )

.model nch_ff_14 nmos (
+ level = 54
+ poxedge = 1
+ binunit = 2
+ scref = 1e-6
+ toxref = 3e-9
+ pigcd = 2.621
+ aigsd = 0.010772879
+ wags = 1.2013302e-6
+ lvoff = -2.0718068800000003e-9
+ pkvth0we = -1.3e-19
+ wcit = 1.2011066e-10
+ tvfbsdoff = 0.022
+ voff = -0.13980004150000003
+ lvsat = 0.0010644048900000005
+ lvth0 = 2.7772229100000004e-9
+ acde = 0.4
+ delta = 0.007595625
+ vsat = 89163.73610000002
+ laigc = -2.2637509e-11
+ wint = 0
+ vfbsdoff = 0.02
+ vth0 = 0.29349447529999995
+ ltvoff = 1.2509019e-10
+ wkt1 = 8.1830806e-8
+ wkt2 = 1.6147625e-8
+ rnoia = 0
+ rnoib = 0
+ wmax = 8.9974e-6
+ aigc = 0.011714263
+ wmin = 8.974e-7
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ pketa = 8.4378567e-15
+ ngate = 8e+20
+ paramchk = 1
+ ngcon = 1
+ wpclm = 3.4675908e-7
+ wua1 = -1.154179e-16
+ wub1 = 3.1505286e-27
+ wuc1 = 9.7519251e-17
+ lku0we = 2.5e-11
+ a0 = -0.035582299999999956
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ bigc = 0.001442
+ gbmin = 1e-12
+ epsrox = 3.9
+ at = 65883.509
+ cf = 8.720500000000001e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = -0.036587969000000005
+ k3 = -1.8419
+ wvfbsdoff = 0
+ em = 1000000.0
+ wwlc = 0
+ jswgd = 1.28e-13
+ lvfbsdoff = 0
+ jswgs = 1.28e-13
+ ll = 0
+ lw = 0
+ u0 = 0.007422836099999999
+ w0 = 0
+ ua = -2.421907e-9
+ ub = 1.9130826320999997e-18
+ uc = 4.338735e-12
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 2.33e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ rdsmod = 0
+ cdsc = 0
+ igbmod = 1
+ cgbo = 0
+ cgdl = 3.5522823e-12
+ cgdo = 5.2490134000000004e-11
+ xtid = 3
+ xtis = 3
+ ijthdfwd = 0.01
+ cgsl = 3.5522823e-12
+ cgso = 5.2490134000000004e-11
+ cigc = 0.000625
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ pbswgd = 0.95
+ pbswgs = 0.95
+ njtsswg = 9
+ igcmod = 1
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ ijthdrev = 0.01
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.006833075
+ pdiblcb = -0.3
+ tvoff = -0.00053245355
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ lpdiblc2 = 7.1362462e-15
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ k2we = 5e-5
+ paigsd = 1.5255572e-23
+ dsub = 0.75
+ dtox = 2.7e-10
+ ku0we = -0.0007
+ bigbacc = 0.002588
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ beta0 = 13
+ leta0 = 2.6128654e-9
+ letab = -2.2297043e-8
+ permod = 1
+ kvth0we = 0.00018
+ ppclm = -2.5569374e-14
+ eta0 = 0.27220356
+ etab = -0.011678893
+ lkvth0we = -2e-12
+ dlcig = 2.5e-9
+ lintnoi = -1.5e-8
+ bgidl = 2320000000.0
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ acnqsmod = 0
+ voffcv = -0.16942
+ wpemod = 1
+ dmcgt = 0
+ tcjsw = 0.000357
+ rbodymod = 0
+ bigsd = 0.00125
+ ags = 2.4574722
+ wvoff = 8.241506600000007e-9
+ cjd = 0.0012620099999999998
+ cit = 0.00079415993
+ cjs = 0.0012620099999999998
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 3.26497e-9
+ tpbswg = 0.0009
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ wvsat = -0.011322354899999998
+ nfactor = 1
+ wvth0 = -1.4059849099999998e-8
+ wpdiblc2 = 7.4309162e-10
+ waigc = -2.4473999e-12
+ la0 = 2.94419216e-8
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.0005899833300000001
+ kt1 = -0.41803712
+ lk2 = -5.0446112e-10
+ kt2 = -0.10268076
+ llc = 0
+ lln = 1
+ lu0 = 1.3321008000000002e-10
+ mjd = 0.26
+ lua = 3.6827721e-17
+ mjs = 0.26
+ lub = -1.9895881809999996e-26
+ luc = 1.827009e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ ptvoff = -1.5034232e-16
+ njd = 1.02
+ njs = 1.02
+ pa0 = 7.627786000000002e-15
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 9.5987885e-10
+ pbs = 0.52
+ pk2 = 1.6131306e-16
+ waigsd = 3.0714121e-12
+ lketa = 2.8547804e-8
+ pu0 = -1.7664274e-16
+ prt = 0
+ pua = -1.4490045e-23
+ xpart = 1
+ pub = 2.3973370000000036e-34
+ puc = 4.0045874e-24
+ pud = 0
+ rsh = 17.5
+ keta = -0.51555907
+ tcj = 0.00076
+ ua1 = 9.0255397e-10
+ ub1 = -8.0270486e-19
+ uc1 = -7.4218809e-11
+ diomod = 1
+ tpb = 0.0014
+ nigbacc = 10
+ wa0 = 1.203209e-7
+ egidl = 0.29734
+ ute = -1
+ wat = -0.011948694
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -5.5751276e-9
+ pditsd = 0
+ pditsl = 0
+ wlc = 0
+ wln = 1
+ wkvth0we = 2e-12
+ wu0 = 1.5300184999999998e-9
+ cjswgd = 2.6226e-10
+ pku0we = -1.5e-18
+ xgl = -1.09e-8
+ cjswgs = 2.6226e-10
+ xgw = 0
+ wua = 1.5882075e-16
+ wub = -5.862147e-26
+ wuc = -7.6599643e-17
+ wud = 0
+ wwc = 0
+ jswd = 1.28e-13
+ wwl = 0
+ wwn = 1
+ jsws = 1.28e-13
+ lcit = 1.0447464e-10
+ kt1l = 0
+ trnqsmod = 0
+ nigbinv = 10
+ lint = 0
+ mjswgd = 0.85
+ mjswgs = 0.85
+ lkt1 = 9.504028e-9
+ lkt2 = 1.0192413e-9
+ pvfbsdoff = 0
+ lmax = 9.167e-8
+ tcjswg = 0.001
+ lmin = 5.567e-8
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ minv = -0.3
+ rgatemod = 0
+ lua1 = -1.8750406e-17
+ wtvfbsdoff = 0
+ lub1 = -7.6940068e-27
+ luc1 = 1.062175e-17
+ pvoff = -1.135113399999999e-16
+ tnjtsswg = 1
+ fnoimod = 1
+ ndep = 1e+18
+ eigbinv = 1.1
+ cdscb = 0
+ cdscd = 0
+ lwlc = 0
+ moin = 5.1
+ pvsat = 7.102800199999998e-10
+ wk2we = 5e-12
+ pvth0 = -4.295049219999997e-16
+ ltvfbsdoff = 0
+ drout = 0.56
+ nigc = 3.083
+ paigc = 1.8938113e-18
+ fprout = 300
+ voffl = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ weta0 = -3.9858587e-8
+ wetab = 2.7041872e-8
+ lpclm = -8.5343289e-9
+ wtvoff = 1.7320676e-9
+ cigbacc = 0.32875
+ ntox = 2.029
+ pcit = -3.2574433e-17
+ pclm = 1.1824913
+ cgidl = 0.22
+ ptvfbsdoff = 0
+ tnoimod = 0
+ phin = 0.15
+ capmod = 2
+ pkt1 = -7.2665907e-15
+ pkt2 = -2.0869621e-15
+ wku0we = 2e-11
+ cigbinv = 0.006
+ pbswd = 0.8
+ pbsws = 0.8
+ mobmod = 0
+ rbdb = 50
+ pua1 = 1.2507395e-23
+ prwb = 0
+ prwg = 0
+ pub1 = -4.2778592e-33
+ puc1 = -7.7010123e-24
+ version = 4.5
+ pdits = 0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ cigsd = 0.069865
+ tempmod = 0
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ rdsw = 100
+ ijthsfwd = 0.01
+ aigbacc = 0.02
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ laigsd = -1.6939346e-18
+ tnoia = 0
+ ijthsrev = 0.01
+ rshg = 15.6
+ peta0 = 3.7467072e-15
+ aigbinv = 0.0163
+ petab = -3.4888335e-15
+ wketa = -1.1526014e-7
+ tpbsw = 0.0019
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ cjswd = 7.625999999999999e-11
+ cjsws = 7.625999999999999e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ ppdiblc2 = -4.5980291e-21
+ tnom = 25
+ toxe = 2.3900000000000002e-9
+ toxm = 2.43e-9
+ )

.model nch_ff_15 nmos (
+ level = 54
+ fnoimod = 1
+ ltvoff = -2.8596488e-10
+ eigbinv = 1.1
+ pvfbsdoff = 0
+ lku0we = 2.5e-11
+ epsrox = 3.9
+ pvoff = 8.85540199999999e-16
+ cdscb = 0
+ cdscd = 0
+ rdsmod = 0
+ cigbacc = 0.32875
+ pvsat = -2.6073073e-9
+ igbmod = 1
+ wk2we = 5e-12
+ pvth0 = -1.0527000000001127e-17
+ drout = 0.56
+ ijthsfwd = 0.01
+ paigc = 1.0773556e-18
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ tnoimod = 0
+ voffl = 0
+ pbswgd = 0.95
+ pbswgs = 0.95
+ keta = 0.067264197
+ cigbinv = 0.006
+ weta0 = 3.2678994e-7
+ igcmod = 1
+ wetab = -1.4667966e-7
+ lpclm = -8.0899178e-8
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 2.1355174e-10
+ ijthsrev = 0.01
+ kt1l = 0
+ cgidl = 0.22
+ version = 4.5
+ a0 = 5.6809619
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = -70591.59300000001
+ cf = 8.720500000000001e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = -0.016951152
+ k3 = -1.8419
+ em = 1000000.0
+ ll = 0
+ tempmod = 0
+ lw = 0
+ lint = 0
+ u0 = 0.00081555646
+ w0 = 0
+ ua = -3.0786989e-9
+ ub = 2.197681248e-18
+ uc = -5.08518e-12
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 2.33e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ lkt1 = -1.7073163e-8
+ lkt2 = 1.223943e-9
+ lmax = 5.567e-8
+ lmin = 4.667e-8
+ paigsd = -3.180948e-23
+ pbswd = 0.8
+ lpe0 = 9.2e-8
+ pbsws = 0.8
+ lpeb = 2.5e-7
+ aigbacc = 0.02
+ minv = -0.3
+ permod = 1
+ lua1 = 1.293984e-17
+ lub1 = 2.65765339e-26
+ luc1 = 1.702510023e-17
+ ndep = 1e+18
+ pdits = 0
+ lwlc = 0
+ cigsd = 0.069865
+ moin = 5.1
+ aigbinv = 0.0163
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ nigc = 3.083
+ voffcv = -0.16942
+ wpemod = 1
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ pkvth0we = -1.3e-19
+ tnoia = 0
+ ntox = 2.029
+ pcit = 1.39981203e-16
+ pclm = 2.4301611
+ peta0 = -1.7518907e-14
+ petab = 6.5870154e-15
+ vfbsdoff = 0.02
+ wketa = 1.9475197e-7
+ poxedge = 1
+ tpbsw = 0.0019
+ phin = 0.15
+ cjswd = 7.625999999999999e-11
+ cjsws = 7.625999999999999e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ binunit = 2
+ pkt1 = 1.2886179999999999e-14
+ pkt2 = 7.7933247e-16
+ tpbswg = 0.0009
+ paramchk = 1
+ rbdb = 50
+ pua1 = -3.7208869e-24
+ prwb = 0
+ prwg = 0
+ pub1 = -5.9613729e-32
+ puc1 = -1.1133321e-23
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ ptvoff = 3.472697e-16
+ waigsd = 3.0722235e-12
+ rdsw = 100
+ ijthdfwd = 0.01
+ scref = 1e-6
+ diomod = 1
+ pigcd = 2.621
+ aigsd = 0.010772879
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ pditsd = 0
+ pditsl = 0
+ lvoff = -3.7179500799999983e-9
+ cjswgd = 2.6226e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.6226e-10
+ tvfbsdoff = 0.022
+ lvsat = 0.0008510027900000004
+ ijthdrev = 0.01
+ lvth0 = 2.5627522400000005e-9
+ rshg = 15.6
+ delta = 0.007595625
+ laigc = -2.1310273e-11
+ wtvfbsdoff = 0
+ mjswgd = 0.85
+ mjswgs = 0.85
+ rnoia = 0
+ rnoib = 0
+ tcjswg = 0.001
+ ltvfbsdoff = 0
+ pketa = -9.5428465e-15
+ ngate = 8e+20
+ ngcon = 1
+ wpclm = -1.3405624e-6
+ njtsswg = 9
+ tnom = 25
+ wvfbsdoff = 0
+ gbmin = 1e-12
+ lvfbsdoff = 0
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ jswgd = 1.28e-13
+ toxe = 2.3900000000000002e-9
+ jswgs = 1.28e-13
+ toxm = 2.43e-9
+ ckappad = 0.6
+ lkvth0we = -2e-12
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.0068331981
+ pdiblcb = -0.3
+ fprout = 300
+ ptvfbsdoff = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ acnqsmod = 0
+ wags = 1.2013302e-6
+ wcit = -2.8549931e-9
+ wtvoff = -6.84745e-9
+ bigbacc = 0.002588
+ rbodymod = 0
+ voff = -0.111418263
+ acde = 0.4
+ vsat = 92843.10940000002
+ tvoff = 0.0065547027
+ kvth0we = 0.00018
+ wint = 0
+ vth0 = 0.297192242
+ wkt1 = -2.6563076e-7
+ wkt2 = -3.3271248e-8
+ xjbvd = 1
+ xjbvs = 1
+ wmax = 8.9974e-6
+ lk2we = -1.5e-12
+ capmod = 2
+ aigc = 0.011691379
+ wmin = 8.974e-7
+ lintnoi = -1.5e-8
+ bigbinv = 0.004953
+ wku0we = 2e-11
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ mobmod = 0
+ ku0we = -0.0007
+ wua1 = 1.6438006e-16
+ wub1 = 9.572171599999999e-25
+ wuc1 = 1.56696984e-16
+ beta0 = 13
+ wpdiblc2 = 7.4301235e-10
+ leta0 = 1.0110619e-10
+ letab = 3.9727723e-8
+ bigc = 0.001442
+ wwlc = 0
+ ppclm = 7.229527e-14
+ cdsc = 0
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ cgbo = 0
+ cgdl = 3.5522823e-12
+ cgdo = 5.2490134000000004e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.5522823e-12
+ cgso = 5.2490134000000004e-11
+ cigc = 0.000625
+ laigsd = 3.532034e-18
+ dmcgt = 0
+ wkvth0we = 2e-12
+ tcjsw = 0.000357
+ nfactor = 1
+ ags = 2.4574722
+ trnqsmod = 0
+ cjd = 0.0012620099999999998
+ cit = -0.0010864838
+ cjs = 0.0012620099999999998
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ dlc = 3.26497e-9
+ k3b = 1.9326
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ bigsd = 0.00125
+ k2we = 5e-5
+ wvoff = -8.983524000000003e-9
+ la0 = -3.0211764e-7
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = 0.0073255742000000006
+ dsub = 0.75
+ kt1 = 0.040190302
+ lk2 = -1.6433965e-9
+ kt2 = -0.1062101
+ dtox = 2.7e-10
+ llc = 0
+ lln = 1
+ lu0 = 5.1643238e-10
+ mjd = 0.26
+ nigbacc = 10
+ lua = 7.492165e-17
+ mjs = 0.26
+ lub = -3.6402602300000003e-26
+ luc = 2.373596e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ wvsat = 0.045877431999999996
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ njd = 1.02
+ njs = 1.02
+ pa0 = -1.230232e-13
+ rgatemod = 0
+ wvth0 = -2.1283431999999998e-8
+ nsd = 1e+20
+ pbd = 0.52
+ pat = -7.180893900000001e-9
+ pbs = 0.52
+ pk2 = 5.8185614e-16
+ tnjtsswg = 1
+ pu0 = -3.9034275e-17
+ prt = 0
+ pua = 3.4306982e-23
+ pub = -6.0757564e-32
+ puc = -7.1571349e-24
+ pud = 0
+ waigc = 1.1629424e-11
+ eta0 = 0.31550975
+ rsh = 17.5
+ etab = -1.0810714
+ tcj = 0.00076
+ ua1 = 3.5617042e-10
+ ub1 = -1.393576019e-18
+ uc1 = -1.8462139999999999e-10
+ tpb = 0.0014
+ wa0 = 2.372924e-6
+ ute = -1
+ wat = 0.12840945
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -1.282587e-8
+ nigbinv = 10
+ lketa = -5.2559457e-9
+ toxref = 3e-9
+ wlc = 0
+ wln = 1
+ wu0 = -8.425413540000001e-10
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -6.825073e-16
+ wub = 9.9305604e-25
+ wuc = 1.1584384e-16
+ wud = 0
+ wwc = 0
+ xpart = 1
+ wwl = 0
+ wwn = 1
+ egidl = 0.29734
+ )

.model nch_ff_16 nmos (
+ level = 54
+ pketa = 8.7750313e-15
+ pkt1 = -9.8484796e-16
+ pkt2 = 1.5926682e-15
+ ngate = 8e+20
+ lku0we = 2.5e-11
+ ngcon = 1
+ wpclm = -1.03603352e-6
+ epsrox = 3.9
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ wpdiblc2 = 7.4301235e-10
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ rdsmod = 0
+ bigbacc = 0.002588
+ rbdb = 50
+ pua1 = -1.9060214e-23
+ prwb = 0
+ prwg = 0
+ pub1 = 2.6550731000000005e-32
+ puc1 = 1.47310838e-23
+ igbmod = 1
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ rdsw = 100
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ kvth0we = 0.00018
+ pbswgd = 0.95
+ pbswgs = 0.95
+ lintnoi = -1.5e-8
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ igcmod = 1
+ wkvth0we = 2e-12
+ rshg = 15.6
+ trnqsmod = 0
+ tvoff = 0.002919136
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ paigsd = 4.3875156e-23
+ ku0we = -0.0007
+ permod = 1
+ beta0 = 13
+ rgatemod = 0
+ leta0 = 1.5743207e-8
+ tnom = 25
+ letab = 3.0329695e-8
+ tnjtsswg = 1
+ toxe = 2.3900000000000002e-9
+ toxm = 2.43e-9
+ nfactor = 1
+ ppclm = 5.7373356e-14
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ voffcv = -0.16942
+ wpemod = 1
+ a0 = 3.2177147
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 97840.91
+ cf = 8.720500000000001e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.023015951
+ k3 = -1.8419
+ em = 1000000.0
+ ll = 0
+ lw = 0
+ ags = 2.4574722
+ u0 = 0.0036279722999999994
+ w0 = 0
+ ua = -2.19661343e-9
+ ub = 1.4860819409999996e-18
+ uc = 2.2595638e-10
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ wags = 1.2013302e-6
+ xl = 2.33e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ cjd = 0.0012620099999999998
+ cit = -0.0084826049
+ cjs = 0.0012620099999999998
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dmcgt = 0
+ dlc = 3.26497e-9
+ wcit = 1.1098639999999993e-10
+ tcjsw = 0.000357
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ nigbacc = 10
+ voff = -0.04075972859999999
+ acde = 0.4
+ la0 = -1.8141853e-7
+ vsat = 64987.781699999985
+ wint = 0
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.0009276249
+ vth0 = 0.37735216059999993
+ kt1 = -0.20813859
+ lk2 = -3.6017846e-9
+ kt2 = -0.11042259
+ llc = 0
+ lln = 1
+ lu0 = 3.7862393e-10
+ wkt1 = 1.7451446e-8
+ wkt2 = -4.9869936e-8
+ mjd = 0.26
+ bigsd = 0.00125
+ lua = 3.1699464000000005e-17
+ mjs = 0.26
+ lub = -1.5342368999999952e-27
+ luc = -8.94744e-18
+ lud = 0
+ wmax = 8.9974e-6
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ aigc = 0.011397597
+ wmin = 8.974e-7
+ njs = 1.02
+ pa0 = -1.9996651e-13
+ nsd = 1e+20
+ nigbinv = 10
+ pbd = 0.52
+ pat = -9.658699e-10
+ pbs = 0.52
+ pk2 = 3.3250012e-16
+ tpbswg = 0.0009
+ pu0 = -3.9242668999999997e-17
+ prt = 0
+ pua = 2.7971342e-23
+ pub = -4.5926045000000006e-32
+ puc = -7.6781524e-24
+ pud = 0
+ wvoff = 8.333983999999995e-9
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 4.3071269e-10
+ ub1 = -7.468433610000001e-19
+ uc1 = 5.294111900000001e-10
+ wua1 = 4.7742754e-16
+ tpb = 0.0014
+ wub1 = -8.0124139e-25
+ wuc1 = -3.71148e-16
+ wvsat = 0.037473207999999994
+ wa0 = 3.9431957e-6
+ wvth0 = -5.0348026999999994e-8
+ ute = -1
+ wat = 0.0015722129999999994
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -7.7369724e-9
+ bigc = 0.001442
+ wlc = 0
+ wln = 1
+ wu0 = -8.3828936e-10
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -5.5320853e-16
+ wub = 6.903720200000001e-25
+ wuc = 1.2647685e-16
+ wud = 0
+ wwlc = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ waigc = -9.3979847e-11
+ ptvoff = -3.4317401e-17
+ waigsd = 3.0706789e-12
+ fnoimod = 1
+ cdsc = 0
+ eigbinv = 1.1
+ cgbo = 0
+ cgdl = 3.5522823e-12
+ cgdo = 5.2490134000000004e-11
+ xtid = 3
+ lketa = -2.4929909e-8
+ xtis = 3
+ ijthsfwd = 0.01
+ diomod = 1
+ cgsl = 3.5522823e-12
+ cgso = 5.2490134000000004e-11
+ xpart = 1
+ wtvfbsdoff = 0
+ cigc = 0.000625
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 2.6226e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.6226e-10
+ egidl = 0.29734
+ ltvfbsdoff = 0
+ ijthsrev = 0.01
+ mjswgd = 0.85
+ mjswgs = 0.85
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ cigbacc = 0.32875
+ pvfbsdoff = 0
+ tcjswg = 0.001
+ tnoimod = 0
+ k2we = 5e-5
+ dsub = 0.75
+ dtox = 2.7e-10
+ ptvfbsdoff = 0
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ cigbinv = 0.006
+ pvoff = 3.698261999999959e-17
+ cdscb = 0
+ cdscd = 0
+ eta0 = -0.003716791
+ etab = -0.88927493
+ pvsat = -2.1955010499999996e-9
+ wk2we = 5e-12
+ pvth0 = 1.41363016e-15
+ drout = 0.56
+ version = 4.5
+ fprout = 300
+ paigc = 6.2522098e-18
+ tempmod = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ voffl = 0
+ weta0 = 2.2378028e-8
+ pkvth0we = -1.3e-19
+ wetab = 3.831648e-8
+ aigbacc = 0.02
+ wtvoff = 9.4004181e-10
+ lpclm = -7.043921000000001e-8
+ cgidl = 0.22
+ vfbsdoff = 0.02
+ capmod = 2
+ aigbinv = 0.0163
+ wku0we = 2e-11
+ mobmod = 0
+ pbswd = 0.8
+ pbsws = 0.8
+ paramchk = 1
+ pdits = 0
+ cigsd = 0.069865
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ poxedge = 1
+ ijthdfwd = 0.01
+ laigsd = -2.6649547e-17
+ pk2we = -1e-19
+ keta = 0.46877367
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ binunit = 2
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ tnoia = 0
+ lcit = 5.7596243e-10
+ ijthdrev = 0.01
+ kt1l = 0
+ peta0 = -2.6027237e-15
+ petab = -2.4777955e-15
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ wketa = -1.7908228e-7
+ tpbsw = 0.0019
+ lint = 0
+ cjswd = 7.625999999999999e-11
+ cjsws = 7.625999999999999e-11
+ lkt1 = -4.905047e-9
+ lkt2 = 1.4303548e-9
+ mjswd = 0.11
+ lmax = 4.667e-8
+ mjsws = 0.11
+ agidl = 9.41e-8
+ lmin = 3.6e-8
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ minv = -0.3
+ lua1 = 9.2872684e-18
+ lub1 = -5.113301800000003e-27
+ luc1 = -1.796249619e-17
+ ndep = 1e+18
+ lwlc = 0
+ lkvth0we = -2e-12
+ moin = 5.1
+ toxref = 3e-9
+ nigc = 3.083
+ scref = 1e-6
+ pigcd = 2.621
+ aigsd = 0.01077288
+ acnqsmod = 0
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ lvoff = -7.180218279999999e-9
+ tvfbsdoff = 0.022
+ njtsswg = 9
+ rbodymod = 0
+ lvsat = 0.002215917613
+ lvth0 = -1.3650739699999994e-9
+ ntox = 2.029
+ ltvoff = -1.0782211e-10
+ pcit = -5.351009999999994e-18
+ pclm = 2.21669238
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ delta = 0.007595625
+ laigc = -6.9149623e-12
+ ckappad = 0.6
+ ckappas = 0.6
+ rnoia = 0
+ rnoib = 0
+ pdiblc1 = 0
+ pdiblc2 = 0.0068331981
+ phin = 0.15
+ pdiblcb = -0.3
+ )

.model nch_ff_17 nmos (
+ level = 54
+ cgbo = 0
+ cgdl = 3.5522823e-12
+ cgdo = 5.2490134000000004e-11
+ xtid = 3
+ pbswgd = 0.95
+ xtis = 3
+ pbswgs = 0.95
+ ijthdfwd = 0.01
+ cgsl = 3.5522823e-12
+ cgso = 5.2490134000000004e-11
+ aigbinv = 0.0163
+ cigc = 0.000625
+ voffl = 0
+ igcmod = 1
+ weta0 = -1.09928e-7
+ wetab = 2.7482e-8
+ ijthdrev = 0.01
+ cgidl = 0.22
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ poxedge = 1
+ k2we = 5e-5
+ pbswd = 0.8
+ pbsws = 0.8
+ dsub = 0.75
+ permod = 1
+ dtox = 2.7e-10
+ binunit = 2
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ pdits = 0
+ eta0 = 0.42133333
+ cigsd = 0.069865
+ etab = -0.29033333
+ lkvth0we = -2e-12
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ voffcv = -0.16942
+ wpemod = 1
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ acnqsmod = 0
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ tnoia = 0
+ rbodymod = 0
+ peta0 = 0
+ wketa = -3.7974654e-8
+ tpbsw = 0.0019
+ cjswd = 7.625999999999999e-11
+ tpbswg = 0.0009
+ cjsws = 7.625999999999999e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ wtvfbsdoff = 0
+ a0 = 2.2098167
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 72000
+ cf = 8.720500000000001e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.014686228
+ k3 = -1.8419
+ em = 1000000.0
+ wpdiblc2 = -6.449088e-9
+ ll = 0
+ lw = 0
+ u0 = 0.0151465
+ w0 = 0
+ ua = -1.7855187e-9
+ ub = 2.0636167e-18
+ uc = 7.8391667e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 2.33e-9
+ ptvoff = 0
+ ww = 0
+ xw = 8.600000000000001e-9
+ njtsswg = 9
+ ltvfbsdoff = 0
+ waigsd = 3.0876027e-12
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ diomod = 1
+ scref = 1e-6
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.025656394
+ pigcd = 2.621
+ pdiblcb = -0.3
+ pditsd = 0
+ pditsl = 0
+ aigsd = 0.010772862
+ cjswgd = 2.6226e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.6226e-10
+ keta = 0.015093331
+ tvfbsdoff = 0.022
+ lvoff = -2e-11
+ wkvth0we = 2e-12
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lvsat = -0.0003
+ lcit = -1e-11
+ lvth0 = -1e-10
+ ptvfbsdoff = 0
+ kt1l = 0
+ mjswgd = 0.85
+ mjswgs = 0.85
+ trnqsmod = 0
+ delta = 0.007595625
+ bigbacc = 0.002588
+ tcjswg = 0.001
+ rnoia = 0
+ rnoib = 0
+ lint = 6.5375218e-9
+ kvth0we = 0.00018
+ lkt1 = -1.1e-9
+ lmax = 2.001e-5
+ lmin = 9.00077e-6
+ ngate = 8e+20
+ lintnoi = -1.5e-8
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ ngcon = 1
+ bigbinv = 0.004953
+ wpclm = 5.7423639e-7
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ rgatemod = 0
+ minv = -0.3
+ lub1 = 0
+ gbmin = 1e-12
+ tnjtsswg = 1
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ ndep = 1e+18
+ lwlc = 0
+ moin = 5.1
+ fprout = 300
+ nigc = 3.083
+ xrcrg1 = 12
+ xrcrg2 = 1
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ wtvoff = 9.3503662e-10
+ ntox = 2.029
+ pcit = -1.5e-17
+ pclm = 0.629885
+ tvoff = 5.0359625e-5
+ capmod = 2
+ nfactor = 1
+ wku0we = 2e-11
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ phin = 0.15
+ mobmod = 0
+ pkt1 = -5e-17
+ ku0we = -0.0007
+ beta0 = 13
+ leta0 = 0
+ nigbacc = 10
+ rbdb = 50
+ prwb = 0
+ prwg = 0
+ pub1 = 0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ ags = 0.58720097
+ dlcig = 2.5e-9
+ rdsw = 100
+ bgidl = 2320000000.0
+ cjd = 0.0012620099999999998
+ cit = 6.2896875e-5
+ cjs = 0.0012620099999999998
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 9.8024918e-9
+ ijthsfwd = 0.01
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ nigbinv = 10
+ la0 = 0
+ jsd = 6.11e-7
+ dmcgt = 0
+ jss = 6.11e-7
+ lat = -0.0001
+ kt1 = -0.28314411
+ kt2 = -0.074391698
+ tcjsw = 0.000357
+ llc = 0
+ lln = 1
+ lu0 = 6e-12
+ mjd = 0.26
+ mjs = 0.26
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 0
+ ijthsrev = 0.01
+ nsd = 1e+20
+ pbd = 0.52
+ pat = -2.8e-11
+ pbs = 0.52
+ rshg = 15.6
+ pu0 = 2e-18
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ prt = 0
+ pud = 0
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = -6.8749055e-10
+ ub1 = 1.0341951e-18
+ uc1 = 4.5339833e-11
+ fnoimod = 1
+ bigsd = 0.00125
+ tpb = 0.0014
+ wa0 = 7.159061e-7
+ eigbinv = 1.1
+ ute = -2.01925
+ wat = 0
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 3.760485e-9
+ wlc = 0
+ wln = 1
+ wu0 = -1.59669e-10
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -7.132277e-17
+ wub = 7.28273e-26
+ wuc = -1.167985e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ wvoff = 1.0181215e-9
+ wvsat = -0.0045771271
+ wvth0 = -1.27727395e-8
+ tnom = 25
+ toxe = 2.3900000000000002e-9
+ waigc = 5.0140497e-11
+ toxm = 2.43e-9
+ toxref = 3e-9
+ cigbacc = 0.32875
+ xpart = 1
+ tnoimod = 0
+ wags = 9.993247e-8
+ egidl = 0.29734
+ pkvth0we = -1.3e-19
+ wcit = 4.9907306e-10
+ cigbinv = 0.006
+ voff = -0.11158375
+ ltvoff = 0
+ acde = 0.4
+ vsat = 106133.02
+ vfbsdoff = 0.02
+ wint = 0
+ pvfbsdoff = 0
+ vth0 = 0.31972953
+ wkt1 = 3.2075481e-8
+ wkt2 = 1.5939759e-8
+ wmax = 8.974e-7
+ aigc = 0.011740211
+ wmin = 5.374e-7
+ version = 4.5
+ tempmod = 0
+ lku0we = 2.5e-11
+ epsrox = 3.9
+ paramchk = 1
+ wua1 = 1.0731531e-15
+ wub1 = -9.2968455e-25
+ wuc1 = -1.4414309e-17
+ aigbacc = 0.02
+ rdsmod = 0
+ bigc = 0.001442
+ pvoff = 0
+ wute = 5.565105e-7
+ wwlc = 0
+ igbmod = 1
+ cdscb = 0
+ cdscd = 0
+ pvsat = -1.8e-11
+ wk2we = 5e-12
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ pvth0 = -2.3e-16
+ cdsc = 0
+ drout = 0.56
+ )

.model nch_ff_18 nmos (
+ level = 54
+ kt1l = 0
+ nigbacc = 10
+ tvoff = -0.0002433276
+ paigsd = 1.3573222e-22
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ lint = 6.5375218e-9
+ lkt1 = 8.5146405e-8
+ lkt2 = 5.1456509e-9
+ lmax = 9.00077e-6
+ lmin = 9.0075e-7
+ permod = 1
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ nigbinv = 10
+ ags = 0.5416128899999999
+ ku0we = -0.0007
+ ppdiblc2 = 1.9760389e-14
+ beta0 = 13
+ cjd = 0.0012620099999999998
+ leta0 = 0
+ cit = -0.00011782923
+ cjs = 0.0012620099999999998
+ minv = -0.3
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ lua1 = 1.38467e-15
+ lub1 = -1.4892591e-24
+ luc1 = 1.0686128e-16
+ dlc = 9.8024918e-9
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ ndep = 1e+18
+ lute = 1.0068051e-6
+ lwlc = 0
+ moin = 5.1
+ dlcig = 2.5e-9
+ voffcv = -0.16942
+ wpemod = 1
+ bgidl = 2320000000.0
+ la0 = -1.1479603e-6
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ nigc = 3.083
+ lat = 0.085245067
+ kt1 = -0.2927377
+ lk2 = -1.3507419e-8
+ kt2 = -0.074964073
+ llc = 0
+ lln = 1
+ lu0 = -1.9944396e-9
+ fnoimod = 1
+ mjd = 0.26
+ lua = -1.5028094e-16
+ mjs = 0.26
+ lub = -1.4426347e-25
+ luc = -5.2935673e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = -5.1713984e-13
+ eigbinv = 1.1
+ nsd = 1e+20
+ pbd = 0.52
+ pat = -2.8e-11
+ pbs = 0.52
+ pk2 = -1.6553107e-15
+ pu0 = 1.5573224e-17
+ prt = 0
+ noff = 2.7195
+ pua = -3.5916841e-23
+ pub = 6.5823852e-32
+ puc = 3.1761344e-23
+ pud = 0
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ pkvth0we = -1.3e-19
+ dmcgt = 0
+ rsh = 17.5
+ tcjsw = 0.000357
+ tcj = 0.00076
+ ua1 = -8.4151391e-10
+ ub1 = 1.1998524e-18
+ uc1 = 3.3453151e-11
+ tpb = 0.0014
+ wa0 = 7.7343e-7
+ pags = -1.4569295e-13
+ ute = -2.1312417
+ wtvfbsdoff = 0
+ wat = 0
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 3.944613e-9
+ wlc = 0
+ wln = 1
+ ntox = 2.029
+ wu0 = -1.6117881e-10
+ pcit = -6.4447523e-16
+ xgl = -1.09e-8
+ pclm = 0.629885
+ xgw = 0
+ wua = -6.7327571e-17
+ wub = 6.5505403e-26
+ wuc = -1.5212814e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ vfbsdoff = 0.02
+ tpbswg = 0.0009
+ bigsd = 0.00125
+ ltvfbsdoff = 0
+ phin = 0.15
+ cigbacc = 0.32875
+ wvoff = 8.2208115e-10
+ pkt1 = -6.957314e-14
+ pkt2 = -1.5079533e-14
+ paramchk = 1
+ tnoimod = 0
+ wvsat = -0.0045771271
+ wvth0 = -1.3076090100000001e-8
+ ptvoff = -2.0299898e-15
+ waigsd = 3.0875876e-12
+ waigc = 5.030718e-11
+ rbdb = 50
+ pua1 = -1.044071e-21
+ prwb = 0
+ prwg = 0
+ pub1 = 9.8799081e-31
+ cigbinv = 0.006
+ puc1 = -4.3746501e-23
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ pute = -5.4971558e-13
+ diomod = 1
+ rdsw = 100
+ ptvfbsdoff = 0
+ lketa = -1.3350472e-7
+ ijthdfwd = 0.01
+ pditsd = 0
+ xpart = 1
+ pditsl = 0
+ cjswgd = 2.6226e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.6226e-10
+ version = 4.5
+ tempmod = 0
+ egidl = 0.29734
+ mjswgd = 0.85
+ mjswgs = 0.85
+ ijthdrev = 0.01
+ aigbacc = 0.02
+ a0 = 2.3375097
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ rshg = 15.6
+ at = 62506.667
+ cf = 8.720500000000001e-11
+ tcjswg = 0.001
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.016188722000000003
+ k3 = -1.8419
+ em = 1000000.0
+ pvfbsdoff = 0
+ ll = 0
+ lw = 0
+ u0 = 0.015369018
+ lpdiblc2 = -2.2119558e-8
+ w0 = 0
+ ua = -1.7688022e-9
+ ub = 2.0796638e-18
+ uc = 8.4279951e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 2.33e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ aigbinv = 0.0163
+ tnom = 25
+ pvoff = 1.7624031e-15
+ toxe = 2.3900000000000002e-9
+ toxm = 2.43e-9
+ cdscb = 0
+ cdscd = 0
+ fprout = 300
+ pvsat = -1.8e-11
+ lkvth0we = -2e-12
+ wk2we = 5e-12
+ pvth0 = 2.4971227e-15
+ drout = 0.56
+ xrcrg1 = 12
+ xrcrg2 = 1
+ paigc = -1.4984839e-18
+ voffl = 0
+ poxedge = 1
+ acnqsmod = 0
+ wtvoff = 1.1608419e-9
+ wags = 1.1613858999999999e-7
+ weta0 = -1.09928e-7
+ wetab = 2.7482e-8
+ wcit = 5.6909255e-10
+ binunit = 2
+ rbodymod = 0
+ voff = -0.1094379
+ acde = 0.4
+ capmod = 2
+ cgidl = 0.22
+ vsat = 106133.02
+ wint = 0
+ wku0we = 2e-11
+ vth0 = 0.31394058999999996
+ wkt1 = 3.9808867e-8
+ wkt2 = 1.7617127e-8
+ wmax = 8.974e-7
+ mobmod = 0
+ aigc = 0.011757817
+ wmin = 5.374e-7
+ pbswd = 0.8
+ pbsws = 0.8
+ wua1 = 1.1892901e-15
+ wub1 = -1.0395834e-24
+ wuc1 = -9.5481798e-18
+ wpdiblc2 = -8.647129e-9
+ bigc = 0.001442
+ wute = 6.1765795e-7
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ wwlc = 0
+ pdits = 0
+ cigsd = 0.069865
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ laigsd = -2.4859383e-16
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.5522823e-12
+ cgdo = 5.2490134000000004e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.5522823e-12
+ cgso = 5.2490134000000004e-11
+ cigc = 0.000625
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ wkvth0we = 2e-12
+ tnoia = 0
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ trnqsmod = 0
+ peta0 = 0
+ njtsswg = 9
+ wketa = -4.7550208e-8
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ tpbsw = 0.0019
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ cjswd = 7.625999999999999e-11
+ cjsws = 7.625999999999999e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.028116857
+ k2we = 5e-5
+ pdiblcb = -0.3
+ dsub = 0.75
+ dtox = 2.7e-10
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ rgatemod = 0
+ tnjtsswg = 1
+ toxref = 3e-9
+ eta0 = 0.42133333
+ etab = -0.29033333
+ bigbacc = 0.002588
+ scref = 1e-6
+ pigcd = 2.621
+ aigsd = 0.010772862
+ kvth0we = 0.00018
+ tvfbsdoff = 0.022
+ lvoff = -1.9311251e-8
+ lintnoi = -1.5e-8
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ ltvoff = 2.6402481e-9
+ lvsat = -0.0003
+ lvth0 = 5.1942566e-8
+ delta = 0.007595625
+ laigc = -1.5827875e-10
+ rnoia = 0
+ rnoib = 0
+ lku0we = 2.5e-11
+ pketa = 8.6084224e-14
+ epsrox = 3.9
+ ngate = 8e+20
+ ngcon = 1
+ wvfbsdoff = 0
+ wpclm = 5.7423639e-7
+ lvfbsdoff = 0
+ rdsmod = 0
+ gbmin = 1e-12
+ igbmod = 1
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ pbswgd = 0.95
+ pbswgs = 0.95
+ nfactor = 1
+ ijthsfwd = 0.01
+ igcmod = 1
+ keta = 0.029943688
+ lags = 4.0983681e-7
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 1.6147277e-9
+ ijthsrev = 0.01
+ )

.model nch_ff_19 nmos (
+ level = 54
+ rgatemod = 0
+ tnom = 25
+ tnjtsswg = 1
+ toxe = 2.3900000000000002e-9
+ toxm = 2.43e-9
+ pdits = 0
+ cigsd = 0.069865
+ voffcv = -0.16942
+ wpemod = 1
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ njtsswg = 9
+ wtvfbsdoff = 0
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ ltvfbsdoff = 0
+ ckappad = 0.6
+ ckappas = 0.6
+ wags = -7.98542e-7
+ pdiblc1 = 0
+ pdiblc2 = -0.019237439
+ pdiblcb = -0.3
+ wcit = -4.0548514e-10
+ tnoia = 0
+ voff = -0.12566406
+ acde = 0.4
+ peta0 = 0
+ vsat = 106133.02
+ wketa = 9.2259042e-8
+ wint = 0
+ tpbswg = 0.0009
+ vth0 = 0.37214179
+ tpbsw = 0.0019
+ wkt1 = -7.1953249e-8
+ wkt2 = 3.7202325e-9
+ wmax = 8.974e-7
+ bigbacc = 0.002588
+ cjswd = 7.625999999999999e-11
+ aigc = 0.01160027
+ cjsws = 7.625999999999999e-11
+ wmin = 5.374e-7
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ ptvfbsdoff = 0
+ kvth0we = 0.00018
+ ptvoff = 9.96032e-16
+ wua1 = 1.1798319e-17
+ wub1 = 1.8760115e-25
+ wuc1 = -8.2926019e-17
+ lintnoi = -1.5e-8
+ waigsd = 3.0878745e-12
+ bigbinv = 0.004953
+ bigc = 0.001442
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ wwlc = 0
+ diomod = 1
+ cdsc = 0
+ cgbo = 0
+ pditsd = 0
+ pditsl = 0
+ cgdl = 3.5522823e-12
+ cgdo = 5.2490134000000004e-11
+ xtid = 3
+ xtis = 3
+ cjswgd = 2.6226e-10
+ ijthsfwd = 0.01
+ scref = 1e-6
+ pku0we = -1.5e-18
+ cjswgs = 2.6226e-10
+ cgsl = 3.5522823e-12
+ cgso = 5.2490134000000004e-11
+ cigc = 0.000625
+ pigcd = 2.621
+ tvfbsdoff = 0.022
+ aigsd = 0.010772861
+ lvoff = -4.8699703e-9
+ mjswgd = 0.85
+ mjswgs = 0.85
+ lvsat = -0.0003
+ lvth0 = 1.4349239999999998e-10
+ ijthsrev = 0.01
+ tcjswg = 0.001
+ delta = 0.007595625
+ laigc = -1.8062176e-11
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ rnoia = 0
+ rnoib = 0
+ nfactor = 1
+ pketa = -3.8346008e-14
+ ngate = 8e+20
+ k2we = 5e-5
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ ngcon = 1
+ dsub = 0.75
+ wpclm = 5.7423639e-7
+ dtox = 2.7e-10
+ ppdiblc2 = -1.3176269e-14
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ fprout = 300
+ eta0 = 0.42133333
+ etab = -0.29033333
+ xrcrg1 = 12
+ xrcrg2 = 1
+ nigbacc = 10
+ a0 = 1.6362276
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 209176.65
+ cf = 8.720500000000001e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.012938798
+ k3 = -1.8419
+ em = 1000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.014847274
+ w0 = 0
+ ua = -1.7708735e-9
+ ub = 1.8600147e-18
+ uc = 2.580063e-11
+ ud = 0
+ wtvoff = -2.2391826e-9
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 2.33e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ pkvth0we = -1.3e-19
+ nigbinv = 10
+ capmod = 2
+ wku0we = 2e-11
+ tvoff = 0.004406442
+ vfbsdoff = 0.02
+ mobmod = 0
+ ags = 2.4075610000000003
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ cjd = 0.0012620099999999998
+ cit = 0.0020125208
+ cjs = 0.0012620099999999998
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 9.8024918e-9
+ k3b = 1.9326
+ fnoimod = 1
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ eigbinv = 1.1
+ paramchk = 1
+ ku0we = -0.0007
+ beta0 = 13
+ la0 = -5.2381924e-7
+ leta0 = 0
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.04529122
+ kt1 = -0.12585017
+ lk2 = -1.0614987e-8
+ kt2 = -0.061139846
+ llc = 0
+ lln = 1
+ lu0 = -1.5300873e-9
+ mjd = 0.26
+ lua = -1.4843753e-16
+ mjs = 0.26
+ lub = 5.1224193e-26
+ luc = -8.8907704e-19
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 9.5948774e-14
+ nsd = 1e+20
+ pbd = 0.52
+ pat = -5.002413e-9
+ pbs = 0.52
+ laigsd = 2.1900591e-16
+ pk2 = -1.0578878e-15
+ pu0 = 1.3957723999999998e-17
+ dlcig = 2.5e-9
+ prt = 0
+ pua = 5.0063903e-23
+ pub = -8.0709098e-32
+ puc = -9.2074471e-24
+ pud = 0
+ bgidl = 2320000000.0
+ ijthdfwd = 0.01
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 7.2552224e-10
+ ub1 = -4.8701436e-19
+ uc1 = 1.8003493e-10
+ tpb = 0.0014
+ wa0 = 8.4566389e-8
+ ute = -1
+ wat = 0.0055892281
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 3.2733514e-9
+ keta = -0.17327473
+ cigbacc = 0.32875
+ wlc = 0
+ wln = 1
+ wu0 = -1.5936364000000001e-10
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -1.6393515e-16
+ wub = 2.3014917e-25
+ wuc = 3.0819536e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ dmcgt = 0
+ tcjsw = 0.000357
+ lags = -1.250857e-6
+ tnoimod = 0
+ jswd = 1.28e-13
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ jsws = 1.28e-13
+ lcit = -2.812838e-10
+ ijthdrev = 0.01
+ kt1l = 0
+ cigbinv = 0.006
+ lpdiblc2 = 2.0025765e-8
+ bigsd = 0.00125
+ lint = 6.5375218e-9
+ lkt1 = -6.3383496e-8
+ lkt2 = -7.1579117e-9
+ lmax = 9.0075e-7
+ lmin = 4.5075e-7
+ wvoff = 5.2999378e-9
+ lpe0 = 9.2e-8
+ version = 4.5
+ lpeb = 2.5e-7
+ tempmod = 0
+ wvsat = -0.0045771271
+ wvth0 = -1.15199227e-8
+ minv = -0.3
+ lua1 = -9.9922063e-18
+ lub1 = 1.2052288e-26
+ luc1 = -2.3596511e-17
+ toxref = 3e-9
+ waigc = 6.3350032e-11
+ ndep = 1e+18
+ aigbacc = 0.02
+ lwlc = 0
+ lkvth0we = -2e-12
+ moin = 5.1
+ lketa = 4.735968e-8
+ nigc = 3.083
+ xpart = 1
+ acnqsmod = 0
+ aigbinv = 0.0163
+ egidl = 0.29734
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ ltvoff = -1.4980468e-9
+ rbodymod = 0
+ pags = 6.6837277e-13
+ ntox = 2.029
+ pvfbsdoff = 0
+ pcit = 2.2289891e-16
+ pclm = 0.629885
+ phin = 0.15
+ lku0we = 2.5e-11
+ epsrox = 3.9
+ pkt1 = 2.9895144e-14
+ pkt2 = -2.7112972e-15
+ poxedge = 1
+ rdsmod = 0
+ igbmod = 1
+ wpdiblc2 = 2.8360352e-8
+ pvoff = -2.2228894e-15
+ binunit = 2
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ rbdb = 50
+ pua1 = 3.8966634e-24
+ prwb = 0
+ prwg = 0
+ pub1 = -1.0420346e-31
+ cdscb = 0
+ cdscd = 0
+ puc1 = 2.1559776e-23
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ pvsat = -1.8e-11
+ rbsb = 50
+ pvag = 1.2
+ pbswgd = 0.95
+ pbswgs = 0.95
+ wk2we = 5e-12
+ pvth0 = 1.1121337e-15
+ drout = 0.56
+ rdsw = 100
+ igcmod = 1
+ paigc = -1.3106622e-17
+ voffl = 0
+ weta0 = -1.09928e-7
+ wetab = 2.7482e-8
+ wkvth0we = 2e-12
+ trnqsmod = 0
+ cgidl = 0.22
+ rshg = 15.6
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ paigsd = -1.1957726e-22
+ permod = 1
+ pbswd = 0.8
+ pbsws = 0.8
+ )

.model nch_ff_20 nmos (
+ level = 54
+ rgatemod = 0
+ tnom = 25
+ tnjtsswg = 1
+ toxe = 2.3900000000000002e-9
+ toxm = 2.43e-9
+ pdits = 0
+ cigsd = 0.069865
+ voffcv = -0.16942
+ wpemod = 1
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ njtsswg = 9
+ wtvfbsdoff = 0
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ ltvfbsdoff = 0
+ ckappad = 0.6
+ ckappas = 0.6
+ wags = 2.499663e-6
+ pdiblc1 = 0
+ pdiblc2 = 0.041730695
+ pdiblcb = -0.3
+ wcit = 2.0646633e-10
+ tnoia = 0
+ voff = -0.11119538
+ acde = 0.4
+ peta0 = 0
+ vsat = 99029.765
+ wketa = 8.4379468e-9
+ wint = 0
+ tpbswg = 0.0009
+ vth0 = 0.38049988999999995
+ tpbsw = 0.0019
+ wkt1 = 8.316763e-9
+ wkt2 = -6.4493333e-9
+ wmax = 8.974e-7
+ bigbacc = 0.002588
+ cjswd = 7.625999999999999e-11
+ aigc = 0.011620363
+ cjsws = 7.625999999999999e-11
+ wmin = 5.374e-7
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ ptvfbsdoff = 0
+ kvth0we = 0.00018
+ ptvoff = -1.0913215e-16
+ wua1 = 2.6150731e-17
+ wub1 = -7.4432483e-26
+ wuc1 = -3.5091334e-17
+ lintnoi = -1.5e-8
+ waigsd = 3.0877293e-12
+ bigbinv = 0.004953
+ bigc = 0.001442
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ wwlc = 0
+ diomod = 1
+ cdsc = 0
+ cgbo = 0
+ pditsd = 0
+ pditsl = 0
+ cgdl = 3.5522823e-12
+ cgdo = 5.2490134000000004e-11
+ xtid = 3
+ xtis = 3
+ cjswgd = 2.6226e-10
+ ijthsfwd = 0.01
+ scref = 1e-6
+ pku0we = -1.5e-18
+ cjswgs = 2.6226e-10
+ cgsl = 3.5522823e-12
+ cgso = 5.2490134000000004e-11
+ cigc = 0.000625
+ pigcd = 2.621
+ tvfbsdoff = 0.022
+ aigsd = 0.010772861
+ lvoff = -1.123619e-8
+ mjswgd = 0.85
+ mjswgs = 0.85
+ lvsat = 0.0028254309
+ lvth0 = -3.534068e-9
+ ijthsrev = 0.01
+ tcjswg = 0.001
+ delta = 0.007595625
+ laigc = -2.6902885e-11
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ rnoia = 0
+ rnoib = 0
+ nfactor = 1
+ pketa = -1.4647263e-15
+ ngate = 8e+20
+ k2we = 5e-5
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ ngcon = 1
+ dsub = 0.75
+ wpclm = 5.7423639e-7
+ dtox = 2.7e-10
+ ppdiblc2 = 1.3236303e-15
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ fprout = 300
+ eta0 = 0.42133333
+ etab = -0.29033333
+ xrcrg1 = 12
+ xrcrg2 = 1
+ nigbacc = 10
+ a0 = -0.63009793
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 152816.98
+ cf = 8.720500000000001e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.01190817
+ k3 = -1.8419
+ em = 1000000.0
+ ll = -1.18e-13
+ lw = 0
+ u0 = 0.012770665
+ w0 = 0
+ ua = -2.0345741e-9
+ ub = 2.0265059e-18
+ uc = 2.0750138e-11
+ ud = 0
+ wtvoff = 2.7255415e-10
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 2.33e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ pkvth0we = -1.3e-19
+ nigbinv = 10
+ capmod = 2
+ wku0we = 2e-11
+ tvoff = 0.001369836
+ vfbsdoff = 0.02
+ mobmod = 0
+ ags = -5.5534702000000005
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ cjd = 0.0012620099999999998
+ cit = 0.0010906361
+ cjs = 0.0012620099999999998
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 1.30529375e-8
+ k3b = 1.9326
+ fnoimod = 1
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ eigbinv = 1.1
+ paramchk = 1
+ ku0we = -0.0007
+ beta0 = 13
+ la0 = 4.73364e-7
+ leta0 = 0
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.020492964
+ kt1 = -0.257877
+ lk2 = -1.0161511e-8
+ kt2 = -0.061294719
+ llc = -1.18e-13
+ lln = 0.7
+ lu0 = -6.1637936e-10
+ mjd = 0.26
+ lua = -3.2409276e-17
+ mjs = 0.26
+ lub = -2.2031936e-26
+ luc = 1.3331392e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = -5.6835585e-13
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 5.4600900999999995e-9
+ pbs = 0.52
+ laigsd = 6.148791e-17
+ pk2 = 5.7885716e-16
+ pu0 = 7.5708054e-18
+ dlcig = 2.5e-9
+ prt = 0
+ pua = 1.3198419e-23
+ pub = -1.7542132e-32
+ puc = -4.6237685e-24
+ pud = 0
+ bgidl = 2320000000.0
+ ijthdfwd = 0.01
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 7.2295613e-10
+ ub1 = -3.1143135e-19
+ uc1 = 1.5561971e-10
+ tpb = 0.0014
+ wa0 = 1.5943496e-6
+ ute = -1
+ wat = -0.018189188
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -4.4652352e-10
+ keta = -0.031454297
+ cigbacc = 0.32875
+ wlc = 0
+ wln = 1
+ wu0 = -1.4484792e-10
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -8.0149958e-17
+ wub = 8.6587882e-26
+ wuc = 2.0402085e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ dmcgt = 0
+ tcjsw = 0.000357
+ lags = 2.2519967e-6
+ tnoimod = 0
+ jswd = 1.28e-13
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ jsws = 1.28e-13
+ lcit = 1.2434545e-10
+ ijthdrev = 0.01
+ kt1l = 0
+ cigbinv = 0.006
+ lpdiblc2 = -6.8002141e-9
+ bigsd = 0.00125
+ lint = 9.7879675e-9
+ lkt1 = -5.2916909e-9
+ lkt2 = -7.0897675e-9
+ lmax = 4.5075e-7
+ lmin = 2.1744e-7
+ wvoff = -5.5871857e-9
+ lpe0 = 9.2e-8
+ version = 4.5
+ lpeb = 2.5e-7
+ tempmod = 0
+ wvsat = 0.0018584193
+ wvth0 = -1.04953081e-8
+ minv = -0.3
+ lua1 = -8.8631172e-18
+ lub1 = -6.5204234e-26
+ luc1 = -1.2853813e-17
+ toxref = 3e-9
+ waigc = 3.2137522e-11
+ ndep = 1e+18
+ aigbacc = 0.02
+ lwlc = 0
+ lkvth0we = -2e-12
+ moin = 5.1
+ lketa = -1.5041313e-8
+ nigc = 3.083
+ xpart = 1
+ acnqsmod = 0
+ aigbinv = 0.0163
+ egidl = 0.29734
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ ltvoff = -1.6194017e-10
+ rbodymod = 0
+ pags = -7.8283743e-13
+ ntox = 2.029
+ pvfbsdoff = 0
+ pcit = -4.6359735e-17
+ pclm = 0.629885
+ phin = 0.15
+ lku0we = 2.5e-11
+ epsrox = 3.9
+ pkt1 = -5.4236613e-15
+ pkt2 = 1.7633117e-15
+ poxedge = 1
+ rdsmod = 0
+ igbmod = 1
+ wpdiblc2 = -4.5939646e-9
+ pvoff = 2.567445e-15
+ binunit = 2
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ rbdb = 50
+ pua1 = -2.4183981e-24
+ prwb = 0
+ prwg = 0
+ pub1 = 1.1091342e-32
+ cdscb = 0
+ cdscd = 0
+ puc1 = 5.125141e-25
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ pvsat = -2.8496404000000002e-9
+ rbsb = 50
+ pvag = 1.2
+ pbswgd = 0.95
+ pbswgs = 0.95
+ wk2we = 5e-12
+ pvth0 = 6.613032399999999e-16
+ drout = 0.56
+ rdsw = 100
+ igcmod = 1
+ paigc = 6.2688273e-19
+ voffl = 0
+ weta0 = -1.09928e-7
+ wetab = 2.7482e-8
+ wkvth0we = 2e-12
+ trnqsmod = 0
+ cgidl = 0.22
+ rshg = 15.6
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ paigsd = -5.5708045e-23
+ permod = 1
+ pbswd = 0.8
+ pbsws = 0.8
+ )

.model nch_ff_21 nmos (
+ level = 54
+ acnqsmod = 0
+ dmcgt = 0
+ version = 4.5
+ tcjsw = 0.000357
+ ptvfbsdoff = 0
+ tempmod = 0
+ rbodymod = 0
+ tpbswg = 0.0009
+ aigbacc = 0.02
+ bigsd = 0.00125
+ wvoff = 4.2089489999999885e-10
+ ptvoff = 6.7086074e-18
+ wvsat = -0.0116031636
+ waigsd = 3.0872445e-12
+ aigbinv = 0.0163
+ wvth0 = 4.2902145900000014e-9
+ wpdiblc2 = 3.4958017e-9
+ waigc = 1.7847398e-12
+ diomod = 1
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 2.6226e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.6226e-10
+ lketa = -3.6124213e-8
+ xpart = 1
+ keta = 0.068466797
+ egidl = 0.29734
+ mjswgd = 0.85
+ mjswgs = 0.85
+ wkvth0we = 2e-12
+ poxedge = 1
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ tcjswg = 0.001
+ lcit = 5.1521194000000004e-11
+ pvfbsdoff = 0
+ kt1l = 0
+ trnqsmod = 0
+ binunit = 2
+ lint = 9.7879675e-9
+ lkt1 = -3.8411747999999995e-10
+ lkt2 = 9.4878496e-10
+ lmax = 2.1744e-7
+ lmin = 9.167e-8
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ rgatemod = 0
+ minv = -0.3
+ lua1 = 1.428412e-17
+ pvoff = 1.2997136100000001e-15
+ lub1 = -6.3260104e-26
+ luc1 = -5.9196014e-18
+ tnjtsswg = 1
+ fprout = 300
+ ndep = 1e+18
+ cdscb = 0
+ cdscd = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ pvsat = -9.247134000000162e-12
+ lwlc = 0
+ wk2we = 5e-12
+ pvth0 = -2.4584174400000003e-15
+ moin = 5.1
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ drout = 0.56
+ nigc = 3.083
+ paigc = 7.0313197e-18
+ wtvoff = -2.7645419e-10
+ voffl = 0
+ noff = 2.7195
+ weta0 = -1.09928e-7
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ wetab = 2.7482e-8
+ lpclm = 5.9671804e-8
+ capmod = 2
+ wku0we = 2e-11
+ ntox = 2.029
+ cgidl = 0.22
+ pcit = -4.8161006999999996e-17
+ pclm = 0.34708024
+ mobmod = 0
+ njtsswg = 9
+ phin = 0.15
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ pkt1 = -1.1550175e-15
+ pkt2 = -1.739649e-15
+ pbswd = 0.8
+ pbsws = 0.8
+ a0 = 1.2892878
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 51380.779
+ cf = 8.720500000000001e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = -0.035282087000000004
+ k3 = -1.8419
+ em = 1000000.0
+ ckappad = 0.6
+ ckappas = 0.6
+ ll = -1.18e-13
+ lw = 0
+ u0 = 0.010899764000000001
+ w0 = 0
+ ua = -2.2703742e-9
+ ub = 2.053795462e-18
+ uc = 5.2246809e-11
+ ud = 0
+ pdiblc1 = 0
+ pdiblc2 = 0.010471563
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 2.33e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ pdiblcb = -0.3
+ rbdb = 50
+ pua1 = -9.0422848e-24
+ prwb = 0
+ pdits = 0
+ laigsd = -6.8373623e-17
+ prwg = 0
+ pub1 = 1.3277736e-32
+ puc1 = 4.9546192e-24
+ cigsd = 0.069865
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ rdsw = 100
+ ijthsfwd = 0.01
+ bigbacc = 0.002588
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ kvth0we = 0.00018
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ tnoia = 0
+ ijthsrev = 0.01
+ lintnoi = -1.5e-8
+ bigbinv = 0.004953
+ peta0 = 0
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ rshg = 15.6
+ wketa = -5.2502872e-8
+ tpbsw = 0.0019
+ cjswd = 7.625999999999999e-11
+ cjsws = 7.625999999999999e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ ppdiblc2 = -3.8331042e-16
+ toxref = 3e-9
+ tnom = 25
+ toxe = 2.3900000000000002e-9
+ toxm = 2.43e-9
+ scref = 1e-6
+ tvfbsdoff = 0.022
+ pigcd = 2.621
+ aigsd = 0.010772862
+ nfactor = 1
+ ltvoff = 9.6416574e-11
+ wags = -1.210467e-6
+ lvoff = -9.078213999999999e-10
+ pkvth0we = -1.3e-19
+ wcit = 2.1500316e-10
+ lvsat = -0.0005381747100000002
+ lvth0 = -6.296310299999999e-9
+ voff = -0.16014500000000004
+ acde = 0.4
+ delta = 0.007595625
+ laigc = -1.4310771e-11
+ vfbsdoff = 0.02
+ vsat = 114971.1026
+ wint = 0
+ vth0 = 0.39359110699999994
+ rnoia = 0
+ rnoib = 0
+ lku0we = 2.5e-11
+ wkt1 = -1.19137768e-8
+ wkt2 = 1.0152376e-8
+ nigbacc = 10
+ wmax = 8.974e-7
+ epsrox = 3.9
+ aigc = 0.011560684
+ wmin = 5.374e-7
+ wvfbsdoff = 0
+ pketa = 1.139354e-14
+ lvfbsdoff = 0
+ ngate = 8e+20
+ rdsmod = 0
+ ngcon = 1
+ paramchk = 1
+ wpclm = 8.9560432e-7
+ igbmod = 1
+ wua1 = 5.7543559e-17
+ wub1 = -8.4794537e-26
+ wuc1 = -5.6143964e-17
+ gbmin = 1e-12
+ nigbinv = 10
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ bigc = 0.001442
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ wwlc = 0
+ pbswgd = 0.95
+ pbswgs = 0.95
+ cdsc = 0
+ igcmod = 1
+ cgbo = 0
+ cgdl = 3.5522823e-12
+ cgdo = 5.2490134000000004e-11
+ xtid = 3
+ ijthdfwd = 0.01
+ xtis = 3
+ cgsl = 3.5522823e-12
+ cgso = 5.2490134000000004e-11
+ cigc = 0.000625
+ fnoimod = 1
+ eigbinv = 1.1
+ ags = 5.1194999999999995
+ ijthdrev = 0.01
+ cjd = 0.0012620099999999998
+ cit = 0.0014357747
+ cjs = 0.0012620099999999998
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 1.30529375e-8
+ paigsd = 4.6587859e-23
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ tvoff = 0.00014539643
+ lpdiblc2 = -2.045371e-10
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ permod = 1
+ la0 = 6.8373618e-8
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = 0.0009100743
+ kt1 = -0.28113564
+ lk2 = -2.0436616e-10
+ kt2 = -0.099392124
+ llc = -1.18e-13
+ lln = 0.7
+ wtvfbsdoff = 0
+ lu0 = -2.2161917e-10
+ mjd = 0.26
+ lua = 1.7344554e-17
+ mjs = 0.26
+ lub = -2.7790142600000004e-26
+ luc = -5.3126584e-18
+ lud = 0
+ k2we = 5e-5
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = -4.6587862e-14
+ nsd = 1e+20
+ dsub = 0.75
+ pbd = 0.52
+ pat = -1.8212972999999999e-9
+ pbs = 0.52
+ pk2 = -1.7344476e-15
+ cigbacc = 0.32875
+ dtox = 2.7e-10
+ ku0we = -0.0007
+ pu0 = 5.028211e-18
+ beta0 = 13
+ prt = 0
+ pua = 1.2335294e-23
+ pub = -1.88032504e-32
+ puc = -1.1996375e-24
+ pud = 0
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ leta0 = 0
+ ltvfbsdoff = 0
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 6.1325358e-10
+ ub1 = -3.2064524e-19
+ uc1 = 1.2275615e-10
+ tnoimod = 0
+ tpb = 0.0014
+ ppclm = -6.7808634e-14
+ wa0 = -8.7848444e-7
+ voffcv = -0.16942
+ wpemod = 1
+ ute = -1
+ wat = 0.016319757
+ eta0 = 0.42133333
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 1.0517006e-8
+ lkvth0we = -2e-12
+ etab = -0.29033333
+ wlc = 0
+ wln = 1
+ wu0 = -1.32797711e-10
+ xgl = -1.09e-8
+ xgw = 0
+ dlcig = 2.5e-9
+ wua = -7.6059319e-17
+ wub = 9.256491399999999e-26
+ wuc = 4.1739756e-18
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ bgidl = 2320000000.0
+ cigbinv = 0.006
+ )

.model nch_ff_22 nmos (
+ level = 54
+ phin = 0.15
+ cjswd = 7.625999999999999e-11
+ cjsws = 7.625999999999999e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ pkt1 = -2.497551e-15
+ pkt2 = 8.0276583e-16
+ ptvoff = -9.1490879e-17
+ nfactor = 1
+ paramchk = 1
+ waigsd = 3.0879615e-12
+ diomod = 1
+ rbdb = 50
+ pua1 = -1.6477593e-25
+ prwb = 0
+ prwg = 0
+ pub1 = 1.4533022e-32
+ puc1 = 1.092524e-23
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ pditsd = 0
+ pditsl = 0
+ rbsb = 50
+ pvag = 1.2
+ cjswgd = 2.6226e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.6226e-10
+ rdsw = 100
+ ijthdfwd = 0.01
+ scref = 1e-6
+ tvfbsdoff = 0.022
+ nigbacc = 10
+ pigcd = 2.621
+ aigsd = 0.010772861
+ mjswgd = 0.85
+ mjswgs = 0.85
+ lvoff = -5.168304999999995e-10
+ tcjswg = 0.001
+ lvsat = 0.0014805949840000002
+ ijthdrev = 0.01
+ lvth0 = 9.500104000000002e-10
+ nigbinv = 10
+ delta = 0.007595625
+ rshg = 15.6
+ laigc = -8.7106488e-12
+ lpdiblc2 = -4.1841324e-15
+ rnoia = 0
+ rnoib = 0
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ pketa = -2.7052976e-14
+ ngate = 8e+20
+ ngcon = 1
+ wpclm = 4.0103412e-7
+ fnoimod = 1
+ fprout = 300
+ eigbinv = 1.1
+ gbmin = 1e-12
+ tnom = 25
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ xrcrg1 = 12
+ xrcrg2 = 1
+ toxe = 2.3900000000000002e-9
+ toxm = 2.43e-9
+ lkvth0we = -2e-12
+ wtvoff = 7.682212e-10
+ ags = 5.1194999999999995
+ cjd = 0.0012620099999999998
+ cit = 0.00080536553
+ cjs = 0.0012620099999999998
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ acnqsmod = 0
+ dlc = 3.26497e-9
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ wags = -1.210467e-6
+ capmod = 2
+ wcit = 1.0996029000000003e-10
+ cigbacc = 0.32875
+ rbodymod = 0
+ wku0we = 2e-11
+ la0 = -1.9182963e-7
+ voff = -0.164304478
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.00179425008
+ acde = 0.4
+ kt1 = -0.33033037
+ lk2 = -1.3785596e-9
+ kt2 = -0.066210327
+ mobmod = 0
+ llc = 0
+ lln = 1
+ lu0 = -3.818681899999999e-11
+ tnoimod = 0
+ mjd = 0.26
+ tvoff = 0.00053139469
+ lua = 2.7860169e-17
+ mjs = 0.26
+ lub = -2.7395085e-26
+ luc = 1.41139916e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ vsat = 93494.81899999999
+ njs = 1.02
+ pa0 = 2.0809981e-13
+ wint = 0
+ vth0 = 0.316502588
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 2.0509444199999998e-9
+ pbs = 0.52
+ pk2 = 9.5324632e-16
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ wkt1 = 2.3684939e-9
+ wkt2 = -1.689459e-8
+ pu0 = -2.13571417e-17
+ wmax = 8.974e-7
+ prt = 0
+ pua = -6.3654423e-24
+ pub = 7.034010899999999e-33
+ puc = -7.127418999999999e-24
+ pud = 0
+ cigbinv = 0.006
+ aigc = 0.011501109
+ wmin = 5.374e-7
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 8.1588744e-10
+ ub1 = -6.9089562e-19
+ uc1 = 1.6549472299999998e-10
+ tpb = 0.0014
+ wa0 = -3.5879278e-6
+ ute = -1
+ wat = -0.024874303599999998
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -1.8075483e-8
+ ku0we = -0.0007
+ wlc = 0
+ wln = 1
+ wu0 = 1.4789755199999998e-10
+ xgl = -1.09e-8
+ xgw = 0
+ beta0 = 13
+ wua = 1.2288469e-16
+ wub = -1.8229956900000002e-25
+ wua1 = -3.6898024e-17
+ wuc = 6.7235478e-17
+ wud = 0
+ wub1 = -9.8148649e-26
+ wuc1 = -1.19661208e-16
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ leta0 = -1.0826782e-8
+ wpdiblc2 = -5.8202891e-10
+ letab = -2.2164189e-8
+ version = 4.5
+ bigc = 0.001442
+ laigsd = 3.8113519e-17
+ tempmod = 0
+ wwlc = 0
+ ppclm = -2.1319035e-14
+ dlcig = 2.5e-9
+ cdsc = 0
+ bgidl = 2320000000.0
+ cgbo = 0
+ cgdl = 3.5522823e-12
+ cgdo = 5.2490134000000004e-11
+ xtid = 3
+ aigbacc = 0.02
+ xtis = 3
+ cgsl = 3.5522823e-12
+ cgso = 5.2490134000000004e-11
+ cigc = 0.000625
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ dmcgt = 0
+ tcjsw = 0.000357
+ wkvth0we = 2e-12
+ aigbinv = 0.0163
+ a0 = 4.0574074
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 80150.18699999999
+ cf = 8.720500000000001e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = -0.022790667
+ k3 = -1.8419
+ em = 1000000.0
+ ll = 0
+ lw = 0
+ trnqsmod = 0
+ u0 = 0.008948356000000001
+ w0 = 0
+ ua = -2.3822425e-9
+ ub = 2.049592666e-18
+ uc = -1.5441968e-10
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 2.33e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ bigsd = 0.00125
+ wvoff = 3.044252900000001e-8
+ k2we = 5e-5
+ dsub = 0.75
+ dtox = 2.7e-10
+ wvsat = -0.015246289999999996
+ toxref = 3e-9
+ wvth0 = -3.4905183000000016e-8
+ rgatemod = 0
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ tnjtsswg = 1
+ poxedge = 1
+ waigc = 1.9067031e-10
+ eta0 = 0.53651186
+ etab = -0.054544089
+ binunit = 2
+ lketa = 6.7720908e-8
+ xpart = 1
+ ltvoff = 6.0132739e-11
+ egidl = 0.29734
+ pvfbsdoff = 0
+ lku0we = 2.5e-11
+ epsrox = 3.9
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ rdsmod = 0
+ igbmod = 1
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ pvoff = -1.5223199999999999e-15
+ pbswgd = 0.95
+ pbswgs = 0.95
+ cdscb = 0
+ cdscd = 0
+ pvsat = 3.332095999999998e-10
+ wk2we = 5e-12
+ igcmod = 1
+ pvth0 = 1.2259500000000001e-15
+ drout = 0.56
+ paigc = -1.0723924e-17
+ ijthsfwd = 0.01
+ njtsswg = 9
+ voffl = 0
+ keta = -1.0362685
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ weta0 = -2.7932191e-7
+ wetab = 6.5877739e-8
+ wtvfbsdoff = 0
+ lpclm = -1.3225653e-8
+ ckappad = 0.6
+ ckappas = 0.6
+ jswd = 1.28e-13
+ pdiblc1 = 0
+ jsws = 1.28e-13
+ pdiblc2 = 0.0082956805
+ lcit = 1.1077991e-10
+ paigsd = -2.0809977e-23
+ pdiblcb = -0.3
+ ijthsrev = 0.01
+ kt1l = 0
+ cgidl = 0.22
+ ltvfbsdoff = 0
+ permod = 1
+ lint = 0
+ lkt1 = 4.2401869e-9
+ lkt2 = -2.1703039e-9
+ lmax = 9.167e-8
+ lmin = 5.567e-8
+ pbswd = 0.8
+ pbsws = 0.8
+ bigbacc = 0.002588
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ ppdiblc2 = 5.6582339e-21
+ minv = -0.3
+ kvth0we = 0.00018
+ lua1 = -4.7634626e-18
+ lub1 = -2.8456569e-26
+ luc1 = -9.937027189999999e-18
+ voffcv = -0.16942
+ wpemod = 1
+ pdits = 0
+ ndep = 1e+18
+ lintnoi = -1.5e-8
+ cigsd = 0.069865
+ ptvfbsdoff = 0
+ lwlc = 0
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ moin = 5.1
+ vtsswgs = 4.2
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ nigc = 3.083
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ pkvth0we = -1.3e-19
+ tnoia = 0
+ tpbswg = 0.0009
+ peta0 = 1.5923028e-14
+ ntox = 2.029
+ pcit = -3.82869215e-17
+ petab = -3.6091995e-15
+ pclm = 1.1225851
+ vfbsdoff = 0.02
+ wketa = 3.5650261e-7
+ tpbsw = 0.0019
+ )

.model nch_ff_23 nmos (
+ level = 54
+ pditsl = 0
+ cjswgd = 2.6226e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.6226e-10
+ cdsc = 0
+ lketa = -2.0578185e-8
+ cgbo = 0
+ cgdl = 3.5522823e-12
+ cgdo = 5.2490134000000004e-11
+ ijthsfwd = 0.01
+ xtid = 3
+ xtis = 3
+ xpart = 1
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ cgsl = 3.5522823e-12
+ cgso = 5.2490134000000004e-11
+ cigc = 0.000625
+ mjswgd = 0.85
+ mjswgs = 0.85
+ egidl = 0.29734
+ tcjswg = 0.001
+ pvfbsdoff = 0
+ ijthsrev = 0.01
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ njtsswg = 9
+ k2we = 5e-5
+ dsub = 0.75
+ dtox = 2.7e-10
+ fprout = 300
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ xrcrg1 = 12
+ xrcrg2 = 1
+ pvoff = -3.925098540000001e-15
+ ckappad = 0.6
+ ckappas = 0.6
+ cdscb = 0
+ pdiblc1 = 0
+ pdiblc2 = 0.0082956083
+ cdscd = 0
+ pdiblcb = -0.3
+ pvsat = 3.926533010999999e-9
+ eta0 = 0.49180426
+ etab = -1.1686036
+ wk2we = 5e-12
+ pvth0 = 5.3812269e-15
+ drout = 0.56
+ wtvoff = -4.625476e-9
+ paigc = -1.7630641e-18
+ voffl = 0
+ weta0 = 1.6706711e-7
+ capmod = 2
+ bigbacc = 0.002588
+ wetab = -6.7375536e-8
+ pkvth0we = -1.3e-19
+ lpclm = -4.9784452e-8
+ wku0we = 2e-11
+ mobmod = 0
+ kvth0we = 0.00018
+ cgidl = 0.22
+ vfbsdoff = 0.02
+ lintnoi = -1.5e-8
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ pbswd = 0.8
+ pbsws = 0.8
+ paramchk = 1
+ laigsd = -3.1577826e-17
+ pdits = 0
+ cigsd = 0.069865
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ ijthdfwd = 0.01
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ keta = 0.48612964
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ nfactor = 1
+ tnoia = 0
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ ijthdrev = 0.01
+ lcit = 3.8417159999999997e-10
+ peta0 = -9.9675358e-15
+ kt1l = 0
+ petab = 4.1194905e-15
+ wketa = -1.8474011e-7
+ tpbsw = 0.0019
+ lint = 0
+ cjswd = 7.625999999999999e-11
+ cjsws = 7.625999999999999e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ lkt1 = -1.5974128000000002e-8
+ lkt2 = -1.4213753e-9
+ lmax = 5.567e-8
+ lmin = 4.667e-8
+ nigbacc = 10
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ toxref = 3e-9
+ minv = -0.3
+ lua1 = 7.7308837e-17
+ lub1 = -1.39757062e-25
+ luc1 = -7.236573999999998e-18
+ ndep = 1e+18
+ lkvth0we = -2e-12
+ nigbinv = 10
+ lwlc = 0
+ moin = 5.1
+ a0 = 11.080765
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 31524.241299999994
+ cf = 8.720500000000001e-11
+ ef = 1.0
+ k1 = 0.274
+ tvfbsdoff = 0.022
+ k2 = 0.011147898
+ k3 = -1.8419
+ em = 1000000.0
+ ll = 0
+ lw = 0
+ u0 = -0.0017551457400000001
+ scref = 1e-6
+ nigc = 3.083
+ w0 = 0
+ ua = -5.2066121e-9
+ ub = 5.20056154e-18
+ uc = 2.7090556e-10
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 2.33e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ pigcd = 2.621
+ aigsd = 0.010772862
+ ltvoff = -1.4697355e-10
+ acnqsmod = 0
+ lvoff = 1.5918058999999963e-9
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ fnoimod = 1
+ lvsat = -0.0063607503699999995
+ rbodymod = 0
+ lvth0 = -3.388415299999997e-9
+ eigbinv = 1.1
+ ntox = 2.029
+ delta = 0.007595625
+ pcit = -1.4599822999999998e-17
+ lku0we = 2.5e-11
+ pclm = 1.7529092
+ laigc = -1.8175152e-11
+ epsrox = 3.9
+ rnoia = 0
+ rnoib = 0
+ wvfbsdoff = 0
+ phin = 0.15
+ lvfbsdoff = 0
+ rdsmod = 0
+ pketa = 4.339103e-15
+ igbmod = 1
+ ngate = 8e+20
+ pkt1 = 1.1890454999999999e-14
+ pkt2 = 3.1759909e-15
+ ngcon = 1
+ wpclm = -7.2697212e-7
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ wpdiblc2 = -5.8193135e-10
+ pbswgd = 0.95
+ gbmin = 1e-12
+ pbswgs = 0.95
+ cigbacc = 0.32875
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ ags = 5.1194999999999995
+ rbdb = 50
+ pua1 = -6.2039198e-23
+ prwb = 0
+ prwg = 0
+ pub1 = 9.108448899999999e-32
+ puc1 = 1.0847755599999997e-23
+ igcmod = 1
+ wtvfbsdoff = 0
+ cjd = 0.0012620099999999998
+ cit = -0.0039082693
+ cjs = 0.0012620099999999998
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ dlc = 3.26497e-9
+ k3b = 1.9326
+ tnoimod = 0
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ rdsw = 100
+ ltvfbsdoff = 0
+ cigbinv = 0.006
+ la0 = -5.9918439e-7
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = 0.0010260548200000004
+ kt1 = 0.018192305
+ lk2 = -3.3469964e-9
+ kt2 = -0.079122889
+ llc = 0
+ lln = 1
+ lu0 = 5.8261626e-10
+ mjd = 0.26
+ lua = 1.9167361e-16
+ mjs = 0.26
+ lub = -2.101512744e-25
+ luc = -1.0554871600000002e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 1.4611928e-13
+ wkvth0we = 2e-12
+ nsd = 1e+20
+ pbd = 0.52
+ pat = -1.47353358e-9
+ pbs = 0.52
+ pk2 = 2.1253177e-15
+ paigsd = 1.0451534e-29
+ pu0 = -9.8996924e-17
+ prt = 0
+ pua = -7.1470289e-23
+ pub = 9.665873609999999e-32
+ puc = 4.556057900000002e-24
+ pud = 0
+ version = 4.5
+ rsh = 17.5
+ trnqsmod = 0
+ tcj = 0.00076
+ ua1 = -5.9915221e-10
+ ub1 = 1.22807897e-18
+ uc1 = 1.1893518999999988e-10
+ rshg = 15.6
+ tempmod = 0
+ tvoff = 0.0041021928
+ tpb = 0.0014
+ wa0 = -2.5192978e-6
+ permod = 1
+ ute = -1
+ wat = 0.035892558
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -3.8283609e-8
+ xjbvd = 1
+ xjbvs = 1
+ wlc = 0
+ wln = 1
+ lk2we = -1.5e-12
+ wu0 = 1.4865129000000002e-9
+ xgl = -1.09e-8
+ xgw = 0
+ wua = 1.2453821e-15
+ wub = -1.72755342e-24
+ wuc = -1.3420376999999993e-16
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ ptvfbsdoff = 0
+ aigbacc = 0.02
+ ku0we = -0.0007
+ beta0 = 13
+ rgatemod = 0
+ leta0 = -8.2337409e-9
+ letab = 4.245126e-8
+ voffcv = -0.16942
+ wpemod = 1
+ tnom = 25
+ tnjtsswg = 1
+ toxe = 2.3900000000000002e-9
+ toxm = 2.43e-9
+ aigbinv = 0.0163
+ ppclm = 4.4105328e-14
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ wags = -1.210467e-6
+ dmcgt = 0
+ tcjsw = 0.000357
+ wcit = -2.9844526e-10
+ tpbswg = 0.0009
+ voff = -0.20066027000000003
+ acde = 0.4
+ poxedge = 1
+ vsat = 228690.634
+ wint = 0
+ vth0 = 0.39130301399999995
+ bigsd = 0.00125
+ binunit = 2
+ wkt1 = -2.4570057999999997e-7
+ wkt2 = -5.7812263e-8
+ wmax = 8.974e-7
+ aigc = 0.01166429
+ wmin = 5.374e-7
+ ptvoff = 2.2134356e-16
+ wvoff = 7.186973409999998e-8
+ waigsd = 3.0876027e-12
+ wvsat = -0.07720017247000001
+ wua1 = 1.0299024e-15
+ wub1 = -1.41800181e-24
+ wuc1 = -1.1832528899999998e-16
+ wvth0 = -1.0654783200000001e-7
+ diomod = 1
+ bigc = 0.001442
+ waigc = 3.6172725e-11
+ wwlc = 0
+ pditsd = 0
+ )

.model nch_ff_24 nmos (
+ level = 54
+ lvsat = -0.002008701199999999
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lvth0 = 3.3387407000000002e-9
+ lcit = 4.669948800000001e-10
+ trnqsmod = 0
+ kt1l = 0
+ cigbacc = 0.32875
+ delta = 0.007595625
+ laigc = -7.4258513e-12
+ rnoia = 0
+ rnoib = 0
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ tnoimod = 0
+ lint = 0
+ lkt1 = -8.858509999999989e-11
+ lkt2 = 6.4873536e-9
+ lmax = 4.667e-8
+ pketa = 3.05233408e-14
+ ags = 5.1194999999999995
+ ngate = 8e+20
+ lmin = 3.6e-8
+ cigbinv = 0.006
+ ngcon = 1
+ lpe0 = 9.2e-8
+ cjd = 0.0012620099999999998
+ cit = -0.005598636000000001
+ fprout = 300
+ cjs = 0.0012620099999999998
+ clc = 1e-7
+ wpclm = 9.524622100000001e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ lpeb = 2.5e-7
+ dlc = 3.26497e-9
+ k3b = 1.9326
+ xrcrg1 = 12
+ xrcrg2 = 1
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ rgatemod = 0
+ gbmin = 1e-12
+ minv = -0.3
+ tnjtsswg = 1
+ lua1 = -6.7547343e-17
+ lub1 = 1.1659735399999998e-25
+ luc1 = 1.834266e-17
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ ndep = 1e+18
+ la0 = -5.581062559999999e-7
+ version = 4.5
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.00276593679
+ wtvoff = -5.6534448e-10
+ lwlc = 0
+ kt1 = -0.30600245
+ lk2 = -3.4047834e-9
+ kt2 = -0.24052552
+ llc = 0
+ moin = 5.1
+ lln = 1
+ lu0 = 8.8489725e-10
+ tempmod = 0
+ mjd = 0.26
+ lua = 1.9963428e-16
+ mjs = 0.26
+ lub = -1.86515944e-25
+ luc = -1.3855022100000003e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 1.41312605e-13
+ nigc = 3.083
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 6.996441899999999e-10
+ pbs = 0.52
+ pk2 = 1.540171e-16
+ pu0 = -4.9792621e-16
+ prt = 0
+ pua = -1.24177601e-22
+ pub = 1.2166737845000001e-31
+ puc = -3.231882900000001e-24
+ pud = 0
+ aigbacc = 0.02
+ capmod = 2
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 2.3570964e-9
+ ub1 = -4.0036457e-18
+ uc1 = -4.0308999999999995e-10
+ tpb = 0.0014
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ wku0we = 2e-11
+ wa0 = -2.4212027299999997e-6
+ ute = -1
+ wat = -0.008457981
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 1.947015e-9
+ wlc = 0
+ wln = 1
+ wu0 = 9.627935500000001e-9
+ xgl = -1.09e-8
+ mobmod = 0
+ xgw = 0
+ wua = 2.32104147e-15
+ wub = -2.2379339299999998e-24
+ wuc = 2.4733810000000014e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ ntox = 2.029
+ pcit = 9.3372643e-17
+ pclm = 0.021884800000000038
+ tvoff = 0.0045807103
+ aigbinv = 0.0163
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ phin = 0.15
+ pkt1 = -5.3485624e-15
+ pkt2 = -2.9889728e-15
+ ku0we = -0.0007
+ beta0 = 13
+ laigsd = 2.1777751e-17
+ leta0 = 6.023777099999999e-9
+ letab = 3.2196399e-8
+ ppclm = -3.8186956000000005e-14
+ rbdb = 50
+ pua1 = 5.0551945e-23
+ prwb = 0
+ prwg = 0
+ pub1 = -8.3719216e-32
+ puc1 = -1.81613879e-23
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ poxedge = 1
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ rdsw = 100
+ ijthsfwd = 0.01
+ binunit = 2
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ dmcgt = 0
+ tcjsw = 0.000357
+ ijthsrev = 0.01
+ rshg = 15.6
+ bigsd = 0.00125
+ wvoff = -2.5396920999999984e-8
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ toxref = 3e-9
+ wvsat = -0.030373111000000005
+ wvth0 = 6.1396173e-8
+ tnom = 25
+ waigc = -1.3685053e-10
+ toxe = 2.3900000000000002e-9
+ toxm = 2.43e-9
+ lketa = -4.89346675e-8
+ xpart = 1
+ ltvoff = -1.7042091e-10
+ egidl = 0.29734
+ njtsswg = 9
+ wags = -1.210467e-6
+ pkvth0we = -1.3e-19
+ pvfbsdoff = 0
+ wcit = -2.5020114e-9
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ voff = -0.003529144999999956
+ lku0we = 2.5e-11
+ acde = 0.4
+ ckappad = 0.6
+ epsrox = 3.9
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.0082956083
+ vfbsdoff = 0.02
+ pdiblcb = -0.3
+ vsat = 139873.196
+ wint = 0
+ vth0 = 0.2540148649999999
+ wkt1 = 1.0611611e-7
+ wkt2 = 6.8003321e-8
+ rdsmod = 0
+ wtvfbsdoff = 0
+ wmax = 8.974e-7
+ aigc = 0.011444916
+ wmin = 5.374e-7
+ igbmod = 1
+ a0 = 10.24243689
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 108911.802
+ cf = 8.720500000000001e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.012327223
+ k3 = -1.8419
+ em = 1000000.0
+ ll = 0
+ lw = 0
+ u0 = -0.0079241478
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ paramchk = 1
+ w0 = 0
+ ua = -5.369074800000001e-9
+ ub = 4.718207719999999e-18
+ uc = 3.3825556e-10
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 2.33e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ ltvfbsdoff = 0
+ pbswgd = 0.95
+ pbswgs = 0.95
+ wua1 = -1.2678761e-15
+ wub1 = 2.1494207099999998e-24
+ wuc1 = 4.7369808e-16
+ bigbacc = 0.002588
+ pvoff = 8.409683299999991e-16
+ bigc = 0.001442
+ igcmod = 1
+ wwlc = 0
+ cdscb = 0
+ cdscd = 0
+ kvth0we = 0.00018
+ pvsat = 1.63200933e-9
+ wk2we = 5e-12
+ pvth0 = -2.8480257000000006e-15
+ drout = 0.56
+ cdsc = 0
+ lintnoi = -1.5e-8
+ paigc = 6.7150752e-18
+ cgbo = 0
+ ijthdfwd = 0.01
+ cgdl = 3.5522823e-12
+ cgdo = 5.2490134000000004e-11
+ xtid = 3
+ xtis = 3
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ cgsl = 3.5522823e-12
+ cgso = 5.2490134000000004e-11
+ voffl = 0
+ cigc = 0.000625
+ ptvfbsdoff = 0
+ weta0 = -1.6294544599999998e-7
+ wetab = 1.0177792e-7
+ paigsd = 4.9710031e-30
+ lpclm = 3.5035747999999996e-8
+ ijthdrev = 0.01
+ cgidl = 0.22
+ permod = 1
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ pbswd = 0.8
+ pbsws = 0.8
+ k2we = 5e-5
+ dsub = 0.75
+ dtox = 2.7e-10
+ voffcv = -0.16942
+ wpemod = 1
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ nfactor = 1
+ pdits = 0
+ cigsd = 0.069865
+ eta0 = 0.20083450200000003
+ lkvth0we = -2e-12
+ etab = -0.95932067
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ acnqsmod = 0
+ nigbacc = 10
+ tpbswg = 0.0009
+ tnoia = 0
+ rbodymod = 0
+ peta0 = 6.20307972e-15
+ petab = -4.1690291e-15
+ wketa = -7.1911233e-7
+ tpbsw = 0.0019
+ nigbinv = 10
+ cjswd = 7.625999999999999e-11
+ cjsws = 7.625999999999999e-11
+ ptvoff = 2.2397114e-17
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ waigsd = 3.0876027e-12
+ diomod = 1
+ wpdiblc2 = -5.8193135e-10
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 2.6226e-10
+ pku0we = -1.5e-18
+ fnoimod = 1
+ cjswgs = 2.6226e-10
+ eigbinv = 1.1
+ tvfbsdoff = 0.022
+ scref = 1e-6
+ pigcd = 2.621
+ mjswgd = 0.85
+ aigsd = 0.010772861
+ mjswgs = 0.85
+ keta = 1.06483334
+ tcjswg = 0.001
+ lvoff = -8.067620000000001e-9
+ wkvth0we = 2e-12
+ )

.model nch_ff_25 nmos (
+ level = 54
+ fprout = 300
+ xrcrg1 = 12
+ xrcrg2 = 1
+ pvoff = 0
+ tnom = 25
+ cdscb = 0
+ cdscd = 0
+ toxe = 2.3900000000000002e-9
+ toxm = 2.43e-9
+ wtvoff = 0
+ pvsat = -1.8e-11
+ lkvth0we = -2e-12
+ wk2we = 5e-12
+ pvth0 = -2.3e-16
+ drout = 0.56
+ voffl = 0
+ capmod = 2
+ acnqsmod = 0
+ wku0we = 2e-11
+ weta0 = -1.1162667e-8
+ wags = -8.046904e-8
+ wetab = 2.2325333e-8
+ mobmod = 0
+ wcit = 3.463688e-10
+ rbodymod = 0
+ nfactor = 1
+ voff = -0.13478422
+ acde = 0.4
+ cgidl = 0.22
+ vsat = 102889.02
+ wint = 0
+ vth0 = 0.33620511999999997
+ wkt1 = -2.097059387e-9
+ wkt2 = -5.3296152e-9
+ wmax = 5.374e-7
+ aigc = 0.011779434
+ wmin = 2.674e-7
+ pbswd = 0.8
+ pbsws = 0.8
+ wua1 = -1.874362e-16
+ nigbacc = 10
+ wub1 = 1.1464267e-25
+ wuc1 = -2.7527136e-17
+ wpdiblc2 = 4.9914968e-9
+ bigc = 0.001442
+ pdits = 0
+ wwlc = 0
+ cigsd = 0.069865
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.5522823e-12
+ cgdo = 5.2490134000000004e-11
+ xtid = 3
+ nigbinv = 10
+ xtis = 3
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ cgsl = 3.5522823e-12
+ cgso = 5.2490134000000004e-11
+ cigc = 0.000625
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ wkvth0we = 2e-12
+ tnoia = 0
+ trnqsmod = 0
+ peta0 = 0
+ fnoimod = 1
+ wketa = 1.6322115e-8
+ eigbinv = 1.1
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ tpbsw = 0.0019
+ dmdg = 0
+ cjswd = 7.625999999999999e-11
+ cjsws = 7.625999999999999e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ toxref = 3e-9
+ k2we = 5e-5
+ dsub = 0.75
+ dtox = 2.7e-10
+ rgatemod = 0
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ tnjtsswg = 1
+ tvfbsdoff = 0.022
+ eta0 = 0.24044444
+ etab = -0.28088889
+ cigbacc = 0.32875
+ ltvoff = 0
+ scref = 1e-6
+ pigcd = 2.621
+ tnoimod = 0
+ aigsd = 0.010772818
+ wtvfbsdoff = 0
+ lvoff = -2e-11
+ cigbinv = 0.006
+ lvsat = -0.0003
+ lku0we = 2.5e-11
+ lvth0 = -1e-10
+ ltvfbsdoff = 0
+ epsrox = 3.9
+ delta = 0.007595625
+ ags = 0.9176066700000001
+ wvfbsdoff = 0
+ cjd = 0.0012620099999999998
+ cit = 0.000342575
+ version = 4.5
+ cjs = 0.0012620099999999998
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ lvfbsdoff = 0
+ rnoia = 0
+ rnoib = 0
+ rdsmod = 0
+ dlc = 9.8024918e-9
+ k3b = 1.9326
+ tempmod = 0
+ igbmod = 1
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ ngate = 8e+20
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ ngcon = 1
+ la0 = 0
+ wpclm = 9.3989653e-8
+ pbswgd = 0.95
+ jsd = 6.11e-7
+ pbswgs = 0.95
+ jss = 6.11e-7
+ lat = -0.0001
+ aigbacc = 0.02
+ kt1 = -0.22055704
+ kt2 = -0.0354368
+ llc = 0
+ lln = 1
+ lu0 = 6e-12
+ mjd = 0.26
+ mjs = 0.26
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ gbmin = 1e-12
+ njs = 1.02
+ pa0 = 0
+ igcmod = 1
+ nsd = 1e+20
+ pbd = 0.52
+ pat = -2.8e-11
+ jswgd = 1.28e-13
+ ptvfbsdoff = 0
+ pbs = 0.52
+ jswgs = 1.28e-13
+ pu0 = 2e-18
+ prt = 0
+ pud = 0
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 1.6212811e-9
+ ub1 = -8.7849211e-19
+ uc1 = 6.9356e-11
+ tpb = 0.0014
+ aigbinv = 0.0163
+ wa0 = -1.17208e-8
+ ijthsfwd = 0.01
+ ute = -1
+ wat = 0.071441067
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 1.8596306e-9
+ wlc = 0
+ wln = 1
+ wu0 = -1.3197067000000002e-9
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -1.3097991e-16
+ wub = 9.54408e-26
+ wuc = -2.4557867e-18
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ keta = -0.084351302
+ a0 = 3.5424667
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = -58844.444
+ cf = 8.720500000000001e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.018167646000000003
+ k3 = -1.8419
+ em = 1000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.017271111
+ jswd = 1.28e-13
+ w0 = 0
+ jsws = 1.28e-13
+ ijthsrev = 0.01
+ ua = -1.6762565e-9
+ ub = 2.0222e-18
+ uc = 6.1497778e-11
+ ud = 0
+ lcit = -1e-11
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 2.33e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ permod = 1
+ kt1l = 0
+ tvoff = 0.0017628809
+ xjbvd = 1
+ xjbvs = 1
+ poxedge = 1
+ lk2we = -1.5e-12
+ lint = 6.5375218e-9
+ lkt1 = -1.1e-9
+ lmax = 2.001e-5
+ binunit = 2
+ lmin = 9.00077e-6
+ lpe0 = 9.2e-8
+ voffcv = -0.16942
+ wpemod = 1
+ lpeb = 2.5e-7
+ ku0we = -0.0007
+ beta0 = 13
+ leta0 = 0
+ minv = -0.3
+ lub1 = 0
+ ndep = 1e+18
+ lwlc = 0
+ dlcig = 2.5e-9
+ moin = 5.1
+ bgidl = 2320000000.0
+ nigc = 3.083
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ noff = 2.7195
+ dmcgt = 0
+ noia = 3.11e+42
+ noib = 1.22e+22
+ pkvth0we = -1.3e-19
+ noic = 45200000.0
+ tpbswg = 0.0009
+ tcjsw = 0.000357
+ ntox = 2.029
+ pcit = -1.5e-17
+ pclm = 1.5094578
+ vfbsdoff = 0.02
+ bigsd = 0.00125
+ ptvoff = 0
+ phin = 0.15
+ waigsd = 3.1112026e-12
+ wvoff = 1.3685577e-8
+ pkt1 = -5e-17
+ paramchk = 1
+ diomod = 1
+ wvsat = -0.0028059037
+ wvth0 = -2.1768414e-8
+ njtsswg = 9
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 2.6226e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.6226e-10
+ waigc = 2.8724444e-11
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ rbdb = 50
+ prwb = 0
+ prwg = 0
+ pub1 = 0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.0047029422
+ rdsw = 100
+ pdiblcb = -0.3
+ ijthdfwd = 0.01
+ mjswgd = 0.85
+ xpart = 1
+ mjswgs = 0.85
+ tcjswg = 0.001
+ egidl = 0.29734
+ pvfbsdoff = 0
+ bigbacc = 0.002588
+ ijthdrev = 0.01
+ rshg = 15.6
+ kvth0we = 0.00018
+ lintnoi = -1.5e-8
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ )

.model nch_ff_26 nmos (
+ level = 54
+ poxedge = 1
+ capmod = 2
+ wku0we = 2e-11
+ binunit = 2
+ mobmod = 0
+ pkvth0we = -1.3e-19
+ tvoff = 0.0019388906
+ vfbsdoff = 0.02
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ laigsd = -2.019482e-16
+ paramchk = 1
+ ku0we = -0.0007
+ beta0 = 13
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ leta0 = 0
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ ijthdfwd = 0.01
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ keta = -0.091670067
+ dmcgt = 0
+ tcjsw = 0.000357
+ lags = -1.7808411e-7
+ njtsswg = 9
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ ijthdrev = 0.01
+ lcit = 6.5778289e-10
+ kt1l = 0
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ lpdiblc2 = 2.6261368e-8
+ bigsd = 0.00125
+ ckappad = 0.6
+ ckappas = 0.6
+ lint = 6.5375218e-9
+ pdiblc1 = 0
+ pdiblc2 = 0.0017817666
+ toxref = 3e-9
+ pdiblcb = -0.3
+ lkt1 = 7.9572759e-9
+ lkt2 = -2.1662043e-8
+ lmax = 9.00077e-6
+ wvoff = 1.395365e-8
+ lmin = 9.0075e-7
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ wvsat = -0.0028059037
+ wvth0 = -2.2116317e-8
+ minv = -0.3
+ wtvfbsdoff = 0
+ lua1 = -8.9279603e-16
+ lub1 = 6.8544226e-25
+ luc1 = -5.9256432e-18
+ waigc = 2.989874e-11
+ bigbacc = 0.002588
+ ndep = 1e+18
+ lkvth0we = -2e-12
+ lwlc = 0
+ moin = 5.1
+ ltvoff = -1.582327e-9
+ ltvfbsdoff = 0
+ lketa = 6.5795695e-8
+ kvth0we = 0.00018
+ nigc = 3.083
+ xpart = 1
+ lintnoi = -1.5e-8
+ acnqsmod = 0
+ pvfbsdoff = 0
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ egidl = 0.29734
+ vtsswgs = 4.2
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ lku0we = 2.5e-11
+ rbodymod = 0
+ epsrox = 3.9
+ pags = 1.7531187e-13
+ ntox = 2.029
+ pcit = -1.2198337e-16
+ pclm = 1.5094578
+ rdsmod = 0
+ ptvfbsdoff = 0
+ igbmod = 1
+ phin = 0.15
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ pbswgd = 0.95
+ pkt1 = -2.7427875e-14
+ pkt2 = -4.4253241e-16
+ pbswgs = 0.95
+ igcmod = 1
+ wpdiblc2 = 5.7318301e-9
+ pvoff = -2.4099793e-15
+ cdscb = 0
+ cdscd = 0
+ rbdb = 50
+ pua1 = 1.9942546e-22
+ prwb = 0
+ prwg = 0
+ pub1 = -1.9939615e-31
+ puc1 = 1.7835157e-23
+ nfactor = 1
+ pvsat = -1.8e-11
+ rbpb = 50
+ rbpd = 50
+ wk2we = 5e-12
+ rbps = 50
+ pvth0 = 2.8976502e-15
+ rbsb = 50
+ pvag = 1.2
+ drout = 0.56
+ rdsw = 100
+ paigc = -1.0556924e-17
+ voffl = 0
+ paigsd = 1.1026372e-22
+ weta0 = -1.1162667e-8
+ wetab = 2.2325333e-8
+ wkvth0we = 2e-12
+ nigbacc = 10
+ permod = 1
+ trnqsmod = 0
+ cgidl = 0.22
+ rshg = 15.6
+ nigbinv = 10
+ pbswd = 0.8
+ pbsws = 0.8
+ voffcv = -0.16942
+ wpemod = 1
+ rgatemod = 0
+ tnjtsswg = 1
+ tnom = 25
+ pdits = 0
+ toxe = 2.3900000000000002e-9
+ toxm = 2.43e-9
+ a0 = 3.8452644
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ cigsd = 0.069865
+ b1 = 0
+ at = -81312.781
+ cf = 8.720500000000001e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.019723392
+ k3 = -1.8419
+ em = 1000000.0
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ ll = 0
+ lw = 0
+ u0 = 0.017524559999999998
+ w0 = 0
+ fnoimod = 1
+ ua = -1.6436128e-9
+ ub = 2.0158412e-18
+ uc = 5.8736458e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 2.33e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ eigbinv = 1.1
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ tpbswg = 0.0009
+ wags = -9.9969804e-8
+ wcit = 3.5826906e-10
+ tnoia = 0
+ voff = -0.13348839
+ peta0 = 0
+ acde = 0.4
+ wketa = 1.8850903e-8
+ vsat = 102889.02
+ ptvoff = 2.7553621e-16
+ wint = 0
+ tpbsw = 0.0019
+ vth0 = 0.33049777999999996
+ cigbacc = 0.32875
+ waigsd = 3.1111904e-12
+ wkt1 = 9.483104999999998e-10
+ wkt2 = -5.2803902e-9
+ cjswd = 7.625999999999999e-11
+ cjsws = 7.625999999999999e-11
+ wmax = 5.374e-7
+ mjswd = 0.11
+ aigc = 0.011795195
+ mjsws = 0.11
+ wmin = 2.674e-7
+ agidl = 9.41e-8
+ diomod = 1
+ tnoimod = 0
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 2.6226e-10
+ pku0we = -1.5e-18
+ wua1 = -2.0961923e-16
+ wub1 = 1.3682244e-25
+ cjswgs = 2.6226e-10
+ wuc1 = -2.9511024e-17
+ cigbinv = 0.006
+ bigc = 0.001442
+ wwlc = 0
+ tvfbsdoff = 0.022
+ cdsc = 0
+ mjswgd = 0.85
+ mjswgs = 0.85
+ scref = 1e-6
+ version = 4.5
+ ijthsfwd = 0.01
+ cgbo = 0
+ cgdl = 3.5522823e-12
+ cgdo = 5.2490134000000004e-11
+ xtid = 3
+ xtis = 3
+ pigcd = 2.621
+ cgsl = 3.5522823e-12
+ tcjswg = 0.001
+ cgso = 5.2490134000000004e-11
+ tempmod = 0
+ aigsd = 0.010772818
+ cigc = 0.000625
+ ags = 0.9374157999999999
+ lvoff = -1.1669524999999999e-8
+ cjd = 0.0012620099999999998
+ cit = 0.00026829437
+ cjs = 0.0012620099999999998
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ aigbacc = 0.02
+ dlc = 9.8024918e-9
+ lvsat = -0.0003
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ lvth0 = 5.1208999e-8
+ ijthsrev = 0.01
+ delta = 0.007595625
+ laigc = -1.416882e-10
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ la0 = -2.722152e-6
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ rnoia = 0
+ rnoib = 0
+ dmdg = 0
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = 0.20189035000000002
+ kt1 = -0.22156452
+ lk2 = -1.3986155e-8
+ kt2 = -0.033027229
+ llc = 0
+ lln = 1
+ lu0 = -2.2725025999999998e-9
+ mjd = 0.26
+ aigbinv = 0.0163
+ lua = -2.9346741e-16
+ mjs = 0.26
+ lub = 5.7165214e-26
+ luc = 2.4824263e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 3.4236885e-13
+ fprout = 300
+ nsd = 1e+20
+ pbd = 0.52
+ pat = -6.371632400000001e-8
+ pbs = 0.52
+ pketa = -2.2733801e-14
+ pk2 = -1.3939214e-15
+ ngate = 8e+20
+ pu0 = 1.6739558e-16
+ xrcrg1 = 12
+ xrcrg2 = 1
+ k2we = 5e-5
+ prt = 0
+ pua = 4.226297e-23
+ pub = -4.4156209e-32
+ puc = -1.0695581e-23
+ pud = 0
+ ngcon = 1
+ wpclm = 9.3989653e-8
+ dsub = 0.75
+ rsh = 17.5
+ tcj = 0.00076
+ dtox = 2.7e-10
+ ua1 = 1.720591e-9
+ ub1 = -9.5473708e-19
+ uc1 = 7.0015137e-11
+ ppdiblc2 = -6.6555967e-15
+ tpb = 0.0014
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ wa0 = -4.9804098e-8
+ gbmin = 1e-12
+ ute = -1
+ wat = 0.078525419
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 2.0146831e-9
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ wtvoff = -3.0649189e-11
+ wlc = 0
+ wln = 1
+ wu0 = -1.3381044000000001e-9
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -1.3568102e-16
+ wub = 1.003525e-25
+ wuc = -1.2660669e-18
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ eta0 = 0.24044444
+ etab = -0.28088889
+ )

.model nch_ff_27 nmos (
+ level = 54
+ ntox = 2.029
+ pcit = -1.3105802e-16
+ pclm = 1.5094578
+ fnoimod = 1
+ phin = 0.15
+ eigbinv = 1.1
+ pbswd = 0.8
+ pbsws = 0.8
+ pkt1 = 4.762844300000001e-15
+ pkt2 = 2.2738921e-15
+ pdits = 0
+ rbdb = 50
+ pua1 = -2.6369043e-23
+ prwb = 0
+ prwg = 0
+ pub1 = 4.8759292e-32
+ cigsd = 0.069865
+ puc1 = 6.8677984e-24
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ dvt0w = 0
+ pvag = 1.2
+ dvt1w = 0
+ dvt2w = 0
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ rdsw = 100
+ ijthsfwd = 0.01
+ cigbacc = 0.32875
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ tnoimod = 0
+ tnoia = 0
+ ijthsrev = 0.01
+ cigbinv = 0.006
+ peta0 = 0
+ rshg = 15.6
+ wketa = -2.2122195e-8
+ wtvfbsdoff = 0
+ tpbsw = 0.0019
+ toxref = 3e-9
+ cjswd = 7.625999999999999e-11
+ cjsws = 7.625999999999999e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ version = 4.5
+ ltvfbsdoff = 0
+ tempmod = 0
+ ppdiblc2 = 1.7501102e-15
+ tnom = 25
+ aigbacc = 0.02
+ tvfbsdoff = 0.022
+ toxe = 2.3900000000000002e-9
+ toxm = 2.43e-9
+ ltvoff = 1.3913801e-9
+ ags = 0.26766657
+ scref = 1e-6
+ cjd = 0.0012620099999999998
+ cit = 0.00059502911
+ cjs = 0.0012620099999999998
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 9.8024918e-9
+ pigcd = 2.621
+ k3b = 1.9326
+ aigsd = 0.010772818
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ ptvfbsdoff = 0
+ aigbinv = 0.0163
+ lvoff = -5.213220300000001e-10
+ wags = 3.6984035999999996e-7
+ lku0we = 2.5e-11
+ pkvth0we = -1.3e-19
+ la0 = 3.6355951e-7
+ epsrox = 3.9
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.052838453
+ kt1 = -0.19312528
+ lk2 = -1.4722356e-8
+ kt2 = -0.039065148
+ wcit = 3.6846529999999997e-10
+ lvsat = -0.0003
+ llc = 0
+ lln = 1
+ lu0 = -1.7456993e-9
+ mjd = 0.26
+ lvth0 = -8.315815599999999e-9
+ lua = -1.1159069e-16
+ mjs = 0.26
+ lub = -2.3732546e-26
+ luc = -2.9405776e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ voff = -0.14601446
+ njs = 1.02
+ pa0 = -3.8856002e-13
+ nsd = 1e+20
+ delta = 0.007595625
+ acde = 0.4
+ pbd = 0.52
+ wvfbsdoff = 0
+ pat = -8.8162363e-10
+ pbs = 0.52
+ rdsmod = 0
+ pk2 = 1.1847359e-15
+ lvfbsdoff = 0
+ laigc = -3.3762752e-11
+ pu0 = 1.3168191e-16
+ vfbsdoff = 0.02
+ igbmod = 1
+ prt = 0
+ pua = 2.9945529e-23
+ pub = -3.9782718e-32
+ puc = 6.3626704e-24
+ pud = 0
+ vsat = 102889.02
+ wint = 0
+ rnoia = 0
+ rnoib = 0
+ vth0 = 0.39737958999999995
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 6.6639379e-10
+ ub1 = 1.1665789e-19
+ uc1 = 5.9635906e-11
+ wkt1 = -3.5221037e-8
+ wkt2 = -8.3325526e-9
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ tpb = 0.0014
+ wmax = 5.374e-7
+ wa0 = 7.714643e-7
+ aigc = 0.01167393
+ wmin = 2.674e-7
+ ute = -1
+ wat = 0.0079246317
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -8.8268726e-10
+ pbswgd = 0.95
+ pketa = 1.3732256e-14
+ poxedge = 1
+ pbswgs = 0.95
+ ngate = 8e+20
+ wlc = 0
+ wln = 1
+ wu0 = -1.2979767e-9
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -1.218412e-16
+ wub = 9.5438468e-26
+ wuc = -2.0432641e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ ngcon = 1
+ paramchk = 1
+ wpclm = 9.3989653e-8
+ igcmod = 1
+ binunit = 2
+ wua1 = 4.4082452e-17
+ wub1 = -1.420039e-25
+ wuc1 = -1.718815e-17
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ bigc = 0.001442
+ wwlc = 0
+ cdsc = 0
+ ijthdfwd = 0.01
+ cgbo = 0
+ cgdl = 3.5522823e-12
+ cgdo = 5.2490134000000004e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.5522823e-12
+ cgso = 5.2490134000000004e-11
+ cigc = 0.000625
+ permod = 1
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ ijthdrev = 0.01
+ tvoff = -0.0014023534
+ lpdiblc2 = -7.3119259e-9
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ voffcv = -0.16942
+ wpemod = 1
+ k2we = 5e-5
+ ku0we = -0.0007
+ dsub = 0.75
+ dtox = 2.7e-10
+ beta0 = 13
+ leta0 = 0
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ njtsswg = 9
+ lkvth0we = -2e-12
+ eta0 = 0.24044444
+ etab = -0.28088889
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.039504569
+ pdiblcb = -0.3
+ tpbswg = 0.0009
+ acnqsmod = 0
+ dmcgt = 0
+ tcjsw = 0.000357
+ rbodymod = 0
+ ptvoff = -5.8159511e-16
+ bigbacc = 0.002588
+ waigsd = 3.1113143e-12
+ bigsd = 0.00125
+ a0 = 0.37817284
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 204899.36
+ cf = 8.720500000000001e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.02055059
+ k3 = -1.8419
+ em = 1000000.0
+ kvth0we = 0.00018
+ diomod = 1
+ ll = 0
+ lw = 0
+ u0 = 0.016932646
+ w0 = 0
+ wvoff = 1.6411259e-8
+ ua = -1.8479686e-9
+ ub = 2.1067376e-18
+ uc = 1.1966909e-10
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 2.33e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ lintnoi = -1.5e-8
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 2.6226e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.6226e-10
+ bigbinv = 0.004953
+ wvsat = -0.0028059037
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ wvth0 = -2.5299760999999998e-8
+ wpdiblc2 = -3.7127843e-9
+ waigc = 2.313153e-11
+ mjswgd = 0.85
+ mjswgs = 0.85
+ lketa = -4.8021757e-8
+ tcjswg = 0.001
+ xpart = 1
+ pvfbsdoff = 0
+ keta = 0.03621471
+ egidl = 0.29734
+ wkvth0we = 2e-12
+ lags = 4.1799271e-7
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 3.6698897e-10
+ trnqsmod = 0
+ kt1l = 0
+ nfactor = 1
+ lint = 6.5375218e-9
+ fprout = 300
+ lkt1 = -1.7353643e-8
+ lkt2 = -1.6288295e-8
+ xrcrg1 = 12
+ xrcrg2 = 1
+ lmax = 9.0075e-7
+ lmin = 4.5075e-7
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ rgatemod = 0
+ wtvoff = 9.3241971e-10
+ pvoff = -4.5972513e-15
+ minv = -0.3
+ tnjtsswg = 1
+ lua1 = 4.5439491e-17
+ lub1 = -2.6809927e-25
+ luc1 = 3.3118724e-18
+ cdscb = 0
+ cdscd = 0
+ nigbacc = 10
+ ndep = 1e+18
+ pvsat = -1.8e-11
+ wk2we = 5e-12
+ pvth0 = 5.7309158e-15
+ lwlc = 0
+ drout = 0.56
+ moin = 5.1
+ capmod = 2
+ paigc = -4.5341069e-18
+ nigc = 3.083
+ voffl = 0
+ wku0we = 2e-11
+ nigbinv = 10
+ mobmod = 0
+ weta0 = -1.1162667e-8
+ wetab = 2.2325333e-8
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ pags = -2.4281917e-13
+ cgidl = 0.22
+ )

.model nch_ff_28 nmos (
+ level = 54
+ wuc1 = -1.3268706e-17
+ bigc = 0.001442
+ ppclm = -7.9196439e-14
+ wwlc = 0
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ cdsc = 0
+ bigbacc = 0.002588
+ cgbo = 0
+ cgdl = 3.5522823e-12
+ cgdo = 5.2490134000000004e-11
+ xtid = 3
+ xtis = 3
+ wtvfbsdoff = 0
+ cgsl = 3.5522823e-12
+ cgso = 5.2490134000000004e-11
+ cigc = 0.000625
+ kvth0we = 0.00018
+ dmcgt = 0
+ tcjsw = 0.000357
+ wkvth0we = 2e-12
+ lintnoi = -1.5e-8
+ ltvfbsdoff = 0
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ trnqsmod = 0
+ toxref = 3e-9
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ bigsd = 0.00125
+ wvoff = 5.1767953e-9
+ k2we = 5e-5
+ dsub = 0.75
+ wvsat = -0.0054199005
+ dtox = 2.7e-10
+ ptvfbsdoff = 0
+ wvth0 = -7.6869543e-9
+ rgatemod = 0
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ tnjtsswg = 1
+ waigc = -1.6608588e-12
+ ltvoff = -7.6859018e-11
+ eta0 = 0.24044444
+ etab = -0.28088889
+ lketa = -5.7215427e-9
+ nfactor = 1
+ xpart = 1
+ pvfbsdoff = 0
+ lku0we = 2.5e-11
+ egidl = 0.29734
+ epsrox = 3.9
+ rdsmod = 0
+ igbmod = 1
+ nigbacc = 10
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ pbswgd = 0.95
+ pbswgs = 0.95
+ igcmod = 1
+ nigbinv = 10
+ pvoff = 3.4591262e-16
+ cdscb = 0
+ cdscd = 0
+ pvsat = 1.1321586000000001e-9
+ wk2we = 5e-12
+ pvth0 = -2.0187192e-15
+ drout = 0.56
+ paigc = 6.374544e-18
+ ijthsfwd = 0.01
+ paigsd = 2.2627557e-23
+ voffl = 0
+ fnoimod = 1
+ eigbinv = 1.1
+ keta = -0.05992214
+ weta0 = -1.1162667e-8
+ wetab = 2.2325333e-8
+ permod = 1
+ lpclm = 1.4504842e-7
+ lags = 5.906061e-7
+ jswd = 1.28e-13
+ ijthsrev = 0.01
+ jsws = 1.28e-13
+ lcit = 8.3365571e-11
+ cgidl = 0.22
+ kt1l = 0
+ lint = 9.7879675e-9
+ voffcv = -0.16942
+ wpemod = 1
+ lkt1 = 7.7603069e-9
+ lkt2 = -2.5638367e-9
+ lmax = 4.5075e-7
+ cigbacc = 0.32875
+ pbswd = 0.8
+ pbsws = 0.8
+ lmin = 2.1744e-7
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ ppdiblc2 = -5.242001e-17
+ tnoimod = 0
+ minv = -0.3
+ lua1 = -4.6794128e-17
+ lub1 = -3.2889654e-26
+ luc1 = -2.1335001e-17
+ pdits = 0
+ ndep = 1e+18
+ cigsd = 0.069865
+ cigbinv = 0.006
+ dvt0w = 0
+ lwlc = 0
+ dvt1w = 0
+ dvt2w = 0
+ moin = 5.1
+ nigc = 3.083
+ tpbswg = 0.0009
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ version = 4.5
+ tempmod = 0
+ pkvth0we = -1.3e-19
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ tnoia = 0
+ pags = 1.2428184e-13
+ peta0 = 0
+ ptvoff = -1.5558646e-16
+ aigbacc = 0.02
+ ntox = 2.029
+ pcit = -2.39847229e-17
+ pclm = 1.1798023
+ waigsd = 3.1112628e-12
+ wketa = 2.3981389e-8
+ vfbsdoff = 0.02
+ tpbsw = 0.0019
+ cjswd = 7.625999999999999e-11
+ cjsws = 7.625999999999999e-11
+ diomod = 1
+ mjswd = 0.11
+ phin = 0.15
+ mjsws = 0.11
+ agidl = 9.41e-8
+ pditsd = 0
+ pditsl = 0
+ aigbinv = 0.0163
+ pkt1 = -1.2550052000000001e-14
+ pkt2 = -7.0784646e-16
+ cjswgd = 2.6226e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.6226e-10
+ paramchk = 1
+ ags = -0.12463658400000001
+ cjd = 0.0012620099999999998
+ tvfbsdoff = 0.022
+ cit = 0.0012396277
+ cjs = 0.0012620099999999998
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 1.30529375e-8
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ rbdb = 50
+ pua1 = 1.8291934e-23
+ prwb = 0
+ prwg = 0
+ pub1 = -6.5524188e-33
+ puc1 = 5.143243e-24
+ mjswgd = 0.85
+ mjswgs = 0.85
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ tcjswg = 0.001
+ rdsw = 100
+ scref = 1e-6
+ ijthdfwd = 0.01
+ la0 = -6.0902319e-7
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.015136937999999999
+ kt1 = -0.25020244
+ lk2 = -1.0681005e-8
+ kt2 = -0.070257098
+ pigcd = 2.621
+ llc = -1.18e-13
+ lln = 0.7
+ aigsd = 0.010772818
+ lu0 = -6.9983626e-10
+ mjd = 0.26
+ lua = -1.8564943e-17
+ mjs = 0.26
+ lub = -5.2748233e-26
+ luc = -4.2757753e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 2.2627554e-14
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 2.5357001000000003e-9
+ poxedge = 1
+ pbs = 0.52
+ pk2 = 8.6250113e-16
+ lvoff = -7.167449400000001e-9
+ a0 = 2.5885881
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ pu0 = 5.3138272000000005e-17
+ at = 119214.09
+ cf = 8.720500000000001e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.011365692
+ k3 = -1.8419
+ em = 1000000.0
+ prt = 0
+ pua = 5.6394132e-24
+ pub = -7.710339e-34
+ puc = -1.5613012e-24
+ pud = 0
+ ll = -1.18e-13
+ lw = 0
+ u0 = 0.014555684000000001
+ w0 = 0
+ ua = -2.0593908e-9
+ ub = 2.1726824e-18
+ uc = 6.2555449e-11
+ ud = 0
+ wl = 0
+ rsh = 17.5
+ wr = 1
+ xj = 8.6e-8
+ xl = 2.33e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ tcj = 0.00076
+ ua1 = 8.7601565e-10
+ lvsat = -0.0044672412
+ ub1 = -4.1790941e-19
+ uc1 = 1.1565153e-10
+ binunit = 2
+ lvth0 = 1.374398e-9
+ ijthdrev = 0.01
+ tpb = 0.0014
+ wvfbsdoff = 0
+ wa0 = -1.6305293e-7
+ lvfbsdoff = 0
+ ute = -1
+ wat = 0.00015798693
+ delta = 0.007595625
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -1.5033038e-10
+ laigc = -3.7429738e-11
+ wlc = 0
+ wln = 1
+ rshg = 15.6
+ wu0 = -1.1194684000000002e-9
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -6.6600022e-17
+ wub = 6.7755498e-27
+ wuc = -2.4236148e-18
+ wud = 0
+ lpdiblc2 = -4.2799755e-9
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ rnoia = 0
+ rnoib = 0
+ fprout = 300
+ xrcrg1 = 12
+ xrcrg2 = 1
+ pketa = -6.5533207e-15
+ ngate = 8e+20
+ ngcon = 1
+ wpclm = 2.7398156e-7
+ wtvoff = -3.5781771e-11
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ tnom = 25
+ jswgs = 1.28e-13
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ toxe = 2.3900000000000002e-9
+ toxm = 2.43e-9
+ lkvth0we = -2e-12
+ capmod = 2
+ wku0we = 2e-11
+ mobmod = 0
+ acnqsmod = 0
+ wags = -4.6448013000000004e-7
+ wcit = 1.25116891e-10
+ rbodymod = 0
+ voff = -0.13090963
+ acde = 0.4
+ tvoff = 0.0019345538
+ njtsswg = 9
+ vsat = 112360.02
+ wint = 0
+ xjbvd = 1
+ xjbvs = 1
+ vth0 = 0.37535638
+ lk2we = -1.5e-12
+ wkt1 = 4.1264547999999994e-9
+ wkt2 = -1.5558741e-9
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ wmax = 5.374e-7
+ laigsd = -8.1983894e-17
+ aigc = 0.011682264
+ wmin = 2.674e-7
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.032613772
+ pdiblcb = -0.3
+ ku0we = -0.0007
+ beta0 = 13
+ leta0 = 0
+ wua1 = -5.7419768e-17
+ wpdiblc2 = 3.8387521e-10
+ wub1 = -1.6295463e-26
+ )

.model nch_ff_29 nmos (
+ level = 54
+ keta = 0.0092481698
+ aigbinv = 0.0163
+ tnoia = 0
+ ijthdrev = 0.01
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = -2.3537106e-11
+ peta0 = 0
+ ptvfbsdoff = 0
+ kt1l = 0
+ wketa = -2.0169501e-8
+ toxref = 3e-9
+ lpdiblc2 = -9.0824285e-10
+ tpbsw = 0.0019
+ ags = 2.6744444
+ cjswd = 7.625999999999999e-11
+ cjsws = 7.625999999999999e-11
+ lint = 9.7879675e-9
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ cjd = 0.0012620099999999998
+ cit = 0.0017462755
+ cjs = 0.0012620099999999998
+ clc = 1e-7
+ cle = 0.6
+ lkt1 = -3.6262126e-9
+ bvd = 8.7
+ lkt2 = -3.9513595e-9
+ bvs = 8.7
+ lmax = 2.1744e-7
+ dlc = 1.30529375e-8
+ lmin = 9.167e-8
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ poxedge = 1
+ tvfbsdoff = 0.022
+ la0 = -2.075695e-7
+ minv = -0.3
+ jsd = 6.11e-7
+ ltvoff = 5.8839234e-11
+ jss = 6.11e-7
+ lat = -0.0016937311
+ lua1 = -5.8912951e-18
+ lub1 = -2.9377439e-26
+ luc1 = 1.0640856e-17
+ kt1 = -0.1962379
+ lk2 = -3.2022951e-9
+ kt2 = -0.063681161
+ llc = -1.18e-13
+ binunit = 2
+ lln = 0.7
+ lu0 = -2.4951767000000005e-10
+ mjd = 0.26
+ lua = 5.2959027e-17
+ mjs = 0.26
+ lub = -7.97606935e-26
+ luc = -8.8267893e-18
+ lud = 0
+ lwc = 0
+ ndep = 1e+18
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ lkvth0we = -2e-12
+ njs = 1.02
+ pa0 = 1.0407708e-13
+ nsd = 1e+20
+ lwlc = 0
+ pbd = 0.52
+ pat = -3.9961951e-10
+ pbs = 0.52
+ pk2 = -9.7578421e-17
+ moin = 5.1
+ pu0 = 2.0260797000000002e-17
+ prt = 0
+ pua = -7.1102082e-24
+ pub = 9.57267e-33
+ puc = 7.19078e-25
+ pud = 0
+ scref = 1e-6
+ nigc = 3.083
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 6.8216336e-10
+ pigcd = 2.621
+ ub1 = -4.3455498e-19
+ uc1 = -3.5892821e-11
+ aigsd = 0.010772818
+ tpb = 0.0014
+ lku0we = 2.5e-11
+ wa0 = -5.4906963e-7
+ acnqsmod = 0
+ ute = -1
+ wat = 0.014069454
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 4.3998097e-9
+ epsrox = 3.9
+ lvoff = 2.3123665299999996e-9
+ wlc = 0
+ wln = 1
+ wu0 = -9.6365099e-10
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -6.1752756e-18
+ wub = -4.2246744000000004e-26
+ wuc = -1.3231099e-17
+ wud = 0
+ wwc = 0
+ noff = 2.7195
+ wwl = 0
+ wwn = 1
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ lvsat = -0.0007573482699999999
+ rbodymod = 0
+ rdsmod = 0
+ wvfbsdoff = 0
+ lvth0 = -1.2294990599999999e-8
+ lvfbsdoff = 0
+ igbmod = 1
+ delta = 0.007595625
+ laigc = 2.6175146e-12
+ ntox = 2.029
+ pcit = -7.1791752e-18
+ jtsswgd = 2.3e-7
+ pclm = 2.3689724
+ jtsswgs = 2.3e-7
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ rnoia = 0
+ rnoib = 0
+ pbswgd = 0.95
+ pbswgs = 0.95
+ phin = 0.15
+ pketa = 2.762517e-15
+ ngate = 8e+20
+ igcmod = 1
+ ngcon = 1
+ pkt1 = 6.151664499999999e-16
+ pkt2 = 9.3582987e-16
+ wpclm = -2.0834879e-7
+ wpdiblc2 = 1.3111248e-10
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ rbdb = 50
+ pua1 = 1.9734917e-24
+ prwb = 0
+ prwg = 0
+ pub1 = -5.2222001e-33
+ puc1 = -4.0873907e-24
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ njtsswg = 9
+ paigsd = -9.4615512e-24
+ rdsw = 100
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ permod = 1
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.016633997
+ pdiblcb = -0.3
+ wkvth0we = 2e-12
+ trnqsmod = 0
+ tvoff = 0.0012914341
+ rshg = 15.6
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ voffcv = -0.16942
+ wpemod = 1
+ bigbacc = 0.002588
+ ku0we = -0.0007
+ kvth0we = 0.00018
+ beta0 = 13
+ leta0 = 0
+ rgatemod = 0
+ lintnoi = -1.5e-8
+ tnjtsswg = 1
+ tnom = 25
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ ppclm = 2.2575265e-14
+ vtsswgs = 4.2
+ toxe = 2.3900000000000002e-9
+ toxm = 2.43e-9
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ tpbswg = 0.0009
+ dmcgt = 0
+ wags = 1.2453333e-7
+ tcjsw = 0.000357
+ wcit = 4.54697462e-11
+ ptvoff = 2.7225835e-17
+ voff = -0.175837897
+ waigsd = 3.1114149e-12
+ acde = 0.4
+ vsat = 94777.65030000001
+ wint = 0
+ bigsd = 0.00125
+ vth0 = 0.44014045399999996
+ diomod = 1
+ wkt1 = -5.8267946e-8
+ wkt2 = -9.3458092e-9
+ wmax = 5.374e-7
+ aigc = 0.011492467
+ wmin = 2.674e-7
+ nfactor = 1
+ pditsd = 0
+ pditsl = 0
+ wvoff = 8.989216699999998e-9
+ cjswgd = 2.6226e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.6226e-10
+ wvsat = -0.0005775380999999999
+ wvth0 = -2.1125728e-8
+ wua1 = 1.991882e-17
+ wub1 = -2.2599817e-26
+ wuc1 = 3.0478373e-17
+ waigc = 3.9031408e-11
+ bigc = 0.001442
+ mjswgd = 0.85
+ mjswgs = 0.85
+ wwlc = 0
+ tcjswg = 0.001
+ nigbacc = 10
+ lketa = -2.0316478e-8
+ cdsc = 0
+ ijthsfwd = 0.01
+ cgbo = 0
+ xpart = 1
+ cgdl = 3.5522823e-12
+ cgdo = 5.2490134000000004e-11
+ pvfbsdoff = 0
+ xtid = 3
+ xtis = 3
+ cgsl = 3.5522823e-12
+ cgso = 5.2490134000000004e-11
+ cigc = 0.000625
+ egidl = 0.29734
+ nigbinv = 10
+ ijthsrev = 0.01
+ fprout = 300
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ fnoimod = 1
+ k2we = 5e-5
+ wtvoff = -9.0219076e-10
+ eigbinv = 1.1
+ dsub = 0.75
+ dtox = 2.7e-10
+ ppdiblc2 = 9.1292629e-19
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ pvoff = -4.585090499999998e-16
+ a0 = 0.68596391
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 55502.213
+ cf = 8.720500000000001e-11
+ cdscb = 0
+ cdscd = 0
+ ef = 1.0
+ k1 = 0.274
+ k2 = -0.024078429999999998
+ k3 = -1.8419
+ em = 1000000.0
+ ll = -1.18e-13
+ lw = 0
+ u0 = 0.012421473
+ pvsat = 1.1042156000000004e-10
+ w0 = 0
+ ua = -2.398367e-9
+ ub = 2.300703286e-18
+ uc = 8.4124236e-11
+ ud = 0
+ wk2we = 5e-12
+ capmod = 2
+ wl = 0
+ wr = 1
+ pvth0 = 8.168620000000001e-16
+ xj = 8.6e-8
+ xl = 2.33e-9
+ ww = 0
+ eta0 = 0.24044444
+ xw = 8.600000000000001e-9
+ drout = 0.56
+ etab = -0.28088889
+ wku0we = 2e-11
+ paigc = -2.2115244e-18
+ mobmod = 0
+ voffl = 0
+ cigbacc = 0.32875
+ weta0 = -1.1162667e-8
+ wetab = 2.2325333e-8
+ pkvth0we = -1.3e-19
+ lpclm = -1.0586647e-7
+ tnoimod = 0
+ cgidl = 0.22
+ vfbsdoff = 0.02
+ cigbinv = 0.006
+ laigsd = 3.4280989e-17
+ pbswd = 0.8
+ pbsws = 0.8
+ paramchk = 1
+ version = 4.5
+ wtvfbsdoff = 0
+ tempmod = 0
+ pdits = 0
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ cigsd = 0.069865
+ ltvfbsdoff = 0
+ dvt0w = 0
+ aigbacc = 0.02
+ dvt1w = 0
+ dvt2w = 0
+ ijthdfwd = 0.01
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ )

.model nch_ff_30 nmos (
+ level = 54
+ keta = -0.29566775
+ aigbinv = 0.0163
+ tnoia = 0
+ ijthdrev = 0.01
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 4.1842280000000005e-11
+ peta0 = -9.3037135e-16
+ ptvfbsdoff = 0
+ petab = -1.2138265e-15
+ kt1l = 0
+ wketa = -4.7865407e-8
+ toxref = 3e-9
+ lpdiblc2 = 8.2379047e-15
+ tpbsw = 0.0019
+ ags = 2.6744444
+ cjswd = 7.625999999999999e-11
+ cjsws = 7.625999999999999e-11
+ lint = 0
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ cjd = 0.0012620099999999998
+ cit = 0.0010507473299999999
+ cjs = 0.0012620099999999998
+ clc = 1e-7
+ cle = 0.6
+ lkt1 = -9.5950836e-9
+ bvd = 8.7
+ lkt2 = 3.8424987e-10
+ bvs = 8.7
+ lmax = 9.167e-8
+ dlc = 3.26497e-9
+ lmin = 5.567e-8
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ poxedge = 1
+ tvfbsdoff = 0.022
+ la0 = 3.9829889e-7
+ minv = -0.3
+ jsd = 6.11e-7
+ ltvoff = -2.7237524e-10
+ jss = 6.11e-7
+ lat = 0.0051856049799999995
+ lua1 = -1.2736334e-17
+ lub1 = 1.6085594e-26
+ luc1 = 1.132730421e-17
+ kt1 = -0.13273927
+ lk2 = 1.0502722e-9
+ kt2 = -0.10980467
+ llc = 0
+ binunit = 2
+ lln = 1
+ lu0 = -2.2938506000000001e-10
+ mjd = 0.26
+ lua = -7.6887484e-18
+ mjs = 0.26
+ lub = 6.3606825e-27
+ luc = -3.2720592999999998e-18
+ lud = 0
+ lwc = 0
+ ndep = 1e+18
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ lkvth0we = -2e-12
+ njs = 1.02
+ pa0 = -1.1411036e-13
+ nsd = 1e+20
+ lwlc = 0
+ pbd = 0.52
+ pat = -1.7600563e-9
+ pbs = 0.52
+ pk2 = -3.7289588e-16
+ moin = 5.1
+ pu0 = 8.3037121e-17
+ prt = 0
+ pua = 1.3044266e-23
+ pub = -1.13966382e-32
+ puc = 2.3653651e-24
+ pud = 0
+ scref = 1e-6
+ nigc = 3.083
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 7.5498293e-10
+ pigcd = 2.621
+ ub1 = -9.1820427e-19
+ uc1 = -4.319545900000001e-11
+ aigsd = 0.010772818
+ tpb = 0.0014
+ lku0we = 2.5e-11
+ wa0 = 1.7720733e-6
+ acnqsmod = 0
+ ute = -1
+ wat = 0.028542186400000003
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 7.3287188e-9
+ epsrox = 3.9
+ lvoff = -3.2711798999999994e-9
+ wlc = 0
+ wln = 1
+ wu0 = -1.6314842e-9
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -2.2058458e-16
+ wub = 1.80830997e-25
+ wuc = -3.0744792e-17
+ wud = 0
+ wwc = 0
+ noff = 2.7195
+ wwl = 0
+ wwn = 1
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ lvsat = 0.0024055243000000006
+ rbodymod = 0
+ rdsmod = 0
+ wvfbsdoff = 0
+ lvth0 = 3.4897243e-9
+ lvfbsdoff = 0
+ igbmod = 1
+ delta = 0.007595625
+ laigc = -3.0244582e-11
+ ntox = 2.029
+ pcit = -6.471760000000062e-19
+ jtsswgd = 2.3e-7
+ pclm = 1.7776553
+ jtsswgs = 2.3e-7
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ rnoia = 0
+ rnoib = 0
+ pbswgd = 0.95
+ pbswgs = 0.95
+ phin = 0.15
+ pketa = 5.3659323e-15
+ ngate = 8e+20
+ igcmod = 1
+ ngcon = 1
+ pkt1 = 5.0565068e-15
+ pkt2 = -5.9202052e-16
+ wpclm = 4.3365813e-8
+ wpdiblc2 = 1.4083642e-10
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ rbdb = 50
+ pua1 = 4.1884121e-24
+ prwb = 0
+ prwg = 0
+ pub1 = -9.7869988e-33
+ puc1 = -6.8508479999999965e-25
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ njtsswg = 9
+ rdsw = 100
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ permod = 1
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.0069717513
+ pdiblcb = -0.3
+ wkvth0we = 2e-12
+ trnqsmod = 0
+ tvoff = 0.0048149924
+ rshg = 15.6
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ voffcv = -0.16942
+ wpemod = 1
+ bigbacc = 0.002588
+ ku0we = -0.0007
+ kvth0we = 0.00018
+ beta0 = 13
+ leta0 = 2.0040249e-8
+ rgatemod = 0
+ letab = -2.6551319e-8
+ lintnoi = -1.5e-8
+ tnjtsswg = 1
+ tnom = 25
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ ppclm = -1.085908e-15
+ vtsswgs = 4.2
+ toxe = 2.3900000000000002e-9
+ toxm = 2.43e-9
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ tpbswg = 0.0009
+ dmcgt = 0
+ wags = 1.2453333e-7
+ tcjsw = 0.000357
+ wcit = -2.4019440000000024e-11
+ ptvoff = 9.0058483e-17
+ voff = -0.116438471
+ waigsd = 3.1113143e-12
+ acde = 0.4
+ vsat = 61130.093
+ wint = 0
+ bigsd = 0.00125
+ vth0 = 0.27221795299999996
+ diomod = 1
+ wkt1 = -1.0551625000000001e-7
+ wkt2 = 6.9079183e-9
+ wmax = 5.374e-7
+ aigc = 0.011842064
+ wmin = 2.674e-7
+ nfactor = 1
+ pditsd = 0
+ pditsl = 0
+ wvoff = 4.307686799999997e-9
+ cjswgd = 2.6226e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.6226e-10
+ wvsat = 0.0024248145000000006
+ wvth0 = -1.0725777100000003e-8
+ wua1 = -3.6441631e-18
+ wub1 = 2.5961869999999995e-26
+ wuc1 = -5.7163699999999976e-18
+ waigc = 4.5087747e-12
+ bigc = 0.001442
+ mjswgd = 0.85
+ mjswgs = 0.85
+ wwlc = 0
+ tcjswg = 0.001
+ nigbacc = 10
+ lketa = 8.345618e-9
+ cdsc = 0
+ ijthsfwd = 0.01
+ cgbo = 0
+ xpart = 1
+ cgdl = 3.5522823e-12
+ cgdo = 5.2490134000000004e-11
+ pvfbsdoff = 0
+ xtid = 3
+ xtis = 3
+ cgsl = 3.5522823e-12
+ cgso = 5.2490134000000004e-11
+ cigc = 0.000625
+ egidl = 0.29734
+ nigbinv = 10
+ ijthsrev = 0.01
+ fprout = 300
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ fnoimod = 1
+ k2we = 5e-5
+ wtvoff = -1.5706231e-9
+ eigbinv = 1.1
+ dsub = 0.75
+ dtox = 2.7e-10
+ ppdiblc2 = -1.1241984e-21
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ pvoff = -1.8445117999999986e-17
+ a0 = -5.7594444
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = -17682.2125
+ cf = 8.720500000000001e-11
+ cdscb = 0
+ cdscd = 0
+ ef = 1.0
+ k1 = 0.274
+ k2 = -0.069318509
+ k3 = -1.8419
+ em = 1000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.012207296000000001
+ pvsat = -1.717988000000001e-10
+ w0 = 0
+ ua = -1.7531779e-9
+ ub = 1.3845184050000002e-18
+ uc = 2.5031363e-11
+ ud = 0
+ wk2we = 5e-12
+ capmod = 2
+ wl = 0
+ wr = 1
+ pvth0 = -1.6073333999999955e-16
+ xj = 8.6e-8
+ xl = 2.33e-9
+ ww = 0
+ eta0 = 0.027250304
+ xw = 8.600000000000001e-9
+ drout = 0.56
+ etab = 0.001571952
+ wku0we = 2e-11
+ paigc = 1.0336032e-18
+ mobmod = 0
+ voffl = 0
+ cigbacc = 0.32875
+ weta0 = -1.2650991e-9
+ wetab = 3.5238381e-8
+ pkvth0we = -1.3e-19
+ lpclm = -5.0282662e-8
+ tnoimod = 0
+ cgidl = 0.22
+ vfbsdoff = 0.02
+ cigbinv = 0.006
+ pbswd = 0.8
+ pbsws = 0.8
+ paramchk = 1
+ version = 4.5
+ wtvfbsdoff = 0
+ tempmod = 0
+ pdits = 0
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ cigsd = 0.069865
+ ltvfbsdoff = 0
+ dvt0w = 0
+ aigbacc = 0.02
+ dvt1w = 0
+ dvt2w = 0
+ ijthdfwd = 0.01
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ )

.model nch_ff_31 nmos (
+ level = 54
+ nigbacc = 10
+ wvoff = 2.6164685300000083e-9
+ wvsat = 0.027479414200000003
+ wvth0 = -3.124854300000001e-8
+ ltvoff = 2.6647905e-10
+ waigc = 1.8753243e-11
+ tnom = 25
+ nigbinv = 10
+ toxe = 2.3900000000000002e-9
+ toxm = 2.43e-9
+ lketa = -2.3617222e-8
+ pvfbsdoff = 0
+ xpart = 1
+ lku0we = 2.5e-11
+ epsrox = 3.9
+ egidl = 0.29734
+ fnoimod = 1
+ pkvth0we = -1.3e-19
+ wags = 1.2453333e-7
+ rdsmod = 0
+ eigbinv = 1.1
+ wcit = 6.4454534e-10
+ igbmod = 1
+ voff = -0.07382279000000001
+ acde = 0.4
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ vfbsdoff = 0.02
+ vsat = 36969.44000000001
+ pbswgd = 0.95
+ pbswgs = 0.95
+ wint = 0
+ vth0 = 0.25339229
+ wkt1 = -1.09856149e-7
+ wkt2 = -2.0876247e-8
+ wmax = 5.374e-7
+ igcmod = 1
+ aigc = 0.011696193
+ wmin = 2.674e-7
+ paramchk = 1
+ cigbacc = 0.32875
+ wua1 = -1.1132499e-16
+ wub1 = -4.4080979999999945e-26
+ wuc1 = 1.6593491000000002e-16
+ pvoff = 7.964544000000045e-17
+ bigc = 0.001442
+ cdscb = 0
+ cdscd = 0
+ tnoimod = 0
+ wwlc = 0
+ pvsat = -1.624968e-9
+ wk2we = 5e-12
+ pvth0 = 1.0295868e-15
+ drout = 0.56
+ paigsd = 1.7624612e-23
+ cdsc = 0
+ paigc = 2.0742404e-19
+ cigbinv = 0.006
+ ijthdfwd = 0.01
+ cgbo = 0
+ cgdl = 3.5522823e-12
+ cgdo = 5.2490134000000004e-11
+ xtid = 3
+ xtis = 3
+ voffl = 0
+ cgsl = 3.5522823e-12
+ cgso = 5.2490134000000004e-11
+ cigc = 0.000625
+ permod = 1
+ weta0 = -1.2005104e-7
+ wetab = 5.6750807e-8
+ lpclm = 5.458214e-8
+ version = 4.5
+ tempmod = 0
+ ijthdrev = 0.01
+ cgidl = 0.22
+ voffcv = -0.16942
+ wpemod = 1
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ aigbacc = 0.02
+ pbswd = 0.8
+ pbsws = 0.8
+ k2we = 5e-5
+ dsub = 0.75
+ dtox = 2.7e-10
+ aigbinv = 0.0163
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ pdits = 0
+ cigsd = 0.069865
+ lkvth0we = -2e-12
+ eta0 = 1.0176617
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ etab = -1.3959412
+ tpbswg = 0.0009
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ acnqsmod = 0
+ tnoia = 0
+ ptvoff = -4.401556e-18
+ poxedge = 1
+ rbodymod = 0
+ ags = 2.6744444
+ waigsd = 3.1110104e-12
+ peta0 = 5.9592132e-15
+ cjd = 0.0012620099999999998
+ cit = -0.0056353599
+ cjs = 0.0012620099999999998
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ petab = -2.4615472e-15
+ dlc = 3.26497e-9
+ binunit = 2
+ wketa = -5.877032e-8
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ diomod = 1
+ tpbsw = 0.0019
+ cjswd = 7.625999999999999e-11
+ cjsws = 7.625999999999999e-11
+ mjswd = 0.11
+ pditsd = 0
+ pditsl = 0
+ mjsws = 0.11
+ agidl = 9.41e-8
+ cjswgd = 2.6226e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.6226e-10
+ la0 = -1.4097724e-8
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = 0.0024085122999999986
+ kt1 = -0.23060700999999997
+ lk2 = 7.4338958e-10
+ kt2 = -0.14677127
+ llc = 0
+ lln = 1
+ lu0 = 4.6598268e-10
+ mjd = 0.26
+ lua = 6.4763643e-17
+ mjs = 0.26
+ lub = -2.3096342000000002e-26
+ luc = -1.0931136000000001e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = -1.7333804e-13
+ nsd = 1e+20
+ pbd = 0.52
+ pat = -2.2283547099999997e-9
+ tvfbsdoff = 0.022
+ pbs = 0.52
+ pk2 = -1.0803308e-16
+ wpdiblc2 = 1.4081704e-10
+ pu0 = -3.5315192999999994e-17
+ prt = 0
+ pua = -2.1774501e-24
+ pub = -5.473259300000002e-33
+ puc = 4.761497700000001e-24
+ pud = 0
+ mjswgd = 0.85
+ mjswgs = 0.85
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 1.4910078e-9
+ ub1 = -1.2882590799999998e-18
+ uc1 = -4.0168785999999996e-10
+ tpb = 0.0014
+ tcjswg = 0.001
+ wa0 = 2.7932403e-6
+ ute = -1
+ wat = 0.03661635459999999
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 2.7621189e-9
+ wlc = 0
+ wln = 1
+ wu0 = 4.090729e-10
+ jtsswgd = 2.3e-7
+ xgl = -1.09e-8
+ jtsswgs = 2.3e-7
+ xgw = 0
+ wua = 4.1858808e-17
+ wub = 7.870378029999999e-26
+ wuc = -7.2057435e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ scref = 1e-6
+ pigcd = 2.621
+ aigsd = 0.010772819
+ keta = 0.2554158
+ lvoff = -5.742889800000002e-9
+ wkvth0we = 2e-12
+ wvfbsdoff = 0
+ lvsat = 0.00380682957
+ lvfbsdoff = 0
+ lvth0 = 4.581610599999999e-9
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 4.2963728999999995e-10
+ trnqsmod = 0
+ delta = 0.007595625
+ laigc = -2.1784105e-11
+ kt1l = 0
+ fprout = 300
+ xrcrg1 = 12
+ xrcrg2 = 1
+ rnoia = 0
+ rnoib = 0
+ lint = 0
+ njtsswg = 9
+ lkt1 = -3.918750599999999e-9
+ lkt2 = 2.528313e-9
+ pketa = 5.998417e-15
+ ngate = 8e+20
+ lmax = 5.567e-8
+ lmin = 4.667e-8
+ wtvoff = 5.799816e-11
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ ngcon = 1
+ wpclm = 2.4669208e-7
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ ckappad = 0.6
+ ckappas = 0.6
+ rgatemod = 0
+ gbmin = 1e-12
+ pdiblc1 = 0
+ pdiblc2 = 0.0069718933
+ pdiblcb = -0.3
+ tnjtsswg = 1
+ minv = -0.3
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ lua1 = -5.5425775e-17
+ lub1 = 3.7548779999999994e-26
+ luc1 = 3.2119863e-17
+ capmod = 2
+ ndep = 1e+18
+ wku0we = 2e-11
+ lwlc = 0
+ moin = 5.1
+ mobmod = 0
+ nigc = 3.083
+ bigbacc = 0.002588
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ kvth0we = 0.00018
+ wtvfbsdoff = 0
+ lintnoi = -1.5e-8
+ bigbinv = 0.004953
+ tvoff = -0.0044755986
+ ntox = 2.029
+ vtsswgd = 4.2
+ pcit = -3.9423707e-17
+ vtsswgs = 4.2
+ pclm = -0.030358553
+ laigsd = -6.385731e-17
+ xjbvd = 1
+ a0 = 1.350842
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ xjbvs = 1
+ lk2we = -1.5e-12
+ at = 30198.703000000005
+ cf = 8.720500000000001e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = -0.064027428
+ k3 = -1.8419
+ em = 1000000.0
+ ltvfbsdoff = 0
+ ll = 0
+ lw = 0
+ u0 = 0.00021819504690000002
+ w0 = 0
+ ua = -3.002357e-9
+ ub = 1.89239813e-18
+ uc = 1.5708441000000004e-10
+ ud = 0
+ phin = 0.15
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 2.33e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ pkt1 = 5.308216660000001e-15
+ pkt2 = 1.019461e-15
+ ku0we = -0.0007
+ beta0 = 13
+ leta0 = -3.7403611e-8
+ letab = 5.4504443e-8
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ ppclm = -1.2878832e-14
+ rbdb = 50
+ pua1 = 1.04339e-23
+ prwb = 0
+ prwg = 0
+ pub1 = -5.7245160000000007e-33
+ puc1 = -1.0640858600000001e-23
+ rbpb = 50
+ rbpd = 50
+ dlcig = 2.5e-9
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ bgidl = 2320000000.0
+ ptvfbsdoff = 0
+ rdsw = 100
+ ijthsfwd = 0.01
+ nfactor = 1
+ dmcgt = 0
+ tcjsw = 0.000357
+ ijthsrev = 0.01
+ toxref = 3e-9
+ rshg = 15.6
+ bigsd = 0.00125
+ )

.model nch_ff_32 nmos (
+ level = 54
+ eta0 = -0.25440451
+ etab = -0.81370191
+ scref = 1e-6
+ lku0we = 2.5e-11
+ pigcd = 2.621
+ epsrox = 3.9
+ aigsd = 0.010772817
+ njtsswg = 9
+ lvoff = -6.3467068e-9
+ rdsmod = 0
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ igbmod = 1
+ lvsat = -0.0002660245999999999
+ ckappad = 0.6
+ ckappas = 0.6
+ lvth0 = -2.316650100000001e-9
+ pdiblc1 = 0
+ pdiblc2 = 0.0069718933
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ pdiblcb = -0.3
+ delta = 0.007595625
+ laigc = 9.707156e-12
+ pbswgd = 0.95
+ pbswgs = 0.95
+ rnoia = 0
+ rnoib = 0
+ igcmod = 1
+ pketa = -6.053668000000001e-15
+ ngate = 8e+20
+ ngcon = 1
+ wpclm = 1.6305740000000013e-7
+ bigbacc = 0.002588
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ kvth0we = 0.00018
+ paigsd = -1.2154906e-23
+ lintnoi = -1.5e-8
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ ijthsfwd = 0.01
+ permod = 1
+ keta = -0.59506219
+ ijthsrev = 0.01
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 7.960899999999999e-10
+ tvoff = 0.0034020192
+ kt1l = 0
+ voffcv = -0.16942
+ wpemod = 1
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ lint = 0
+ lkt1 = -1.2951426000000001e-8
+ lkt2 = 1.0897551e-9
+ lmax = 4.667e-8
+ lmin = 3.6e-8
+ ku0we = -0.0007
+ nfactor = 1
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ beta0 = 13
+ leta0 = 2.4927632200000002e-8
+ letab = 2.5974719e-8
+ minv = -0.3
+ lua1 = 7.6118385e-17
+ lub1 = -1.1028845e-25
+ luc1 = -3.7246243e-17
+ ppclm = -8.780734400000002e-15
+ ndep = 1e+18
+ dlcig = 2.5e-9
+ lwlc = 0
+ tpbswg = 0.0009
+ bgidl = 2320000000.0
+ moin = 5.1
+ nigc = 3.083
+ nigbacc = 10
+ dmcgt = 0
+ pkvth0we = -1.3e-19
+ noff = 2.7195
+ tcjsw = 0.000357
+ ptvoff = -5.392468e-18
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ waigsd = 3.1116181e-12
+ nigbinv = 10
+ diomod = 1
+ ntox = 2.029
+ pcit = -8.631339099999999e-17
+ vfbsdoff = 0.02
+ pclm = 1.46768105
+ bigsd = 0.00125
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 2.6226e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.6226e-10
+ phin = 0.15
+ wvoff = 6.255152000000001e-9
+ paramchk = 1
+ pkt1 = 1.6745505000000003e-15
+ pkt2 = -4.1883975e-17
+ wvsat = -0.019571025999999995
+ wvth0 = -1.5130829e-8
+ fnoimod = 1
+ mjswgd = 0.85
+ mjswgs = 0.85
+ eigbinv = 1.1
+ waigc = 7.6854687e-11
+ tcjswg = 0.001
+ rbdb = 50
+ pua1 = -2.7889543e-23
+ prwb = 0
+ prwg = 0
+ pub1 = 4.0160499e-32
+ puc1 = 1.2190153e-23
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ pvfbsdoff = 0
+ lketa = 1.80561909e-8
+ ijthdfwd = 0.01
+ rdsw = 100
+ xpart = 1
+ egidl = 0.29734
+ cigbacc = 0.32875
+ ijthdrev = 0.01
+ fprout = 300
+ rshg = 15.6
+ xrcrg1 = 12
+ xrcrg2 = 1
+ tnoimod = 0
+ cigbinv = 0.006
+ wtvoff = 7.822084e-11
+ pvoff = -9.865003999999993e-17
+ version = 4.5
+ capmod = 2
+ tnom = 25
+ cdscb = 0
+ cdscd = 0
+ tempmod = 0
+ toxe = 2.3900000000000002e-9
+ toxm = 2.43e-9
+ pvsat = 6.805058200000002e-10
+ wku0we = 2e-11
+ lkvth0we = -2e-12
+ wk2we = 5e-12
+ pvth0 = 2.398146000000002e-16
+ drout = 0.56
+ mobmod = 0
+ wtvfbsdoff = 0
+ paigc = -2.6395467e-18
+ aigbacc = 0.02
+ voffl = 0
+ acnqsmod = 0
+ ltvfbsdoff = 0
+ weta0 = 8.5615058e-8
+ wetab = 2.2270081e-8
+ wags = 1.2453333e-7
+ lpclm = -1.8821805999999992e-8
+ wcit = 1.6014509e-9
+ rbodymod = 0
+ aigbinv = 0.0163
+ voff = -0.061499972999999986
+ cgidl = 0.22
+ acde = 0.4
+ laigsd = 4.4039511e-17
+ vsat = 120089.242
+ wint = 0
+ vth0 = 0.39417297100000004
+ wkt1 = -3.5699569999999984e-8
+ wkt2 = 7.8385579e-10
+ wmax = 5.374e-7
+ aigc = 0.011053515
+ wmin = 2.674e-7
+ pbswd = 0.8
+ pbsws = 0.8
+ ptvfbsdoff = 0
+ wpdiblc2 = 1.4081704e-10
+ wua1 = 6.7078609e-16
+ wub1 = -9.805099000000002e-25
+ wuc1 = -3.0000411e-16
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ poxedge = 1
+ bigc = 0.001442
+ pdits = 0
+ wwlc = 0
+ cigsd = 0.069865
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ binunit = 2
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.5522823e-12
+ cgdo = 5.2490134000000004e-11
+ xtid = 3
+ xtis = 3
+ ags = 2.6744444
+ cgsl = 3.5522823e-12
+ pk2we = -1e-19
+ cgso = 5.2490134000000004e-11
+ cigc = 0.000625
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ a0 = 10.55945905
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 152950.757
+ cf = 8.720500000000001e-11
+ cjd = 0.0012620099999999998
+ cit = -0.0131140508
+ cjs = 0.0012620099999999998
+ clc = 1e-7
+ ef = 1.0
+ k1 = 0.274
+ cle = 0.6
+ k2 = 0.037127322
+ k3 = -1.8419
+ em = 1000000.0
+ bvd = 8.7
+ bvs = 8.7
+ ll = 0
+ lw = 0
+ dlc = 3.26497e-9
+ u0 = 0.006973015400000001
+ w0 = 0
+ k3b = 1.9326
+ ua = -1.7148580999999998e-9
+ ub = 1.250859149999999e-18
+ uc = 5.4381728e-10
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 2.33e-9
+ dwb = 0
+ ww = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ xw = 8.600000000000001e-9
+ wkvth0we = 2e-12
+ tnoia = 0
+ toxref = 3e-9
+ peta0 = -4.1184253e-15
+ la0 = -4.65319969e-7
+ trnqsmod = 0
+ petab = -7.719916e-16
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.00360633488
+ kt1 = -0.04626677999999999
+ lk2 = -4.2131932e-9
+ kt2 = -0.11741295
+ wketa = 1.87190595e-7
+ llc = 0
+ lln = 1
+ lu0 = 1.3499632e-10
+ mjd = 0.26
+ lua = 1.6761980000000137e-18
+ mjs = 0.26
+ lub = 8.339062399999967e-27
+ luc = -2.98810456e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ tpbsw = 0.0019
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 9.065128000000001e-14
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 1.15850572e-9
+ pbs = 0.52
+ pk2 = 5.9540883e-16
+ cjswd = 7.625999999999999e-11
+ cjsws = 7.625999999999999e-11
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ pu0 = -8.848033e-17
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ prt = 0
+ pua = -1.6092489999999997e-23
+ pub = 1.5276544400000003e-32
+ puc = 5.518326299999999e-24
+ pud = 0
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = -1.1935669e-9
+ ub1 = 1.7288272299999998e-18
+ uc1 = 1.0139469700000001e-9
+ tpb = 0.0014
+ k2we = 5e-5
+ wa0 = -2.59429679e-6
+ tvfbsdoff = 0.022
+ ute = -1
+ wat = -0.0325032315
+ dsub = 0.75
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -1.1593839e-8
+ ltvoff = -1.1952424e-10
+ dtox = 2.7e-10
+ wlc = 0
+ wln = 1
+ rgatemod = 0
+ wu0 = 1.4940757e-9
+ xgl = -1.09e-8
+ xgw = 0
+ wua = 3.2583921000000013e-16
+ wub = -3.447615700000002e-25
+ wuc = -8.750290400000002e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ tnjtsswg = 1
+ )

.model nch_ff_33 nmos (
+ level = 54
+ rbodymod = 0
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ version = 4.5
+ pbswgd = 0.95
+ pbswgs = 0.95
+ ntox = 2.029
+ pcit = -1.5e-17
+ pclm = 1.8851852
+ tempmod = 0
+ igcmod = 1
+ phin = 0.15
+ aigbacc = 0.02
+ pkt1 = -5e-17
+ wpdiblc2 = -2.9834e-10
+ pvoff = 0
+ cdscb = 0
+ cdscd = 0
+ pvsat = -1.8e-11
+ aigbinv = 0.0163
+ rbdb = 50
+ prwb = 0
+ prwg = 0
+ pub1 = 0
+ wk2we = 5e-12
+ pvth0 = -2.3e-16
+ drout = 0.56
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ rdsw = 100
+ permod = 1
+ voffl = 0
+ weta0 = 0
+ wkvth0we = 2e-12
+ cgidl = 0.22
+ trnqsmod = 0
+ voffcv = -0.16942
+ wpemod = 1
+ poxedge = 1
+ rshg = 15.6
+ binunit = 2
+ pbswd = 0.8
+ pbsws = 0.8
+ rgatemod = 0
+ tnjtsswg = 1
+ tnom = 25
+ pdits = 0
+ ags = 0.6188259300000001
+ cigsd = 0.069865
+ toxe = 2.3900000000000002e-9
+ toxm = 2.43e-9
+ tpbswg = 0.0009
+ cjd = 0.0012620099999999998
+ dvt0w = 0
+ cit = 0.002342713
+ dvt1w = 0
+ cjs = 0.0012620099999999998
+ clc = 1e-7
+ cle = 0.6
+ dvt2w = 0
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 9.8024918e-9
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ jtsswgd = 2.3e-7
+ pk2we = -1e-19
+ jtsswgs = 2.3e-7
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ la0 = 0
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.0001
+ kt1 = -0.21767878
+ kt2 = -0.055117852
+ ptvoff = 0
+ llc = 0
+ lln = 1
+ lu0 = 6e-12
+ wags = 1.9944440000000004e-9
+ mjd = 0.26
+ mjs = 0.26
+ lub = 0
+ lud = 0
+ lwc = 0
+ waigsd = 3.1789128e-12
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 0
+ tnoia = 0
+ nsd = 1e+20
+ pbd = 0.52
+ pat = -2.8e-11
+ wcit = -2.0566928e-10
+ pbs = 0.52
+ pu0 = 2e-18
+ prt = 0
+ pub = 0
+ pud = 0
+ peta0 = 0
+ diomod = 1
+ voff = -0.095952978
+ acde = 0.4
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 9.5347726e-10
+ wketa = -1.1490089e-9
+ ub1 = -5.3850981e-19
+ uc1 = -6.0041111e-11
+ tpb = 0.0014
+ tpbsw = 0.0019
+ pditsd = 0
+ pditsl = 0
+ vsat = 84306.193
+ wa0 = 0
+ cjswgd = 2.6226e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.6226e-10
+ wint = 0
+ ute = -1
+ wat = 0
+ vth0 = 0.28469411
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 3.0219344e-9
+ cjswd = 7.625999999999999e-11
+ cjsws = 7.625999999999999e-11
+ wlc = 0
+ wln = 1
+ wu0 = -1.2693332999999998e-11
+ wkt1 = -2.89145825e-9
+ wkt2 = 1.0235511e-10
+ xgl = -1.09e-8
+ mjswd = 0.11
+ xgw = 0
+ mjsws = 0.11
+ wua = -1.6467997e-17
+ wub = 3.619626e-26
+ wuc = -1.4955111e-18
+ wud = 0
+ agidl = 9.41e-8
+ wmax = 2.674e-7
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ aigc = 0.01181895
+ wmin = 1.08e-7
+ tvfbsdoff = 0.022
+ njtsswg = 9
+ mjswgd = 0.85
+ mjswgs = 0.85
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ wua1 = -3.1223388e-18
+ wub1 = 2.0807554e-26
+ wuc1 = 8.1864667e-18
+ tcjswg = 0.001
+ bigc = 0.001442
+ ckappad = 0.6
+ ckappas = 0.6
+ wwlc = 0
+ pdiblc1 = 0
+ pdiblc2 = 0.023869018
+ pdiblcb = -0.3
+ scref = 1e-6
+ cdsc = 0
+ ijthsfwd = 0.01
+ cgbo = 0
+ cgdl = 3.5522823e-12
+ cgdo = 5.2490134000000004e-11
+ xtid = 3
+ xtis = 3
+ pigcd = 2.621
+ aigsd = 0.010772573
+ cgsl = 3.5522823e-12
+ cgso = 5.2490134000000004e-11
+ cigc = 0.000625
+ lvoff = -2e-11
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ bigbacc = 0.002588
+ lvsat = -0.0003
+ lvth0 = -1e-10
+ fprout = 300
+ ijthsrev = 0.01
+ delta = 0.007595625
+ xrcrg1 = 12
+ xrcrg2 = 1
+ kvth0we = 0.00018
+ rnoia = 0
+ rnoib = 0
+ lintnoi = -1.5e-8
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ wtvoff = 2.5061202e-10
+ ngate = 8e+20
+ wtvfbsdoff = 0
+ ngcon = 1
+ wpclm = -9.7111111e-9
+ k2we = 5e-5
+ dsub = 0.75
+ dtox = 2.7e-10
+ gbmin = 1e-12
+ capmod = 2
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ ltvfbsdoff = 0
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ wku0we = 2e-11
+ mobmod = 0
+ eta0 = 0.2
+ etab = -0.2
+ pkvth0we = -1.3e-19
+ nfactor = 1
+ ptvfbsdoff = 0
+ tvoff = 0.00085486634
+ vfbsdoff = 0.02
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ paramchk = 1
+ nigbacc = 10
+ ku0we = -0.0007
+ beta0 = 13
+ leta0 = 0
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ dlcig = 2.5e-9
+ nigbinv = 10
+ bgidl = 2320000000.0
+ ijthdfwd = 0.01
+ keta = -0.021050128
+ dmcgt = 0
+ tcjsw = 0.000357
+ toxref = 3e-9
+ ijthdrev = 0.01
+ fnoimod = 1
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = -1e-11
+ eigbinv = 1.1
+ kt1l = 0
+ bigsd = 0.00125
+ lint = 6.5375218e-9
+ lkt1 = -1.1e-9
+ wvoff = 2.9681533e-9
+ lmax = 2.001e-5
+ lmin = 9.00077e-6
+ ltvoff = 0
+ lpe0 = 9.2e-8
+ wvsat = 0.002322956
+ lpeb = 2.5e-7
+ wvth0 = -7.551373900000001e-9
+ a0 = 3.5
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 200000
+ cf = 8.720500000000001e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.013956400999999998
+ k3 = -1.8419
+ em = 1000000.0
+ minv = -0.3
+ waigc = 1.7818122e-11
+ ll = 0
+ lw = 0
+ u0 = 0.012535556000000002
+ w0 = 0
+ lub1 = 0
+ ua = -2.0911548e-9
+ ub = 2.2368542e-18
+ uc = 5.8018519e-11
+ ud = 0
+ cigbacc = 0.32875
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 2.33e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ ndep = 1e+18
+ lkvth0we = -2e-12
+ pvfbsdoff = 0
+ lwlc = 0
+ moin = 5.1
+ lku0we = 2.5e-11
+ tnoimod = 0
+ epsrox = 3.9
+ xpart = 1
+ nigc = 3.083
+ cigbinv = 0.006
+ acnqsmod = 0
+ rdsmod = 0
+ egidl = 0.29734
+ igbmod = 1
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ )

.model nch_ff_34 nmos (
+ level = 54
+ paramchk = 1
+ wpclm = -9.7111111e-9
+ gbmin = 1e-12
+ wua1 = -1.7574281e-19
+ wub1 = 1.7597088e-26
+ wuc1 = 8.3134424e-18
+ jswgd = 1.28e-13
+ nfactor = 1
+ jswgs = 1.28e-13
+ paigsd = -3.8370159e-23
+ bigc = 0.001442
+ wwlc = 0
+ permod = 1
+ cdsc = 0
+ ijthdfwd = 0.01
+ cgbo = 0
+ cgdl = 3.5522823e-12
+ cgdo = 5.2490134000000004e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.5522823e-12
+ cgso = 5.2490134000000004e-11
+ cigc = 0.000625
+ nigbacc = 10
+ ijthdrev = 0.01
+ voffcv = -0.16942
+ wpemod = 1
+ tvoff = 0.00082419905
+ lpdiblc2 = -9.2950492e-9
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ nigbinv = 10
+ k2we = 5e-5
+ ku0we = -0.0007
+ beta0 = 13
+ dsub = 0.75
+ leta0 = 0
+ dtox = 2.7e-10
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ tpbswg = 0.0009
+ fnoimod = 1
+ lkvth0we = -2e-12
+ eigbinv = 1.1
+ dlcig = 2.5e-9
+ eta0 = 0.2
+ bgidl = 2320000000.0
+ etab = -0.2
+ acnqsmod = 0
+ ptvoff = -2.3727895e-16
+ waigsd = 3.1789171e-12
+ dmcgt = 0
+ tcjsw = 0.000357
+ rbodymod = 0
+ diomod = 1
+ cigbacc = 0.32875
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 2.6226e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.6226e-10
+ bigsd = 0.00125
+ tnoimod = 0
+ wvoff = 3.141381e-9
+ mjswgd = 0.85
+ mjswgs = 0.85
+ cigbinv = 0.006
+ wvsat = 0.002322956
+ wvth0 = -7.7363659e-9
+ wpdiblc2 = -6.4961636e-10
+ tcjswg = 0.001
+ waigc = 1.8291238e-11
+ pvfbsdoff = 0
+ version = 4.5
+ lketa = -2.7750915e-8
+ tempmod = 0
+ xpart = 1
+ egidl = 0.29734
+ aigbacc = 0.02
+ keta = -0.017963263
+ wkvth0we = 2e-12
+ wtvfbsdoff = 0
+ fprout = 300
+ lags = 4.3821463e-7
+ xrcrg1 = 12
+ xrcrg2 = 1
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = -1.9265105499999997e-11
+ trnqsmod = 0
+ kt1l = 0
+ ltvfbsdoff = 0
+ aigbinv = 0.0163
+ wtvoff = 2.7700567e-10
+ lint = 6.5375218e-9
+ lkt1 = -8.9918468e-8
+ lkt2 = -1.6837724e-8
+ lmax = 9.00077e-6
+ lmin = 9.0075e-7
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ capmod = 2
+ rgatemod = 0
+ pvoff = -1.5573172e-15
+ tnjtsswg = 1
+ wku0we = 2e-11
+ minv = -0.3
+ lua1 = -7.4262143e-17
+ lub1 = -1.4158035e-25
+ luc1 = 6.2830403e-17
+ cdscb = 0
+ cdscd = 0
+ mobmod = 0
+ pvsat = -1.8e-11
+ ndep = 1e+18
+ wk2we = 5e-12
+ pvth0 = 1.4330782e-15
+ ptvfbsdoff = 0
+ drout = 0.56
+ lwlc = 0
+ poxedge = 1
+ moin = 5.1
+ paigc = -4.2533129e-18
+ nigc = 3.083
+ voffl = 0
+ binunit = 2
+ weta0 = 0
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ laigsd = 3.3658034e-16
+ pags = 5.2134206e-15
+ cgidl = 0.22
+ ntox = 2.029
+ pcit = 6.488187400000001e-17
+ pclm = 1.8851852
+ phin = 0.15
+ pbswd = 0.8
+ pbsws = 0.8
+ ags = 0.5700812500000001
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ pkt1 = -4.1416964000000005e-16
+ pkt2 = -1.7740443e-15
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ cjd = 0.0012620099999999998
+ cit = 0.0023437436
+ cjs = 0.0012620099999999998
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 9.8024918e-9
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ pdits = 0
+ cigsd = 0.069865
+ rbdb = 50
+ pua1 = -2.6489898e-23
+ prwb = 0
+ prwg = 0
+ pub1 = 2.886209e-32
+ puc1 = -1.1415122e-24
+ dvt0w = 0
+ la0 = -1.6207075e-6
+ dvt1w = 0
+ dvt2w = 0
+ rbpb = 50
+ rbpd = 50
+ jsd = 6.11e-7
+ rbps = 50
+ jss = 6.11e-7
+ lat = -0.043322769000000004
+ rbsb = 50
+ pvag = 1.2
+ kt1 = -0.20779908
+ lk2 = -1.5849432e-8
+ kt2 = -0.053244913
+ llc = 0
+ lln = 1
+ lu0 = -1.6732432e-9
+ mjd = 0.26
+ lua = -1.2813977e-16
+ mjs = 0.26
+ lub = -8.5009677e-26
+ luc = -2.2547224e-17
+ lud = 0
+ ijthsfwd = 0.01
+ lwc = 0
+ lwl = 0
+ rdsw = 100
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 3.8370159e-14
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 3.9624965e-9
+ pbs = 0.52
+ pk2 = -8.7965669e-16
+ pk2we = -1e-19
+ pu0 = 1.999999999998372e-18
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ prt = 0
+ pua = -3.3674591e-24
+ pub = -4.9159389e-33
+ puc = 2.3789498e-24
+ pud = 0
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 9.6173779e-10
+ ub1 = -5.2276116e-19
+ uc1 = -6.7030033e-11
+ njtsswg = 9
+ tpb = 0.0014
+ toxref = 3e-9
+ wa0 = -4.2680933e-9
+ tnoia = 0
+ ute = -1
+ wat = -0.0004438817
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 3.1197827e-9
+ wlc = 0
+ wln = 1
+ wu0 = -1.2693332999999998e-11
+ ijthsrev = 0.01
+ xgl = -1.09e-8
+ xtsswgd = 0.18
+ xgw = 0
+ xtsswgs = 0.18
+ wua = -1.6093419e-17
+ wub = 3.6743083e-26
+ wuc = -1.7601329e-18
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ peta0 = 0
+ wketa = -1.4921751e-9
+ ckappad = 0.6
+ ckappas = 0.6
+ rshg = 15.6
+ pdiblc1 = 0
+ pdiblc2 = 0.02490295
+ tpbsw = 0.0019
+ pdiblcb = -0.3
+ cjswd = 7.625999999999999e-11
+ cjsws = 7.625999999999999e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ tvfbsdoff = 0.022
+ ltvoff = 2.7569894e-10
+ ppdiblc2 = 3.1579745e-15
+ bigbacc = 0.002588
+ tnom = 25
+ toxe = 2.3900000000000002e-9
+ toxm = 2.43e-9
+ kvth0we = 0.00018
+ lku0we = 2.5e-11
+ epsrox = 3.9
+ scref = 1e-6
+ lintnoi = -1.5e-8
+ pigcd = 2.621
+ bigbinv = 0.004953
+ aigsd = 0.010772573
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ rdsmod = 0
+ wvfbsdoff = 0
+ igbmod = 1
+ lvoff = -1.4758881e-8
+ lvfbsdoff = 0
+ pkvth0we = -1.3e-19
+ wags = 1.4145310000000025e-9
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ lvsat = -0.0003
+ wcit = -2.1455490999999998e-10
+ lvth0 = 5.651542e-8
+ pbswgd = 0.95
+ pbswgs = 0.95
+ voff = -0.094313503
+ delta = 0.007595625
+ laigc = -1.6452737e-10
+ acde = 0.4
+ a0 = 3.6802789
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ vfbsdoff = 0.02
+ igcmod = 1
+ at = 204807.87
+ cf = 8.720500000000001e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.015719407999999997
+ k3 = -1.8419
+ em = 1000000.0
+ rnoia = 0
+ rnoib = 0
+ ll = 0
+ lw = 0
+ vsat = 84306.193
+ u0 = 0.012722346
+ w0 = 0
+ wint = 0
+ ua = -2.0769012e-9
+ ub = 2.2463102e-18
+ uc = 6.0526552e-11
+ ud = 0
+ vth0 = 0.27839651
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 2.33e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ wkt1 = -2.85094995e-9
+ wkt2 = 2.996904e-10
+ wmax = 2.674e-7
+ aigc = 0.011837251
+ wmin = 1.08e-7
+ pketa = 3.0850638e-15
+ ngate = 8e+20
+ ngcon = 1
+ )

.model nch_ff_35 nmos (
+ level = 54
+ a0 = 2.7573663
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ voffl = 0
+ at = 225908.74
+ cf = 8.720500000000001e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.008686581
+ k3 = -1.8419
+ em = 1000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.01231229
+ w0 = 0
+ ua = -2.2251639e-9
+ ub = 2.3450974e-18
+ uc = 3.6825844e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 2.33e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ weta0 = 0
+ keta = -0.063873893
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ voffcv = -0.16942
+ wpemod = 1
+ lags = -4.2829945e-7
+ ijthsrev = 0.01
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ cgidl = 0.22
+ lcit = -6.2890204e-10
+ kt1l = 0
+ ags = 1.5436926
+ cjd = 0.0012620099999999998
+ cit = 0.0030287289
+ cjs = 0.0012620099999999998
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 9.8024918e-9
+ k3b = 1.9326
+ lint = 6.5375218e-9
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ lkt1 = 4.7951427000000004e-8
+ lkt2 = -1.4519819e-8
+ pbswd = 0.8
+ pbsws = 0.8
+ lmax = 9.0075e-7
+ lmin = 4.5075e-7
+ lpe0 = 9.2e-8
+ la0 = -7.9931523e-7
+ lpeb = 2.5e-7
+ jsd = 6.11e-7
+ ppdiblc2 = -1.3141262e-15
+ jss = 6.11e-7
+ lat = -0.062102545
+ kt1 = -0.36270908
+ lk2 = -9.5902228e-9
+ kt2 = -0.0558493
+ llc = 0
+ lln = 1
+ lu0 = -1.3082934e-9
+ njtsswg = 9
+ mjd = 0.26
+ lua = 3.8140531e-18
+ mjs = 0.26
+ lub = -1.7293024e-25
+ luc = -1.4535934e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ tpbswg = 0.0009
+ njd = 1.02
+ minv = -0.3
+ njs = 1.02
+ pa0 = -6.7606598e-14
+ lua1 = -1.6437259e-16
+ lub1 = 2.2818043e-26
+ nsd = 1e+20
+ pdits = 0
+ luc1 = 5.6450349e-17
+ pbd = 0.52
+ pat = 1.6752657e-9
+ pbs = 0.52
+ pk2 = -2.3173279e-16
+ cigsd = 0.069865
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ pu0 = 1.09578742e-17
+ prt = 0
+ ndep = 1e+18
+ pua = -1.9061799e-24
+ pub = 1.3958464e-33
+ puc = -1.352132e-24
+ pud = 0
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ lwlc = 0
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 1.0629855e-9
+ ckappad = 0.6
+ ub1 = -7.0747845e-19
+ moin = 5.1
+ uc1 = -5.9861432e-11
+ ckappas = 0.6
+ tpb = 0.0014
+ pdiblc1 = 0
+ pdiblc2 = 0.01020022
+ pdiblcb = -0.3
+ wa0 = 1.1480691e-7
+ ute = -1
+ nigc = 3.083
+ wat = 0.0021260405
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 2.3917793e-9
+ wlc = 0
+ pk2we = -1e-19
+ ptvoff = -4.8469984e-16
+ wln = 1
+ wu0 = -2.2758359999999998e-11
+ xgl = -1.09e-8
+ dvtp0 = 4e-7
+ xgw = 0
+ dvtp1 = 0.01
+ wua = -1.7735306e-17
+ wub = 2.9651178e-26
+ wuc = 2.4320938e-18
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ waigsd = 3.178874e-12
+ pkvth0we = -1.3e-19
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ tnoia = 0
+ diomod = 1
+ bigbacc = 0.002588
+ peta0 = 0
+ pags = -9.2425378e-15
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 2.6226e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.6226e-10
+ wketa = 5.5022601e-9
+ vfbsdoff = 0.02
+ ntox = 2.029
+ pcit = 1.438079e-16
+ pclm = 1.8851852
+ tpbsw = 0.0019
+ kvth0we = 0.00018
+ cjswd = 7.625999999999999e-11
+ cjsws = 7.625999999999999e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ phin = 0.15
+ tvfbsdoff = 0.022
+ lintnoi = -1.5e-8
+ bigbinv = 0.004953
+ mjswgd = 0.85
+ mjswgs = 0.85
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ paramchk = 1
+ pkt1 = -1.3261355e-14
+ pkt2 = 1.7857928e-15
+ tcjswg = 0.001
+ wtvfbsdoff = 0
+ rbdb = 50
+ pua1 = 3.1539092e-23
+ prwb = 0
+ prwg = 0
+ pub1 = -3.1533886e-32
+ puc1 = -7.798421e-24
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ scref = 1e-6
+ ijthdfwd = 0.01
+ rdsw = 100
+ pigcd = 2.621
+ aigsd = 0.010772573
+ ltvfbsdoff = 0
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ lvoff = -2.8476354e-8
+ fprout = 300
+ lvsat = -0.0003
+ xrcrg1 = 12
+ xrcrg2 = 1
+ lvth0 = 1.8654805999999998e-8
+ ijthdrev = 0.01
+ delta = 0.007595625
+ nfactor = 1
+ laigc = -6.1235169e-11
+ lpdiblc2 = 3.7903799e-9
+ rshg = 15.6
+ rnoia = 0
+ rnoib = 0
+ wtvoff = 5.5500668e-10
+ ptvfbsdoff = 0
+ pketa = -3.1399835e-15
+ ngate = 8e+20
+ ngcon = 1
+ wpclm = -9.7111111e-9
+ capmod = 2
+ wku0we = 2e-11
+ gbmin = 1e-12
+ nigbacc = 10
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ mobmod = 0
+ tnom = 25
+ toxe = 2.3900000000000002e-9
+ toxm = 2.43e-9
+ lkvth0we = -2e-12
+ nigbinv = 10
+ acnqsmod = 0
+ wags = 1.7657181000000002e-8
+ rbodymod = 0
+ wcit = -3.0323584e-10
+ voff = -0.078900611
+ tvoff = -3.4914836e-5
+ acde = 0.4
+ fnoimod = 1
+ xjbvd = 1
+ xjbvs = 1
+ vsat = 84306.193
+ lk2we = -1.5e-12
+ eigbinv = 1.1
+ wint = 0
+ vth0 = 0.32093651999999995
+ wkt1 = 1.158409e-8
+ wkt2 = -3.7001265e-9
+ wmax = 2.674e-7
+ aigc = 0.011721192
+ wmin = 1.08e-7
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ ku0we = -0.0007
+ beta0 = 13
+ leta0 = 0
+ wpdiblc2 = 4.3752159e-9
+ wua1 = -6.5376855e-17
+ wub1 = 8.5457734e-26
+ wuc1 = 1.5793115e-17
+ bigc = 0.001442
+ wwlc = 0
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ cigbacc = 0.32875
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.5522823e-12
+ cgdo = 5.2490134000000004e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.5522823e-12
+ cgso = 5.2490134000000004e-11
+ tnoimod = 0
+ cigc = 0.000625
+ toxref = 3e-9
+ dmcgt = 0
+ tcjsw = 0.000357
+ wkvth0we = 2e-12
+ cigbinv = 0.006
+ trnqsmod = 0
+ bigsd = 0.00125
+ version = 4.5
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ tempmod = 0
+ ltvoff = 1.0403103e-9
+ wvoff = -2.1121636e-9
+ k2we = 5e-5
+ wvsat = 0.002322956
+ aigbacc = 0.02
+ dsub = 0.75
+ wvth0 = -4.2014741000000004e-9
+ dtox = 2.7e-10
+ rgatemod = 0
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ tnjtsswg = 1
+ waigc = 1.00872e-11
+ pvfbsdoff = 0
+ lku0we = 2.5e-11
+ epsrox = 3.9
+ eta0 = 0.2
+ etab = -0.2
+ lketa = 1.3109546e-8
+ aigbinv = 0.0163
+ xpart = 1
+ rdsmod = 0
+ igbmod = 1
+ egidl = 0.29734
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ pbswgd = 0.95
+ pbswgs = 0.95
+ igcmod = 1
+ poxedge = 1
+ binunit = 2
+ pvoff = 3.1183375e-15
+ cdscb = 0
+ cdscd = 0
+ pvsat = -1.8e-11
+ wk2we = 5e-12
+ pvth0 = -1.7129756e-15
+ drout = 0.56
+ permod = 1
+ paigc = 3.0482801e-18
+ ijthsfwd = 0.01
+ )

.model nch_ff_36 nmos (
+ level = 54
+ rshg = 15.6
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ cigbacc = 0.32875
+ tnoimod = 0
+ ku0we = -0.0007
+ a0 = 2.8517872
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ beta0 = 13
+ at = 72186.119
+ cf = 8.720500000000001e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.0021801551
+ k3 = -1.8419
+ em = 1000000.0
+ leta0 = 0
+ rgatemod = 0
+ ll = -1.18e-13
+ lw = 0
+ u0 = 0.010528434000000001
+ tpbswg = 0.0009
+ w0 = 0
+ ua = -2.2247872e-9
+ ub = 2.0937783e-18
+ uc = 7.1203963e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 2.33e-9
+ tnjtsswg = 1
+ ww = 0
+ xw = 8.600000000000001e-9
+ cigbinv = 0.006
+ tnom = 25
+ ppclm = 2.75592e-14
+ toxe = 2.3900000000000002e-9
+ toxm = 2.43e-9
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ ptvoff = 2.8225911e-16
+ version = 4.5
+ waigsd = 3.178874e-12
+ tempmod = 0
+ dmcgt = 0
+ tcjsw = 0.000357
+ diomod = 1
+ wags = 2.3108180000000002e-7
+ aigbacc = 0.02
+ wcit = 2.3683634e-10
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 2.6226e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.6226e-10
+ voff = -0.13810998
+ acde = 0.4
+ bigsd = 0.00125
+ vsat = 84306.193
+ wint = 0
+ vth0 = 0.38355441999999995
+ wtvfbsdoff = 0
+ wkt1 = -4.0570622999999995e-8
+ wkt2 = -4.3121065e-11
+ aigbinv = 0.0163
+ wmax = 2.674e-7
+ mjswgd = 0.85
+ mjswgs = 0.85
+ aigc = 0.011581706
+ wmin = 1.08e-7
+ wvoff = 7.1640927e-9
+ tcjswg = 0.001
+ wvsat = 0.002322956
+ ltvfbsdoff = 0
+ wvth0 = -9.9496131e-9
+ wua1 = 2.3276683e-17
+ wub1 = 1.5603072e-26
+ wuc1 = -5.1034561e-18
+ waigc = 2.6093343e-11
+ pvfbsdoff = 0
+ bigc = 0.001442
+ wwlc = 0
+ lketa = -3.8407777e-8
+ ijthsfwd = 0.01
+ cdsc = 0
+ xpart = 1
+ cgbo = 0
+ cgdl = 3.5522823e-12
+ cgdo = 5.2490134000000004e-11
+ xtid = 3
+ xtis = 3
+ poxedge = 1
+ cgsl = 3.5522823e-12
+ cgso = 5.2490134000000004e-11
+ cigc = 0.000625
+ egidl = 0.29734
+ fprout = 300
+ ptvfbsdoff = 0
+ binunit = 2
+ xrcrg1 = 12
+ xrcrg2 = 1
+ ijthsrev = 0.01
+ wtvoff = -1.1880818e-9
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ capmod = 2
+ k2we = 5e-5
+ wku0we = 2e-11
+ ppdiblc2 = 3.3310302e-16
+ dsub = 0.75
+ dtox = 2.7e-10
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ pvoff = -9.6321526e-16
+ mobmod = 0
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ cdscb = 0
+ cdscd = 0
+ pvsat = -1.8e-11
+ wk2we = 5e-12
+ pvth0 = 8.162056000000001e-16
+ drout = 0.56
+ eta0 = 0.2
+ etab = -0.2
+ paigc = -3.9944226e-18
+ voffl = 0
+ weta0 = 0
+ pkvth0we = -1.3e-19
+ ags = -2.6447884999999998
+ lpclm = -2.4174737e-7
+ cjd = 0.0012620099999999998
+ cit = 0.00083484714
+ cjs = 0.0012620099999999998
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 1.30529375e-8
+ k3b = 1.9326
+ njtsswg = 9
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ cgidl = 0.22
+ vfbsdoff = 0.02
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ la0 = -8.4086042e-7
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = 0.0055354098
+ kt1 = -0.088256509
+ lk2 = -6.7273888e-9
+ kt2 = -0.075738087
+ ckappad = 0.6
+ ckappas = 0.6
+ llc = -1.18e-13
+ lln = 0.7
+ lu0 = -5.2339671e-10
+ mjd = 0.26
+ pdiblc1 = 0
+ pdiblc2 = 0.031716534
+ lua = 3.6483177e-18
+ mjs = 0.26
+ lub = -6.2349821e-26
+ luc = -1.6579966e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ pdiblcb = -0.3
+ njd = 1.02
+ njs = 1.02
+ pa0 = 8.661463e-14
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ pbswd = 0.8
+ pbsws = 0.8
+ nsd = 1e+20
+ pbd = 0.52
+ pat = -3.1698679e-9
+ pbs = 0.52
+ pk2 = -2.2869691e-16
+ paramchk = 1
+ pu0 = 4.4409578e-18
+ prt = 0
+ pua = -4.9144669e-25
+ pub = 1.8790045e-33
+ puc = 1.8346553e-24
+ pud = 0
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 5.8363721e-10
+ ub1 = -5.3348382e-19
+ uc1 = 8.6067289e-11
+ tpb = 0.0014
+ wa0 = -2.3569588e-7
+ ute = -1
+ wat = 0.013137708
+ pdits = 0
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 2.3848778e-9
+ wlc = 0
+ wln = 1
+ cigsd = 0.069865
+ wu0 = -7.947186999999997e-12
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -2.0950609e-17
+ wub = 2.8553091e-26
+ wuc = -4.8106046e-18
+ wud = 0
+ wwc = 0
+ bigbacc = 0.002588
+ wwl = 0
+ wwn = 1
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ ijthdfwd = 0.01
+ kvth0we = 0.00018
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ toxref = 3e-9
+ lintnoi = -1.5e-8
+ keta = 0.053210932
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ tnoia = 0
+ lags = 1.4146322e-6
+ ijthdrev = 0.01
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ peta0 = 0
+ lcit = 3.3640592e-10
+ wketa = -7.2433388e-9
+ kt1l = 0
+ lpdiblc2 = -5.676798e-9
+ tpbsw = 0.0019
+ cjswd = 7.625999999999999e-11
+ cjsws = 7.625999999999999e-11
+ mjswd = 0.11
+ tvfbsdoff = 0.022
+ mjsws = 0.11
+ ltvoff = -1.663256e-9
+ agidl = 9.41e-8
+ lint = 9.7879675e-9
+ lkt1 = -7.280770300000001e-8
+ lkt2 = -5.7687528e-9
+ lmax = 4.5075e-7
+ lmin = 2.1744e-7
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ minv = -0.3
+ lku0we = 2.5e-11
+ lua1 = 4.6540649e-17
+ lub1 = -5.3739597e-26
+ luc1 = -7.7582888e-18
+ epsrox = 3.9
+ lkvth0we = -2e-12
+ ndep = 1e+18
+ nfactor = 1
+ lwlc = 0
+ moin = 5.1
+ scref = 1e-6
+ rdsmod = 0
+ pigcd = 2.621
+ nigc = 3.083
+ igbmod = 1
+ aigsd = 0.010772573
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ acnqsmod = 0
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ lvoff = -2.4242325e-9
+ pbswgd = 0.95
+ noff = 2.7195
+ pbswgs = 0.95
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ lvsat = -0.0003
+ rbodymod = 0
+ lvth0 = -8.897068699999999e-9
+ igcmod = 1
+ nigbacc = 10
+ delta = 0.007595625
+ pags = -1.0314937e-13
+ laigc = 1.3898222e-13
+ ntox = 2.029
+ pcit = -9.382386e-17
+ pclm = 2.434611
+ rnoia = 0
+ rnoib = 0
+ phin = 0.15
+ pketa = 2.46808e-15
+ ngate = 8e+20
+ nigbinv = 10
+ ngcon = 1
+ wpclm = -7.2345657e-8
+ pkt1 = 9.6867187e-15
+ pkt2 = 1.7671038e-16
+ wpdiblc2 = 6.3151306e-10
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ permod = 1
+ rbdb = 50
+ pua1 = -7.4684646e-24
+ prwb = 0
+ prwg = 0
+ pub1 = -7.978346e-34
+ puc1 = 1.3960704e-24
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ fnoimod = 1
+ rdsw = 100
+ eigbinv = 1.1
+ wkvth0we = 2e-12
+ voffcv = -0.16942
+ wpemod = 1
+ trnqsmod = 0
+ tvoff = 0.006109554
+ )

.model nch_ff_37 nmos (
+ level = 54
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ pdits = 0
+ cigsd = 0.069865
+ lkvth0we = -2e-12
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ eta0 = 0.2
+ etab = -0.2
+ ptvoff = -1.8615536e-17
+ waigsd = 3.178874e-12
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ acnqsmod = 0
+ diomod = 1
+ wtvfbsdoff = 0
+ tnoia = 0
+ pditsd = 0
+ pditsl = 0
+ rbodymod = 0
+ cjswgd = 2.6226e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.6226e-10
+ a0 = -2.4455841
+ a1 = 0
+ a2 = 1
+ peta0 = 0
+ b0 = 0
+ b1 = 0
+ ltvfbsdoff = 0
+ at = 121458.51
+ cf = 8.720500000000001e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = -0.007397302
+ k3 = -1.8419
+ em = 1000000.0
+ ll = -1.18e-13
+ wketa = 1.5290605e-8
+ lw = 0
+ u0 = 0.008924213
+ w0 = 0
+ ua = -2.2679307e-9
+ ub = 1.903479518e-18
+ uc = 2.5998306e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 2.33e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ tpbsw = 0.0019
+ nfactor = 1
+ tvfbsdoff = 0.022
+ cjswd = 7.625999999999999e-11
+ cjsws = 7.625999999999999e-11
+ mjswgd = 0.85
+ mjswd = 0.11
+ mjswgs = 0.85
+ mjsws = 0.11
+ agidl = 9.41e-8
+ tcjswg = 0.001
+ wpdiblc2 = 2.0871493e-9
+ ptvfbsdoff = 0
+ nigbacc = 10
+ scref = 1e-6
+ wvfbsdoff = 0
+ pigcd = 2.621
+ lvfbsdoff = 0
+ aigsd = 0.010772573
+ fprout = 300
+ lvoff = 4.451419999999998e-11
+ nigbinv = 10
+ keta = -0.11923047
+ xrcrg1 = 12
+ xrcrg2 = 1
+ wkvth0we = 2e-12
+ lvsat = -0.000689274295
+ lvth0 = -7.9619377e-9
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ trnqsmod = 0
+ delta = 0.007595625
+ lcit = -4.9333293e-11
+ wtvoff = 2.3786433e-10
+ laigc = -6.7426314e-12
+ kt1l = 0
+ rnoia = 0
+ rnoib = 0
+ fnoimod = 1
+ lint = 9.7879675e-9
+ pketa = -2.286582e-15
+ ngate = 8e+20
+ capmod = 2
+ eigbinv = 1.1
+ lkt1 = -5.412061899999999e-10
+ lkt2 = 1.6714521e-10
+ lmax = 2.1744e-7
+ ngcon = 1
+ lmin = 9.167e-8
+ wpclm = 1.5314007e-7
+ wku0we = 2e-11
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ mobmod = 0
+ rgatemod = 0
+ gbmin = 1e-12
+ tnjtsswg = 1
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ minv = -0.3
+ lua1 = -6.7367772e-18
+ lub1 = -3.8361216e-26
+ luc1 = -1.0970607e-17
+ ndep = 1e+18
+ lwlc = 0
+ moin = 5.1
+ nigc = 3.083
+ cigbacc = 0.32875
+ tnoimod = 0
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ cigbinv = 0.006
+ tvoff = -0.0028392003
+ ntox = 2.029
+ pcit = -5.942800000000005e-20
+ pclm = 1.0592301
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ phin = 0.15
+ version = 4.5
+ tempmod = 0
+ pkt1 = -2.3629532999999997e-16
+ pkt2 = -2.0087744e-16
+ ku0we = -0.0007
+ beta0 = 13
+ leta0 = 0
+ ppclm = -2.0018289e-14
+ aigbacc = 0.02
+ rbdb = 50
+ pua1 = 2.2068447e-24
+ prwb = 0
+ prwg = 0
+ pub1 = -2.7426774e-33
+ puc1 = 1.8773731e-24
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ ijthsfwd = 0.01
+ rdsw = 100
+ toxref = 3e-9
+ aigbinv = 0.0163
+ dmcgt = 0
+ tcjsw = 0.000357
+ ijthsrev = 0.01
+ rshg = 15.6
+ bigsd = 0.00125
+ ltvoff = 2.2493116e-10
+ wvoff = 1.8056166e-9
+ poxedge = 1
+ wvsat = 0.00180338308
+ ppdiblc2 = 2.596377e-17
+ wvth0 = -4.284810300000001e-9
+ binunit = 2
+ pvfbsdoff = 0
+ lku0we = 2.5e-11
+ waigc = 5.3999849e-12
+ tnom = 25
+ epsrox = 3.9
+ toxe = 2.3900000000000002e-9
+ toxm = 2.43e-9
+ rdsmod = 0
+ lketa = -2.0226409e-9
+ igbmod = 1
+ xpart = 1
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ egidl = 0.29734
+ pbswgd = 0.95
+ pbswgs = 0.95
+ pkvth0we = -1.3e-19
+ wags = -2.5777778e-7
+ igcmod = 1
+ wcit = -2.0754486e-10
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ voff = -0.149810363
+ acde = 0.4
+ vfbsdoff = 0.02
+ vsat = 86151.12359999999
+ wint = 0
+ vth0 = 0.379122633
+ wkt1 = 6.4578791e-9
+ wkt2 = 1.7463947e-9
+ wmax = 2.674e-7
+ aigc = 0.01161432
+ wmin = 1.08e-7
+ paramchk = 1
+ pvoff = 1.6741822e-16
+ wua1 = -2.2577864e-17
+ wub1 = 2.4820337e-26
+ wuc1 = -7.3845115e-18
+ cdscb = 0
+ cdscd = 0
+ bigc = 0.001442
+ permod = 1
+ pvsat = 9.163312000000007e-11
+ wwlc = 0
+ njtsswg = 9
+ wk2we = 5e-12
+ pvth0 = -3.7906062e-16
+ drout = 0.56
+ ags = 4.0596296
+ paigc = 3.7187593e-19
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ ijthdfwd = 0.01
+ cdsc = 0
+ cjd = 0.0012620099999999998
+ cit = 0.0026629951
+ cgbo = 0
+ cjs = 0.0012620099999999998
+ clc = 1e-7
+ cle = 0.6
+ voffl = 0
+ cgdl = 3.5522823e-12
+ bvd = 8.7
+ cgdo = 5.2490134000000004e-11
+ xtid = 3
+ bvs = 8.7
+ xtis = 3
+ dlc = 1.30529375e-8
+ ckappad = 0.6
+ ckappas = 0.6
+ k3b = 1.9326
+ cgsl = 3.5522823e-12
+ cgso = 5.2490134000000004e-11
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ cigc = 0.000625
+ pdiblc1 = 0
+ pdiblc2 = 0.0095469071
+ pdiblcb = -0.3
+ weta0 = 0
+ voffcv = -0.16942
+ wpemod = 1
+ lpclm = 4.8457997e-8
+ la0 = 2.768849e-7
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.0048610641000000005
+ kt1 = -0.43075175
+ lk2 = -4.7065454e-9
+ kt2 = -0.10387031
+ ijthdrev = 0.01
+ llc = -1.18e-13
+ lln = 0.7
+ lu0 = -1.8490616999999998e-10
+ mjd = 0.26
+ mjs = 0.26
+ lua = 1.2751594e-17
+ lub = -2.21968369e-26
+ cgidl = 0.22
+ luc = -7.0415723e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = -2.9632335e-14
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 4.745644e-10
+ pbs = 0.52
+ pk2 = 3.1759465e-16
+ lpdiblc2 = -9.9900678e-10
+ pu0 = 2.42802262e-18
+ bigbacc = 0.002588
+ prt = 0
+ pua = 3.9870432e-24
+ pub = -6.31495433e-33
+ puc = 2.2635812e-25
+ pud = 0
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 8.3613685e-10
+ ub1 = -6.0636714e-19
+ uc1 = 1.0129155e-10
+ tpb = 0.0014
+ wa0 = 3.1523761e-7
+ kvth0we = 0.00018
+ pbswd = 0.8
+ pbsws = 0.8
+ ute = -1
+ wat = -0.0041344832
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -2.0418175e-10
+ wlc = 0
+ wln = 1
+ wu0 = 1.5927899999999993e-12
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -4.2175679e-17
+ wub = 6.73870221e-26
+ wuc = 2.8116572e-18
+ wud = 0
+ k2we = 5e-5
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ lintnoi = -1.5e-8
+ tpbswg = 0.0009
+ dsub = 0.75
+ bigbinv = 0.004953
+ dtox = 2.7e-10
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ )

.model nch_ff_38 nmos (
+ level = 54
+ dmcgt = 0
+ poxedge = 1
+ pkvth0we = -1.3e-19
+ tcjsw = 0.000357
+ pditsd = 0
+ pditsl = 0
+ noff = 2.7195
+ cjswgd = 2.6226e-10
+ pku0we = -1.5e-18
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ cjswgs = 2.6226e-10
+ binunit = 2
+ vfbsdoff = 0.02
+ ntox = 2.029
+ pcit = 7.2565761e-18
+ pclm = 2.2357699
+ bigsd = 0.00125
+ ptvfbsdoff = 0
+ mjswgd = 0.85
+ mjswgs = 0.85
+ tcjswg = 0.001
+ phin = 0.15
+ wvoff = 4.874463324000002e-9
+ paramchk = 1
+ pkt1 = -1.1181124000000001e-15
+ pkt2 = 3.9546557e-16
+ wvsat = 0.0007260740999999998
+ wvth0 = -5.735803399999999e-9
+ pvfbsdoff = 0
+ waigc = -1.2918923e-11
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ rbdb = 50
+ pua1 = -4.7371604e-25
+ prwb = 0
+ pub1 = -1.1520112000000002e-33
+ prwg = 0
+ puc1 = -4.218097e-24
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ lketa = 2.9224258e-8
+ a0 = 0.7744856
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ ijthdfwd = 0.01
+ at = 96107.1884
+ cf = 8.720500000000001e-11
+ xpart = 1
+ ef = 1.0
+ k1 = 0.274
+ k2 = -0.045338197000000004
+ k3 = -1.8419
+ em = 1000000.0
+ rdsw = 100
+ ll = 0
+ lw = 0
+ u0 = 0.004811909499999999
+ w0 = 0
+ ua = -2.6695158e-9
+ ub = 2.0926996330000003e-18
+ uc = -9.6044814e-11
+ ud = 0
+ fprout = 300
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 2.33e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ xrcrg1 = 12
+ xrcrg2 = 1
+ egidl = 0.29734
+ ijthdrev = 0.01
+ wtvoff = 2.7545299e-10
+ lpdiblc2 = 4.9724259e-14
+ rshg = 15.6
+ njtsswg = 9
+ capmod = 2
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ wku0we = 2e-11
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = -0.0010813536
+ mobmod = 0
+ pdiblcb = -0.3
+ ags = 4.0596296
+ pvoff = -1.2105337000000015e-16
+ cjd = 0.0012620099999999998
+ cit = 0.0019976869999999997
+ cjs = 0.0012620099999999998
+ clc = 1e-7
+ cle = 0.6
+ cdscb = 0
+ cdscd = 0
+ bvd = 8.7
+ tnom = 25
+ bvs = 8.7
+ dlc = 3.26497e-9
+ pvsat = 1.9290050000000003e-10
+ k3b = 1.9326
+ lkvth0we = -2e-12
+ wk2we = 5e-12
+ toxe = 2.3900000000000002e-9
+ dwb = 0
+ dwc = 0
+ toxm = 2.43e-9
+ dwg = 0
+ dwj = 0
+ pvth0 = -2.426664999999999e-16
+ drout = 0.56
+ paigc = 2.0938533e-18
+ bigbacc = 0.002588
+ la0 = -2.5801646e-8
+ voffl = 0
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.00247804025
+ kt1 = -0.57243179
+ kt2 = -0.068117715
+ lk2 = -1.1401013e-9
+ llc = 0
+ lln = 1
+ lu0 = 2.0165036e-10
+ mjd = 0.26
+ acnqsmod = 0
+ mjs = 0.26
+ lua = 5.0500592e-17
+ lub = -3.9983527e-26
+ luc = 4.4304811e-18
+ lud = 0
+ laigsd = 1.06572e-17
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ kvth0we = 0.00018
+ weta0 = 4.2794074e-8
+ pa0 = 2.9413877e-15
+ wetab = -1.5859302e-8
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 3.5510969e-10
+ pbs = 0.52
+ pk2 = 2.316472e-16
+ lpclm = -6.2136744e-8
+ pu0 = -3.5928665e-17
+ wags = -2.5777778e-7
+ prt = 0
+ pua = -3.0159915e-24
+ pub = 1.3943639e-33
+ puc = 2.394639e-25
+ pud = 0
+ lintnoi = -1.5e-8
+ rbodymod = 0
+ wcit = -2.85374837e-10
+ bigbinv = 0.004953
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 7.2026227e-10
+ vtsswgd = 4.2
+ ub1 = -8.527562e-19
+ vtsswgs = 4.2
+ uc1 = -2.7209866e-10
+ cgidl = 0.22
+ tpb = 0.0014
+ wa0 = -3.1291358e-8
+ voff = -0.11849200800000002
+ ute = -1
+ wat = -0.0028636889599999993
+ acde = 0.4
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 7.1015279e-10
+ wlc = 0
+ wln = 1
+ wu0 = 4.0964264e-10
+ xgl = -1.09e-8
+ xgw = 0
+ wua = 3.2324691e-17
+ wub = -1.4627000299999995e-26
+ wuc = 2.6722336e-18
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ vsat = 67284.95300000001
+ wint = 0
+ vth0 = 0.25413830800000003
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ wkt1 = 1.5838826000000005e-8
+ wkt2 = -4.5976799e-9
+ wmax = 2.674e-7
+ aigc = 0.011905208
+ wmin = 1.08e-7
+ pbswd = 0.8
+ pbsws = 0.8
+ wpdiblc2 = 2.3634934e-9
+ wua1 = 5.9387403e-18
+ wub1 = 7.898373999999995e-27
+ wuc1 = 5.7460914e-17
+ pdits = 0
+ bigc = 0.001442
+ cigsd = 0.069865
+ wwlc = 0
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ cdsc = 0
+ nfactor = 1
+ toxref = 3e-9
+ cgbo = 0
+ cgdl = 3.5522823e-12
+ cgdo = 5.2490134000000004e-11
+ xtid = 3
+ xtis = 3
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ cgsl = 3.5522823e-12
+ cgso = 5.2490134000000004e-11
+ cigc = 0.000625
+ wkvth0we = 2e-12
+ tnoia = 0
+ peta0 = -4.0226429e-15
+ trnqsmod = 0
+ petab = 1.4907744e-15
+ wketa = -4.815885e-9
+ tpbsw = 0.0019
+ ltvoff = 1.3417313e-10
+ nigbacc = 10
+ tvfbsdoff = 0.022
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ cjswd = 7.625999999999999e-11
+ cjsws = 7.625999999999999e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ k2we = 5e-5
+ nigbinv = 10
+ dsub = 0.75
+ rgatemod = 0
+ lku0we = 2.5e-11
+ dtox = 2.7e-10
+ tnjtsswg = 1
+ epsrox = 3.9
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ rdsmod = 0
+ eta0 = -0.13238438
+ etab = 0.18670848
+ igbmod = 1
+ scref = 1e-6
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ pigcd = 2.621
+ aigsd = 0.010772573
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ fnoimod = 1
+ pbswgd = 0.95
+ pbswgs = 0.95
+ eigbinv = 1.1
+ lvoff = -2.899411200000001e-9
+ igcmod = 1
+ lvsat = 0.0010841461499999999
+ lvth0 = 3.786589499999999e-9
+ delta = 0.007595625
+ laigc = -3.4086068e-11
+ rnoia = 0
+ rnoib = 0
+ pketa = -3.9657201e-16
+ ngate = 8e+20
+ paigsd = -2.9413875e-24
+ ngcon = 1
+ cigbacc = 0.32875
+ wpclm = -8.3073835e-8
+ gbmin = 1e-12
+ tnoimod = 0
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ permod = 1
+ cigbinv = 0.006
+ ijthsfwd = 0.01
+ voffcv = -0.16942
+ wpemod = 1
+ version = 4.5
+ keta = -0.45164428
+ tempmod = 0
+ ijthsrev = 0.01
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 1.3205699999999998e-11
+ tvoff = -0.0018736893
+ aigbacc = 0.02
+ kt1l = 0
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ lint = 0
+ lkt1 = 1.2776722e-8
+ lkt2 = -3.1935983e-9
+ lmax = 9.167e-8
+ lmin = 5.567e-8
+ tpbswg = 0.0009
+ ku0we = -0.0007
+ aigbinv = 0.0163
+ beta0 = 13
+ lpe0 = 9.2e-8
+ ppdiblc2 = -1.2574432e-20
+ lpeb = 2.5e-7
+ leta0 = 3.1244132e-8
+ letab = -3.6350598e-8
+ wtvfbsdoff = 0
+ minv = -0.3
+ ppclm = 2.1858187e-15
+ lua1 = 4.1554342e-18
+ lub1 = -1.5200603e-26
+ luc1 = 2.4128073e-17
+ ndep = 1e+18
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ ptvoff = -2.2148869e-17
+ lwlc = 0
+ moin = 5.1
+ ltvfbsdoff = 0
+ waigsd = 3.1789053e-12
+ nigc = 3.083
+ diomod = 1
+ )

.model nch_ff_39 nmos (
+ level = 54
+ wkt1 = 9.916755e-9
+ wkt2 = 1.1625249e-8
+ wmax = 2.674e-7
+ aigc = 0.011615807
+ wmin = 1.08e-7
+ fnoimod = 1
+ eigbinv = 1.1
+ wua1 = -1.0774777e-16
+ wub1 = 9.880248999999997e-26
+ wuc1 = 1.606153e-17
+ bigc = 0.001442
+ wwlc = 0
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ scref = 1e-6
+ ijthsfwd = 0.01
+ cdsc = 0
+ fprout = 300
+ pigcd = 2.621
+ cgbo = 0
+ aigsd = 0.010772573
+ cgdl = 3.5522823e-12
+ cgdo = 5.2490134000000004e-11
+ xtid = 3
+ xtis = 3
+ xrcrg1 = 12
+ xrcrg2 = 1
+ cgsl = 3.5522823e-12
+ cgso = 5.2490134000000004e-11
+ cigc = 0.000625
+ lvoff = -6.508439899999999e-9
+ cigbacc = 0.32875
+ lvsat = -0.0025682031000000003
+ wtvoff = 7.91509e-11
+ lvth0 = 8.278550700000002e-9
+ ijthsrev = 0.01
+ tnoimod = 0
+ delta = 0.007595625
+ laigc = -1.730084e-11
+ rnoia = 0
+ rnoib = 0
+ cigbinv = 0.006
+ dmcg = 3.1e-8
+ capmod = 2
+ dmci = 3.1e-8
+ dmdg = 0
+ wku0we = 2e-11
+ pketa = 1.224516e-15
+ ngate = 8e+20
+ a0 = 19.191807
+ a1 = 0
+ a2 = 1
+ ngcon = 1
+ b0 = 0
+ b1 = 0
+ mobmod = 0
+ wpclm = -5.2664346e-8
+ at = 147437.86199999996
+ cf = 8.720500000000001e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = -0.059713829
+ k3 = -1.8419
+ em = 1000000.0
+ k2we = 5e-5
+ ll = 0
+ lw = 0
+ u0 = 0.0023880985
+ w0 = 0
+ ua = -2.3710013e-9
+ ub = 1.4550579529999998e-18
+ uc = -1.4785261e-10
+ ud = 0
+ version = 4.5
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 2.33e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ dsub = 0.75
+ dtox = 2.7e-10
+ gbmin = 1e-12
+ tempmod = 0
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ eta0 = 1.1504337
+ aigbacc = 0.02
+ etab = -1.3364008
+ pkvth0we = -1.3e-19
+ aigbinv = 0.0163
+ tvoff = -0.0045522389
+ vfbsdoff = 0.02
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ paramchk = 1
+ ku0we = -0.0007
+ beta0 = 13
+ leta0 = -4.3159315e-8
+ poxedge = 1
+ letab = 5.198974e-8
+ ppclm = 4.2206835e-16
+ binunit = 2
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ ijthdfwd = 0.01
+ toxref = 3e-9
+ dmcgt = 0
+ keta = 0.16119603
+ tcjsw = 0.000357
+ ijthdrev = 0.01
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 2.6466223e-10
+ ltvoff = 2.8952901e-10
+ kt1l = 0
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ bigsd = 0.00125
+ lint = 0
+ wvoff = -2.2288246e-9
+ lkt1 = 1.8120665000000003e-8
+ lkt2 = 8.1983323e-9
+ lmax = 5.567e-8
+ lmin = 4.667e-8
+ wvsat = 0.0017322021999999996
+ lku0we = 2.5e-11
+ pvfbsdoff = 0
+ lpe0 = 9.2e-8
+ wvth0 = -1.00788921e-8
+ lpeb = 2.5e-7
+ epsrox = 3.9
+ waigc = 4.0939876e-11
+ minv = -0.3
+ lua1 = -3.9796071e-17
+ lub1 = 4.008477099999999e-26
+ luc1 = 1.4911728e-19
+ rdsmod = 0
+ lkvth0we = -2e-12
+ ndep = 1e+18
+ igbmod = 1
+ lwlc = 0
+ lketa = -6.3204807e-9
+ moin = 5.1
+ njtsswg = 9
+ xpart = 1
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ nigc = 3.083
+ pbswgd = 0.95
+ pbswgs = 0.95
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ acnqsmod = 0
+ egidl = 0.29734
+ igcmod = 1
+ ckappad = 0.6
+ ckappas = 0.6
+ noff = 2.7195
+ pdiblc1 = 0
+ pdiblc2 = -0.0010804963
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ pdiblcb = -0.3
+ rbodymod = 0
+ ntox = 2.029
+ pcit = 6.109152999999998e-18
+ pclm = 1.0542662
+ ags = 4.0596296
+ bigbacc = 0.002588
+ phin = 0.15
+ cjd = 0.0012620099999999998
+ cit = -0.0023377727
+ cjs = 0.0012620099999999998
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 3.26497e-9
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ pkt1 = -7.746442400000001e-16
+ pkt2 = -5.454643e-16
+ dwg = 0
+ dwj = 0
+ kvth0we = 0.00018
+ wpdiblc2 = 2.3632766e-9
+ permod = 1
+ pvoff = 2.9093734999999984e-16
+ lintnoi = -1.5e-8
+ la0 = -1.0940063e-6
+ cdscb = 0
+ cdscd = 0
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.005455230580000001
+ bigbinv = 0.004953
+ kt1 = -0.66456841
+ kt2 = -0.26453031
+ lk2 = -3.0631458e-10
+ vtsswgd = 4.2
+ pvsat = 1.3454518000000005e-10
+ vtsswgs = 4.2
+ llc = 0
+ lln = 1
+ lu0 = 3.4223107999999997e-10
+ wk2we = 5e-12
+ pvth0 = 9.236253999999894e-18
+ mjd = 0.26
+ mjs = 0.26
+ lua = 3.3186753e-17
+ lub = -3.0003129999999985e-27
+ luc = 7.435334e-18
+ lud = 0
+ rbdb = 50
+ pua1 = 6.1201017e-24
+ prwb = 0
+ lwc = 0
+ pub1 = -6.424441900000002e-33
+ prwg = 0
+ drout = 0.56
+ lwl = 0
+ puc1 = -1.8169327e-24
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 1.2471671e-13
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ nsd = 1e+20
+ pvag = 1.2
+ pbd = 0.52
+ pat = -5.796346000000003e-11
+ pbs = 0.52
+ pk2 = 1.8168527e-16
+ paigc = -1.0299571e-18
+ pu0 = -1.1596503999999992e-18
+ prt = 0
+ pua = 6.5377716e-24
+ pub = -1.101976303e-32
+ rdsw = 100
+ puc = -3.076481e-25
+ pud = 0
+ voffl = 0
+ rsh = 17.5
+ tcj = 0.00076
+ voffcv = -0.16942
+ wpemod = 1
+ ua1 = 1.4780468e-9
+ ub1 = -1.8059528999999997e-18
+ uc1 = 1.4133161e-10
+ tpb = 0.0014
+ wa0 = -2.130866e-6
+ weta0 = -1.5669611e-7
+ ute = -1
+ wetab = 4.0317659e-8
+ wat = 0.004258294299999999
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 1.5715655e-9
+ wlc = 0
+ wln = 1
+ wu0 = -1.89823297e-10
+ lpclm = 6.3904735e-9
+ xgl = -1.09e-8
+ wkvth0we = 2e-12
+ xgw = 0
+ wua = -1.3239536e-16
+ wub = 1.9940967600000001e-25
+ wuc = 1.2105201e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ cgidl = 0.22
+ trnqsmod = 0
+ rshg = 15.6
+ wtvfbsdoff = 0
+ nfactor = 1
+ pbswd = 0.8
+ pbsws = 0.8
+ tpbswg = 0.0009
+ ltvfbsdoff = 0
+ rgatemod = 0
+ tnjtsswg = 1
+ pdits = 0
+ tnom = 25
+ cigsd = 0.069865
+ toxe = 2.3900000000000002e-9
+ ptvoff = -1.0763348e-17
+ toxm = 2.43e-9
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ waigsd = 3.1788545e-12
+ nigbacc = 10
+ pk2we = -1e-19
+ diomod = 1
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ ptvfbsdoff = 0
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 2.6226e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.6226e-10
+ wags = -2.5777778e-7
+ tnoia = 0
+ nigbinv = 10
+ wcit = -2.6559286000000003e-10
+ peta0 = 7.5477876e-15
+ petab = -1.7674893e-15
+ voff = -0.056267378999999965
+ wketa = -3.2765679e-8
+ acde = 0.4
+ tvfbsdoff = 0.022
+ tpbsw = 0.0019
+ mjswgd = 0.85
+ mjswgs = 0.85
+ vsat = 130256.523
+ wint = 0
+ cjswd = 7.625999999999999e-11
+ cjsws = 7.625999999999999e-11
+ vth0 = 0.17669063899999998
+ tcjswg = 0.001
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ )

.model nch_ff_40 nmos (
+ level = 54
+ wkt1 = 7.369332999999995e-9
+ wkt2 = -1.1473225e-8
+ wmax = 2.674e-7
+ aigc = 0.011144932
+ wmin = 1.08e-7
+ fnoimod = 1
+ eigbinv = 1.1
+ wua1 = 1.9140234e-16
+ wub1 = -2.262572e-25
+ wuc1 = -2.3798265000000004e-17
+ bigc = 0.001442
+ wwlc = 0
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ scref = 1e-6
+ ijthsfwd = 0.01
+ cdsc = 0
+ fprout = 300
+ pigcd = 2.621
+ cgbo = 0
+ aigsd = 0.010772574
+ cgdl = 3.5522823e-12
+ cgdo = 5.2490134000000004e-11
+ xtid = 3
+ xtis = 3
+ xrcrg1 = 12
+ xrcrg2 = 1
+ cgsl = 3.5522823e-12
+ cgso = 5.2490134000000004e-11
+ cigc = 0.000625
+ lvoff = -7.1267393e-9
+ cigbacc = 0.32875
+ lvsat = 0.00543648752
+ wtvoff = -7.2128996e-10
+ lvth0 = -2.7266051999999993e-9
+ ijthsrev = 0.01
+ tnoimod = 0
+ delta = 0.007595625
+ laigc = 5.7720314e-12
+ rnoia = 0
+ rnoib = 0
+ cigbinv = 0.006
+ dmcg = 3.1e-8
+ capmod = 2
+ dmci = 3.1e-8
+ dmdg = 0
+ wku0we = 2e-11
+ pketa = -8.4677334e-15
+ ngate = 8e+20
+ a0 = -5.925916599999999
+ a1 = 0
+ a2 = 1
+ ngcon = 1
+ b0 = 0
+ b1 = 0
+ mobmod = 0
+ wpclm = -7.2101286e-7
+ at = 15266.341999999997
+ cf = 8.720500000000001e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.013523130999999994
+ k3 = -1.8419
+ em = 1000000.0
+ k2we = 5e-5
+ ll = 0
+ lw = 0
+ u0 = 0.013645519
+ w0 = 0
+ ua = -5.589164400000002e-10
+ ub = 8.937269600000036e-20
+ uc = 2.381934e-10
+ ud = 0
+ version = 4.5
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 2.33e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ dsub = 0.75
+ dtox = 2.7e-10
+ gbmin = 1e-12
+ tempmod = 0
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ eta0 = -0.250734997
+ aigbacc = 0.02
+ etab = -0.74723747
+ laigsd = -1.5325105e-17
+ pkvth0we = -1.3e-19
+ aigbinv = 0.0163
+ tvoff = 0.0062987975
+ vfbsdoff = 0.02
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ paramchk = 1
+ ku0we = -0.0007
+ beta0 = 13
+ leta0 = 2.5497954e-8
+ poxedge = 1
+ letab = 2.3120738e-8
+ ppclm = 3.3171145e-14
+ binunit = 2
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ ijthdfwd = 0.01
+ toxref = 3e-9
+ dmcgt = 0
+ keta = -0.51478944
+ tcjsw = 0.000357
+ ijthdrev = 0.01
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 4.819485e-10
+ ltvoff = -2.4217179e-10
+ kt1l = 0
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ bigsd = 0.00125
+ lint = 0
+ wvoff = 1.3282831000000013e-9
+ lkt1 = -4.5298867e-9
+ lkt2 = -1.1864945e-9
+ lmax = 4.667e-8
+ lmin = 3.6e-8
+ wvsat = 0.0227104314
+ lku0we = 2.5e-11
+ pvfbsdoff = 0
+ lpe0 = 9.2e-8
+ wvth0 = -1.7093637e-8
+ lpeb = 2.5e-7
+ epsrox = 3.9
+ waigc = 5.1623453e-11
+ minv = -0.3
+ lua1 = 6.0050187e-18
+ lub1 = 7.877147000000001e-28
+ luc1 = 6.4275095e-18
+ rdsmod = 0
+ lkvth0we = -2e-12
+ ndep = 1e+18
+ igbmod = 1
+ lwlc = 0
+ lketa = 2.6802806000000003e-8
+ moin = 5.1
+ njtsswg = 9
+ xpart = 1
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ nigc = 3.083
+ pbswgd = 0.95
+ pbswgs = 0.95
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ acnqsmod = 0
+ egidl = 0.29734
+ igcmod = 1
+ ckappad = 0.6
+ ckappas = 0.6
+ noff = 2.7195
+ pdiblc1 = 0
+ pdiblc2 = -0.0010804963
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ pdiblcb = -0.3
+ rbodymod = 0
+ ntox = 2.029
+ pcit = 3.904200000000001e-19
+ pclm = 4.6708343
+ ags = 4.0596296
+ bigbacc = 0.002588
+ phin = 0.15
+ paigsd = 4.2297301e-24
+ cjd = 0.0012620099999999998
+ cit = -0.006772191700000001
+ cjs = 0.0012620099999999998
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 3.26497e-9
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ pkt1 = -6.4979764e-16
+ pkt2 = 5.863609e-16
+ dwg = 0
+ dwj = 0
+ kvth0we = 0.00018
+ wpdiblc2 = 2.3632766e-9
+ permod = 1
+ pvoff = 1.1663916e-16
+ lintnoi = -1.5e-8
+ la0 = 1.3676219000000002e-7
+ cdscb = 0
+ cdscd = 0
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = 0.0010211866800000002
+ bigbinv = 0.004953
+ kt1 = -0.20231328
+ kt2 = -0.073003235
+ lk2 = -3.894925700000001e-9
+ vtsswgd = 4.2
+ pvsat = -8.933872599999999e-10
+ vtsswgs = 4.2
+ llc = 0
+ lln = 1
+ lu0 = -2.0938226e-10
+ wk2we = 5e-12
+ pvth0 = 3.5295838999999996e-16
+ mjd = 0.26
+ mjs = 0.26
+ lua = -5.56054081e-17
+ lub = 6.391826569999999e-26
+ luc = -1.14809219e-17
+ lud = 0
+ rbdb = 50
+ pua1 = -8.5382538e-24
+ prwb = 0
+ lwc = 0
+ pub1 = 9.503469000000001e-33
+ prwg = 0
+ drout = 0.56
+ lwl = 0
+ puc1 = 1.361972e-25
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = -7.5523402e-14
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ nsd = 1e+20
+ pvag = 1.2
+ pbd = 0.52
+ pat = -1.1869552000000004e-10
+ pbs = 0.52
+ pk2 = 5.0756697e-16
+ paigc = -1.5534524e-18
+ pu0 = 6.5681068e-18
+ prt = 0
+ pua = -2.8276596999999977e-25
+ pub = -6.331388000000253e-35
+ rdsw = 100
+ puc = 4.398917e-25
+ pud = 0
+ voffl = 0
+ rsh = 17.5
+ tcj = 0.00076
+ voffcv = -0.16942
+ wpemod = 1
+ ua1 = 5.4333072e-10
+ ub1 = -1.00397154e-18
+ uc1 = 1.3201149999999995e-11
+ tpb = 0.0014
+ wa0 = 1.9556670799999998e-6
+ weta0 = 8.4602297e-8
+ ute = -1
+ wetab = 3.9258957e-9
+ wat = 0.005497692499999999
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -5.0790816e-9
+ wlc = 0
+ wln = 1
+ wu0 = -3.4753256999999996e-10
+ lpclm = -1.70821362e-7
+ xgl = -1.09e-8
+ wkvth0we = 2e-12
+ xgw = 0
+ wua = 6.799270000000015e-18
+ wub = -2.4191335000000008e-26
+ wuc = -3.150715e-18
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ cgidl = 0.22
+ trnqsmod = 0
+ rshg = 15.6
+ wtvfbsdoff = 0
+ nfactor = 1
+ pbswd = 0.8
+ pbsws = 0.8
+ tpbswg = 0.0009
+ ltvfbsdoff = 0
+ rgatemod = 0
+ tnjtsswg = 1
+ pdits = 0
+ tnom = 25
+ cigsd = 0.069865
+ toxe = 2.3900000000000002e-9
+ ptvoff = 2.8458255e-17
+ toxm = 2.43e-9
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ waigsd = 3.1787682e-12
+ nigbacc = 10
+ pk2we = -1e-19
+ diomod = 1
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ ptvfbsdoff = 0
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 2.6226e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.6226e-10
+ wags = -2.5777778e-7
+ tnoia = 0
+ nigbinv = 10
+ wcit = -1.4888078000000002e-10
+ peta0 = -4.2758338e-15
+ petab = 1.5707054e-17
+ voff = -0.043649036000000016
+ wketa = 1.65035329e-7
+ acde = 0.4
+ tvfbsdoff = 0.022
+ tpbsw = 0.0019
+ mjswgd = 0.85
+ mjswgs = 0.85
+ vsat = -33104.51799999998
+ wint = 0
+ cjswd = 7.625999999999999e-11
+ cjsws = 7.625999999999999e-11
+ vth0 = 0.401286047
+ tcjswg = 0.001
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ )

.model nch_fs_1 nmos (
+ level = 54
+ fprout = 300
+ xrcrg1 = 12
+ xrcrg2 = 1
+ ags = 0.7875000000000001
+ wtvoff = 0
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ tvoff = 0.0019109629
+ keta = -0.06
+ cjd = 0.001281008
+ cit = 0.0001
+ cjs = 0.001281008
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 9.8024918e-9
+ xjbvd = 1
+ k3b = 1.9326
+ xjbvs = 1
+ lk2we = -1.5e-12
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ tvfbsdoff = 0.022
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = -8e-12
+ capmod = 2
+ la0 = 0
+ kt1l = 0
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.00016
+ kt1 = -0.200226
+ kt2 = -0.05325
+ wku0we = 2e-11
+ wkvth0we = 2e-12
+ llc = 0
+ ku0we = -0.0007
+ lln = 1
+ lu0 = 9.600000000000001e-12
+ mjd = 0.26
+ mjs = 0.26
+ beta0 = 13
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ leta0 = 1.6000000000000003e-9
+ njs = 1.02
+ pa0 = 0
+ mobmod = 0
+ nsd = 1e+20
+ pbd = 0.52
+ pat = -3.04e-11
+ pbs = 0.52
+ lint = 6.5375218e-9
+ trnqsmod = 0
+ pu0 = 1.8400000000000002e-18
+ prt = 0
+ pud = 0
+ lkt1 = -4.8e-10
+ lmax = 2.001e-5
+ lmin = 8.9991e-6
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 1.2299687e-9
+ ub1 = -7.2455506e-19
+ uc1 = 3.028e-11
+ dlcig = 2.5e-9
+ tpb = 0.0014
+ lpe0 = 9.2e-8
+ njtsswg = 9
+ bgidl = 2320000000.0
+ lpeb = 2.5e-7
+ wa0 = 0
+ ute = -1.007
+ wat = 0
+ web = 6843.8
+ wec = -25529.0
+ wlc = 0
+ wln = 1
+ wu0 = -3.6000000000000005e-11
+ xgl = -1.09e-8
+ xgw = 0
+ wud = 0
+ wwc = 0
+ minv = -0.3
+ wwl = 0
+ wwn = 1
+ xtsswgd = 0.18
+ wvfbsdoff = 0
+ xtsswgs = 0.18
+ lvfbsdoff = 0
+ lub1 = -2.4000000000000004e-27
+ ndep = 1e+18
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.018555248
+ lwlc = 0
+ rgatemod = 0
+ dmcgt = 0
+ pdiblcb = -0.3
+ moin = 5.1
+ tcjsw = 0.000357
+ tnjtsswg = 1
+ nigc = 3.083
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ bigsd = 0.00125
+ bigbacc = 0.002588
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ wvoff = 0
+ ntox = 1.0
+ pcit = -1.2000000000000001e-17
+ kvth0we = 0.00018
+ pclm = 1.4
+ wvsat = 0
+ wvth0 = -3.2000000000000005e-9
+ lintnoi = -1.5e-8
+ bigbinv = 0.004953
+ phin = 0.15
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ pkt1 = 5.600000000000001e-17
+ a0 = 3.25
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 72000
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.023001254
+ k3 = -1.8419
+ em = 1000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.01539
+ w0 = 0
+ ua = -1.8237726e-9
+ ub = 2.103696e-18
+ xpart = 1
+ uc = 7.33e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ toxref = 3e-9
+ rbdb = 50
+ prwb = 0
+ prwg = 0
+ pub1 = -3.2e-34
+ egidl = 0.29734
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ rdsw = 100
+ ijthsfwd = 0.01
+ ltvoff = 0
+ nfactor = 1
+ rshg = 15.6
+ ijthsrev = 0.01
+ pvoff = 0
+ lku0we = 2.5e-11
+ cdscb = 0
+ cdscd = 0
+ epsrox = 3.9
+ pvsat = -2.24e-11
+ wk2we = 5e-12
+ pvth0 = -1.2e-16
+ drout = 0.56
+ nigbacc = 10
+ rdsmod = 0
+ igbmod = 1
+ voffl = 0
+ tnom = 25
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ weta0 = 0
+ pbswgd = 0.95
+ pbswgs = 0.95
+ nigbinv = 10
+ igcmod = 1
+ cgidl = 0.22
+ wags = -8e-9
+ wcit = 4.0000000000000004e-11
+ voff = -0.1128204
+ fnoimod = 1
+ pbswd = 0.8
+ pbsws = 0.8
+ acde = 0.4
+ pkvth0we = -1.3e-19
+ eigbinv = 1.1
+ vsat = 102860
+ wint = 0
+ vth0 = 0.32191089
+ wkt1 = -2.5600000000000003e-9
+ pvfbsdoff = 0
+ wmax = 0.00090001
+ aigc = 0.011769394
+ wmin = 8.9974e-6
+ pdits = 0
+ vfbsdoff = 0.02
+ permod = 1
+ cigsd = 0.069865
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ bigc = 0.001442
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ paramchk = 1
+ wwlc = 0
+ cigbacc = 0.32875
+ voffcv = -0.16942
+ wpemod = 1
+ cdsc = 0
+ tnoia = 0
+ tnoimod = 0
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ peta0 = 0.0
+ cigbinv = 0.006
+ tpbsw = 0.0019
+ ijthdfwd = 0.01
+ cjswd = 7.7408e-11
+ cjsws = 7.7408e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ version = 4.5
+ tempmod = 0
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ tpbswg = 0.0009
+ ijthdrev = 0.01
+ aigbacc = 0.02
+ k2we = 5e-5
+ dsub = 0.75
+ dtox = 2.7e-10
+ scref = 1e-6
+ ptvoff = 0
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ pigcd = 2.621
+ aigsd = 0.01077322
+ lvoff = -1.6e-11
+ eta0 = 0.3
+ aigbinv = 0.0163
+ diomod = 1
+ etab = -0.25
+ wtvfbsdoff = 0
+ lvsat = -0.0002
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 2.66208e-10
+ pku0we = -1.5e-18
+ lvth0 = -4.8e-10
+ cjswgs = 2.66208e-10
+ lkvth0we = -2e-12
+ delta = 0.007595625
+ ltvfbsdoff = 0
+ rnoia = 0
+ rnoib = 0
+ mjswgd = 0.85
+ mjswgs = 0.85
+ acnqsmod = 0
+ ngate = 8e+20
+ tcjswg = 0.001
+ ngcon = 1
+ poxedge = 1
+ rbodymod = 0
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ binunit = 2
+ ptvfbsdoff = 0
+ )

.model nch_fs_2 nmos (
+ level = 54
+ wtvoff = 0
+ cgidl = 0.22
+ ijthdfwd = 0.01
+ capmod = 2
+ pbswd = 0.8
+ pbsws = 0.8
+ wku0we = 2e-11
+ rshg = 15.6
+ cigbacc = 0.32875
+ mobmod = 0
+ pvfbsdoff = 0
+ ijthdrev = 0.01
+ tnoimod = 0
+ pdits = 0
+ lpdiblc2 = -5.8501673e-10
+ cigsd = 0.069865
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ cigbinv = 0.006
+ tnom = 25
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ version = 4.5
+ tnoia = 0
+ tempmod = 0
+ lkvth0we = -2e-12
+ peta0 = 0.0
+ tpbsw = 0.0019
+ aigbacc = 0.02
+ wags = -8e-9
+ cjswd = 7.7408e-11
+ cjsws = 7.7408e-11
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ wcit = 4.0000000000000004e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ acnqsmod = 0
+ voff = -0.11120139
+ acde = 0.4
+ vsat = 102860
+ wint = 0
+ rbodymod = 0
+ aigbinv = 0.0163
+ vth0 = 0.31616703
+ wkt1 = -2.5600000000000003e-9
+ wmax = 0.00090001
+ aigc = 0.01178613
+ wmin = 8.9974e-6
+ scref = 1e-6
+ pigcd = 2.621
+ toxref = 3e-9
+ aigsd = 0.01077322
+ bigc = 0.001442
+ wwlc = 0
+ lvoff = -1.4570874e-8
+ poxedge = 1
+ cdsc = 0
+ lvsat = -0.0002
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ lvth0 = 5.1157332e-8
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ delta = 0.007595625
+ binunit = 2
+ laigc = -1.5044982e-10
+ rnoia = 0
+ rnoib = 0
+ ltvoff = -1.4627394e-10
+ a0 = 3.4752469
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ ngate = 8e+20
+ at = 61592.494
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.024488843
+ k3 = -1.8419
+ em = 1000000.0
+ ngcon = 1
+ ll = 0
+ lw = 0
+ u0 = 0.015611951
+ w0 = 0
+ ua = -1.7995884e-9
+ ub = 2.1046515e-18
+ uc = 7.3387901e-11
+ ud = 0
+ wkvth0we = 2e-12
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ lku0we = 2.5e-11
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ trnqsmod = 0
+ epsrox = 3.9
+ k2we = 5e-5
+ rdsmod = 0
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ dsub = 0.75
+ dtox = 2.7e-10
+ igbmod = 1
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ ags = 0.79104901
+ pbswgd = 0.95
+ pbswgs = 0.95
+ eta0 = 0.3
+ cjd = 0.001281008
+ rgatemod = 0
+ etab = -0.25
+ cit = -2.3830864e-5
+ cjs = 0.001281008
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 9.8024918e-9
+ tnjtsswg = 1
+ k3b = 1.9326
+ igcmod = 1
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ tvoff = 0.0019272336
+ la0 = -2.0249698e-6
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = 0.09340348100000001
+ kt1 = -0.19577666
+ lk2 = -1.337342e-8
+ kt2 = -0.051823539
+ xjbvd = 1
+ llc = 0
+ xjbvs = 1
+ lln = 1
+ tvfbsdoff = 0.022
+ lk2we = -1.5e-12
+ lu0 = -1.9857361e-9
+ mjd = 0.26
+ lua = -2.1741579e-16
+ mjs = 0.26
+ lub = -8.5898229e-27
+ luc = -7.902321e-19
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njtsswg = 9
+ njd = 1.02
+ njs = 1.02
+ pa0 = 0
+ nsd = 1e+20
+ pbd = 0.52
+ pat = -3.04e-11
+ pbs = 0.52
+ pu0 = 1.8400000000000002e-18
+ xtsswgd = 0.18
+ prt = 0
+ pud = 0
+ xtsswgs = 0.18
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 1.2713861e-9
+ ub1 = -7.4616446e-19
+ ku0we = -0.0007
+ uc1 = 2.5703642e-11
+ ckappad = 0.6
+ ckappas = 0.6
+ beta0 = 13
+ tpb = 0.0014
+ wa0 = 0
+ leta0 = 1.6000000000000003e-9
+ pdiblc1 = 0
+ pdiblc2 = 0.018620322
+ pdiblcb = -0.3
+ ute = -1.0077691
+ wat = 0
+ web = 6843.8
+ wec = -25529.0
+ wlc = 0
+ wln = 1
+ wu0 = -3.6000000000000005e-11
+ xgl = -1.09e-8
+ xgw = 0
+ permod = 1
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ bigbacc = 0.002588
+ voffcv = -0.16942
+ wpemod = 1
+ dmcgt = 0
+ tcjsw = 0.000357
+ kvth0we = 0.00018
+ lintnoi = -1.5e-8
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ keta = -0.059896633
+ ijthsfwd = 0.01
+ bigsd = 0.00125
+ lags = -3.1905621e-8
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 1.1052395e-9
+ wvoff = 0
+ kt1l = 0
+ tpbswg = 0.0009
+ wvsat = 0
+ wvth0 = -3.2000000000000005e-9
+ ijthsrev = 0.01
+ lint = 6.5375218e-9
+ lkt1 = -4.0479573e-8
+ lkt2 = -1.2823887e-8
+ wtvfbsdoff = 0
+ lmax = 8.9991e-6
+ lmin = 8.9908e-7
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ ptvoff = 0
+ lketa = -9.2926692e-10
+ xpart = 1
+ ltvfbsdoff = 0
+ minv = -0.3
+ lua1 = -3.7234224e-16
+ lub1 = 1.9186851e-25
+ luc1 = 4.1141459e-17
+ nfactor = 1
+ diomod = 1
+ ndep = 1e+18
+ lute = 6.9145309e-9
+ egidl = 0.29734
+ lwlc = 0
+ moin = 5.1
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 2.66208e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.66208e-10
+ nigc = 3.083
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ mjswgd = 0.85
+ mjswgs = 0.85
+ nigbacc = 10
+ ptvfbsdoff = 0
+ tcjswg = 0.001
+ ntox = 1.0
+ pkvth0we = -1.3e-19
+ pcit = -1.2000000000000001e-17
+ pclm = 1.4
+ pvoff = 0
+ nigbinv = 10
+ phin = 0.15
+ cdscb = 0
+ cdscd = 0
+ vfbsdoff = 0.02
+ pvsat = -2.24e-11
+ wk2we = 5e-12
+ pkt1 = 5.600000000000001e-17
+ pvth0 = -1.2e-16
+ drout = 0.56
+ voffl = 0
+ fprout = 300
+ paramchk = 1
+ rbdb = 50
+ prwb = 0
+ prwg = 0
+ pub1 = -3.2e-34
+ xrcrg1 = 12
+ xrcrg2 = 1
+ fnoimod = 1
+ weta0 = 0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ eigbinv = 1.1
+ rdsw = 100
+ )

.model nch_fs_3 nmos (
+ level = 54
+ ku0we = -0.0007
+ beta0 = 13
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ leta0 = 1.6000000000000003e-9
+ ijthsrev = 0.01
+ kvth0we = 0.00018
+ lintnoi = -1.5e-8
+ k2we = 5e-5
+ bigbinv = 0.004953
+ dlcig = 2.5e-9
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ bgidl = 2320000000.0
+ dsub = 0.75
+ wvfbsdoff = 0
+ dtox = 2.7e-10
+ lvfbsdoff = 0
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ eta0 = 0.3
+ dmcgt = 0
+ etab = -0.25
+ tcjsw = 0.000357
+ bigsd = 0.00125
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ wvoff = 0
+ pkvth0we = -1.3e-19
+ nfactor = 1
+ wvsat = 0
+ wvth0 = -3.2000000000000005e-9
+ vfbsdoff = 0.02
+ lketa = -2.6515603e-8
+ toxref = 3e-9
+ xpart = 1
+ nigbacc = 10
+ paramchk = 1
+ egidl = 0.29734
+ nigbinv = 10
+ keta = -0.031147941
+ ltvoff = -6.4393769e-10
+ ijthdfwd = 0.01
+ lags = 4.0889306e-7
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = -1.1851822e-10
+ kt1l = 0
+ lku0we = 2.5e-11
+ fnoimod = 1
+ ijthdrev = 0.01
+ epsrox = 3.9
+ eigbinv = 1.1
+ pvoff = 0
+ lint = 6.5375218e-9
+ cdscb = 0
+ cdscd = 0
+ lkt1 = -1.8244368e-8
+ lkt2 = -1.1493547e-8
+ lmax = 8.9908e-7
+ lpdiblc2 = 3.0380287e-9
+ pvsat = -2.24e-11
+ lmin = 4.4908e-7
+ rdsmod = 0
+ wk2we = 5e-12
+ pvth0 = -1.2e-16
+ drout = 0.56
+ igbmod = 1
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ minv = -0.3
+ voffl = 0
+ lua1 = -1.0281867e-16
+ lub1 = 1.6152992000000002e-26
+ luc1 = 3.7680622e-18
+ pbswgd = 0.95
+ pbswgs = 0.95
+ ndep = 1e+18
+ weta0 = 0
+ lwlc = 0
+ igcmod = 1
+ moin = 5.1
+ a0 = 1.288
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ cigbacc = 0.32875
+ at = 219598.22
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.023410322
+ k3 = -1.8419
+ em = 1000000.0
+ ll = 0
+ nigc = 3.083
+ lw = 0
+ u0 = 0.015110443999999999
+ w0 = 0
+ ua = -1.9429424e-9
+ ub = 2.1566e-18
+ uc = 9.3717778e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ lkvth0we = -2e-12
+ cgidl = 0.22
+ tnoimod = 0
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ cigbinv = 0.006
+ acnqsmod = 0
+ pbswd = 0.8
+ pbsws = 0.8
+ ntox = 1.0
+ pcit = -1.2000000000000001e-17
+ pclm = 1.4
+ pvfbsdoff = 0
+ rbodymod = 0
+ version = 4.5
+ permod = 1
+ phin = 0.15
+ tempmod = 0
+ pdits = 0
+ cigsd = 0.069865
+ pkt1 = 5.600000000000001e-17
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ aigbacc = 0.02
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ voffcv = -0.16942
+ wpemod = 1
+ rbdb = 50
+ prwb = 0
+ pub1 = -3.2e-34
+ prwg = 0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ tnoia = 0
+ rdsw = 100
+ aigbinv = 0.0163
+ peta0 = 0.0
+ tpbsw = 0.0019
+ wtvfbsdoff = 0
+ cjswd = 7.7408e-11
+ cjsws = 7.7408e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ tpbswg = 0.0009
+ rshg = 15.6
+ ltvfbsdoff = 0
+ wkvth0we = 2e-12
+ poxedge = 1
+ trnqsmod = 0
+ ptvoff = 0
+ binunit = 2
+ scref = 1e-6
+ pigcd = 2.621
+ aigsd = 0.01077322
+ tnom = 25
+ diomod = 1
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ ptvfbsdoff = 0
+ lvoff = -1.3784912e-8
+ pditsd = 0
+ rgatemod = 0
+ pditsl = 0
+ cjswgd = 2.66208e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.66208e-10
+ tnjtsswg = 1
+ lvsat = -0.0002
+ lvth0 = 6.9315504e-9
+ delta = 0.007595625
+ laigc = -5.5724245e-11
+ rnoia = 0
+ rnoib = 0
+ mjswgd = 0.85
+ mjswgs = 0.85
+ wags = -8e-9
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ wcit = 4.0000000000000004e-11
+ tcjswg = 0.001
+ ngate = 8e+20
+ voff = -0.1120845
+ acde = 0.4
+ ngcon = 1
+ vsat = 102860
+ wint = 0
+ vth0 = 0.36585892
+ gbmin = 1e-12
+ wkt1 = -2.5600000000000003e-9
+ jswgd = 1.28e-13
+ wmax = 0.00090001
+ jswgs = 1.28e-13
+ aigc = 0.011679696
+ wmin = 8.9974e-6
+ ags = 0.29576959999999997
+ cjd = 0.001281008
+ cit = 0.0013511778
+ cjs = 0.001281008
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 9.8024918e-9
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ fprout = 300
+ dwg = 0
+ dwj = 0
+ njtsswg = 9
+ bigc = 0.001442
+ xrcrg1 = 12
+ xrcrg2 = 1
+ wwlc = 0
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ la0 = -7.832e-8
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.047221618
+ kt1 = -0.22076004
+ kt2 = -0.053318302
+ lk2 = -1.2413537e-8
+ llc = 0
+ cdsc = 0
+ lln = 1
+ lu0 = -1.5393956e-9
+ ckappad = 0.6
+ ckappas = 0.6
+ mjd = 0.26
+ mjs = 0.26
+ lua = -8.9830708e-17
+ lub = -5.4824e-26
+ luc = -1.8883822e-17
+ lud = 0
+ lwc = 0
+ cgbo = 0
+ wtvoff = 0
+ lwl = 0
+ lwn = 1
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ pdiblc1 = 0
+ pdiblc2 = 0.014549485
+ njd = 1.02
+ xtis = 3
+ njs = 1.02
+ pa0 = 0
+ pdiblcb = -0.3
+ nsd = 1e+20
+ pbd = 0.52
+ pat = -3.04e-11
+ pbs = 0.52
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ pu0 = 1.8400000000000002e-18
+ tvoff = 0.0024864064
+ prt = 0
+ pud = 0
+ tvfbsdoff = 0.022
+ rsh = 17.5
+ tcj = 0.00076
+ ijthsfwd = 0.01
+ xjbvd = 1
+ ua1 = 9.685506e-10
+ ub1 = -5.4873129e-19
+ xjbvs = 1
+ uc1 = 6.7696222e-11
+ lk2we = -1.5e-12
+ tpb = 0.0014
+ capmod = 2
+ wa0 = 0
+ ute = -1
+ wat = 0
+ web = 6843.8
+ wec = -25529.0
+ wlc = 0
+ wln = 1
+ wku0we = 2e-11
+ wu0 = -3.6000000000000005e-11
+ xgl = -1.09e-8
+ xgw = 0
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ bigbacc = 0.002588
+ mobmod = 0
+ )

.model nch_fs_4 nmos (
+ level = 54
+ minv = -0.3
+ lua1 = -3.0475764e-17
+ pk2we = -1e-19
+ lub1 = -3.2371927e-26
+ luc1 = -4.3987511e-18
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ ndep = 1e+18
+ rgatemod = 0
+ lwlc = 0
+ moin = 5.1
+ tnjtsswg = 1
+ tnoia = 0
+ nigc = 3.083
+ peta0 = 0.0
+ poxedge = 1
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ tpbsw = 0.0019
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ binunit = 2
+ cjswd = 7.7408e-11
+ cjsws = 7.7408e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ ntox = 1.0
+ pcit = -1.2000000000000001e-17
+ pclm = 1.5439223
+ phin = 0.15
+ pkt1 = 5.600000000000001e-17
+ toxref = 3e-9
+ scref = 1e-6
+ jtsswgd = 2.3e-7
+ pigcd = 2.621
+ jtsswgs = 2.3e-7
+ aigsd = 0.01077322
+ rbdb = 50
+ prwb = 0
+ pub1 = -3.2e-34
+ prwg = 0
+ lvoff = -6.3376134e-9
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ rdsw = 100
+ lvsat = -0.0002
+ lvth0 = -5.170878e-9
+ delta = 0.007595625
+ ltvoff = -1.206053e-10
+ laigc = -1.9935708e-11
+ rnoia = 0
+ rnoib = 0
+ ijthsfwd = 0.01
+ ngate = 8e+20
+ njtsswg = 9
+ ngcon = 1
+ rshg = 15.6
+ lku0we = 2.5e-11
+ ags = -0.025684402000000016
+ epsrox = 3.9
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ cjd = 0.001281008
+ cit = 0.00073144105
+ ijthsrev = 0.01
+ cjs = 0.001281008
+ clc = 1e-7
+ cle = 0.6
+ gbmin = 1e-12
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 1.30529375e-8
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ k3b = 1.9326
+ ckappad = 0.6
+ ckappas = 0.6
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ rdsmod = 0
+ pdiblc1 = 0
+ pdiblc2 = 0.027331777
+ pdiblcb = -0.3
+ igbmod = 1
+ la0 = -2.4730306e-7
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.017025258
+ kt1 = -0.23920434
+ kt2 = -0.070668297
+ lk2 = -9.6174482e-9
+ llc = -1.18e-13
+ lln = 0.7
+ lu0 = -6.147388699999999e-10
+ mjd = 0.26
+ mjs = 0.26
+ lua = -1.0757894e-17
+ lub = -4.7838952e-26
+ luc = -6.6488035e-18
+ lud = 0
+ pbswgd = 0.95
+ pbswgs = 0.95
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ tnom = 25
+ njd = 1.02
+ njs = 1.02
+ pa0 = 0
+ nsd = 1e+20
+ pbd = 0.52
+ pat = -3.04e-11
+ pbs = 0.52
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ pu0 = 1.8400000000000002e-18
+ igcmod = 1
+ prt = 0
+ pud = 0
+ bigbacc = 0.002588
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 8.041349e-10
+ ub1 = -4.3844738e-19
+ uc1 = 8.6257162e-11
+ tpb = 0.0014
+ wa0 = 0
+ ute = -1
+ wat = 0
+ web = 6843.8
+ wec = -25529.0
+ kvth0we = 0.00018
+ wlc = 0
+ wln = 1
+ wu0 = -3.6000000000000005e-11
+ xgl = -1.09e-8
+ xgw = 0
+ tvoff = 0.0012970146
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ tvfbsdoff = 0.022
+ lintnoi = -1.5e-8
+ xjbvd = 1
+ xjbvs = 1
+ wags = -8e-9
+ lk2we = -1.5e-12
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ wcit = 4.0000000000000004e-11
+ voff = -0.12901018
+ acde = 0.4
+ pkvth0we = -1.3e-19
+ ku0we = -0.0007
+ beta0 = 13
+ vsat = 102860
+ wint = 0
+ permod = 1
+ leta0 = 1.6000000000000003e-9
+ vth0 = 0.39336443
+ wkt1 = -2.5600000000000003e-9
+ wmax = 0.00090001
+ aigc = 0.011598359
+ wmin = 8.9974e-6
+ vfbsdoff = 0.02
+ a0 = 1.6720524
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 150970.13
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.017055575
+ k3 = -1.8419
+ em = 1000000.0
+ dlcig = 2.5e-9
+ ll = -1.18e-13
+ wvfbsdoff = 0
+ lw = 0
+ u0 = 0.013008951999999999
+ bgidl = 2320000000.0
+ w0 = 0
+ lvfbsdoff = 0
+ ua = -2.1226533e-9
+ ub = 2.1407249e-18
+ uc = 6.5910917e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ voffcv = -0.16942
+ wpemod = 1
+ bigc = 0.001442
+ paramchk = 1
+ wwlc = 0
+ wtvfbsdoff = 0
+ dmcgt = 0
+ tcjsw = 0.000357
+ nfactor = 1
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ ltvfbsdoff = 0
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ ijthdfwd = 0.01
+ bigsd = 0.00125
+ tpbswg = 0.0009
+ wvoff = 0
+ nigbacc = 10
+ wvsat = 0
+ wvth0 = -3.2000000000000005e-9
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ ijthdrev = 0.01
+ ptvfbsdoff = 0
+ lpdiblc2 = -2.58618e-9
+ ptvoff = 0
+ nigbinv = 10
+ k2we = 5e-5
+ dsub = 0.75
+ lketa = -2.2644187e-8
+ dtox = 2.7e-10
+ xpart = 1
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ diomod = 1
+ pditsd = 0
+ pditsl = 0
+ egidl = 0.29734
+ cjswgd = 2.66208e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.66208e-10
+ eta0 = 0.3
+ etab = -0.25
+ fnoimod = 1
+ eigbinv = 1.1
+ lkvth0we = -2e-12
+ mjswgd = 0.85
+ mjswgs = 0.85
+ tcjswg = 0.001
+ acnqsmod = 0
+ rbodymod = 0
+ pvoff = 0
+ cigbacc = 0.32875
+ cdscb = 0
+ cdscd = 0
+ pvsat = -2.24e-11
+ wk2we = 5e-12
+ pvth0 = -1.2e-16
+ drout = 0.56
+ tnoimod = 0
+ fprout = 300
+ voffl = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ cigbinv = 0.006
+ weta0 = 0
+ lpclm = -6.3325799e-8
+ wtvoff = 0
+ version = 4.5
+ cgidl = 0.22
+ tempmod = 0
+ keta = -0.039946614
+ capmod = 2
+ lags = 5.5033282e-7
+ wku0we = 2e-11
+ aigbacc = 0.02
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 1.5416594e-10
+ pbswd = 0.8
+ mobmod = 0
+ pbsws = 0.8
+ kt1l = 0
+ wkvth0we = 2e-12
+ pvfbsdoff = 0
+ lint = 9.7879675e-9
+ trnqsmod = 0
+ pdits = 0
+ lkt1 = -1.01288734e-8
+ lkt2 = -3.8595493e-9
+ aigbinv = 0.0163
+ lmax = 4.4908e-7
+ cigsd = 0.069865
+ lmin = 2.1577e-7
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ laigsd = -8.1082969e-17
+ )

.model nch_fs_5 nmos (
+ level = 54
+ nigbinv = 10
+ bigsd = 0.00125
+ wags = -8e-9
+ wcit = 4.0000000000000004e-11
+ acnqsmod = 0
+ wvoff = 0
+ voff = -0.15746310460000001
+ acde = 0.4
+ wvsat = 0
+ vsat = 102521.2852
+ wvth0 = -3.2000000000000005e-9
+ rbodymod = 0
+ wint = 0
+ vth0 = 0.4093613742
+ wkt1 = -2.5600000000000003e-9
+ wmax = 0.00090001
+ aigc = 0.011526753
+ wmin = 8.9974e-6
+ fnoimod = 1
+ eigbinv = 1.1
+ toxref = 3e-9
+ lketa = -1.1430034e-8
+ xpart = 1
+ bigc = 0.001442
+ wwlc = 0
+ egidl = 0.29734
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ ltvoff = 1.4850105e-11
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ cigbacc = 0.32875
+ tnoimod = 0
+ lku0we = 2.5e-11
+ cigbinv = 0.006
+ epsrox = 3.9
+ wkvth0we = 2e-12
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ pvoff = 0
+ rdsmod = 0
+ trnqsmod = 0
+ cdscb = 0
+ cdscd = 0
+ igbmod = 1
+ pvsat = -2.24e-11
+ version = 4.5
+ wk2we = 5e-12
+ pvth0 = -1.2e-16
+ k2we = 5e-5
+ drout = 0.56
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ tempmod = 0
+ dsub = 0.75
+ dtox = 2.7e-10
+ pbswgd = 0.95
+ pbswgs = 0.95
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ voffl = 0
+ igcmod = 1
+ aigbacc = 0.02
+ weta0 = 0
+ eta0 = 0.3
+ rgatemod = 0
+ etab = -0.25
+ lpclm = -2.4377173e-8
+ tnjtsswg = 1
+ cgidl = 0.22
+ aigbinv = 0.0163
+ pbswd = 0.8
+ pbsws = 0.8
+ pvfbsdoff = 0
+ permod = 1
+ wtvfbsdoff = 0
+ pdits = 0
+ cigsd = 0.069865
+ dvt0w = 0
+ dvt1w = 0
+ poxedge = 1
+ dvt2w = 0
+ ltvfbsdoff = 0
+ voffcv = -0.16942
+ wpemod = 1
+ binunit = 2
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ tnoia = 0
+ peta0 = 0.0
+ wketa = 0
+ keta = -0.093093889
+ ptvfbsdoff = 0
+ tpbsw = 0.0019
+ ijthsfwd = 0.01
+ cjswd = 7.7408e-11
+ cjsws = 7.7408e-11
+ a0 = 0.66068814
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ mjswd = 0.11
+ lags = 3.3904274e-13
+ mjsws = 0.11
+ agidl = 9.41e-8
+ tpbswg = 0.0009
+ at = 79499.116
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = -0.017712078
+ k3 = -1.8419
+ em = 1000000.0
+ jswd = 1.28e-13
+ ll = -1.18e-13
+ jsws = 1.28e-13
+ lw = 0
+ u0 = 0.011006872
+ w0 = 0
+ lcit = 7.6591162e-11
+ ua = -2.2893587e-9
+ ub = 2.089788886e-18
+ uc = 4.5969231e-11
+ ud = 0
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ kt1l = 0
+ ijthsrev = 0.01
+ lint = 9.7879675e-9
+ ptvoff = 0
+ lkt1 = -3.787522600000001e-9
+ lkt2 = -6.0180086e-10
+ lmax = 2.1577e-7
+ lmin = 9e-8
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ scref = 1e-6
+ diomod = 1
+ pigcd = 2.621
+ minv = -0.3
+ aigsd = 0.01077322
+ lua1 = 7.6861327e-18
+ lub1 = -5.4742256e-26
+ luc1 = -4.2210821e-18
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 2.66208e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.66208e-10
+ ndep = 1e+18
+ lvoff = -3.340626e-10
+ njtsswg = 9
+ lwlc = 0
+ moin = 5.1
+ lvsat = -0.00012851569999999997
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ lvth0 = -8.5462159e-9
+ nigc = 3.083
+ delta = 0.007595625
+ mjswgd = 0.85
+ mjswgs = 0.85
+ laigc = -4.8268328e-12
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.02163037
+ pdiblcb = -0.3
+ tcjswg = 0.001
+ rnoia = 0
+ rnoib = 0
+ ags = 2.5825264
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ cjd = 0.001281008
+ cit = 0.001099094
+ cjs = 0.001281008
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 1.30529375e-8
+ pketa = 0
+ ngate = 8e+20
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ ngcon = 1
+ pkvth0we = -1.3e-19
+ ntox = 1.0
+ pcit = -1.2000000000000001e-17
+ pclm = 1.3593316
+ bigbacc = 0.002588
+ la0 = -3.3904685e-8
+ gbmin = 1e-12
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.0019448735
+ kt1 = -0.26925814
+ kt2 = -0.086107863
+ lk2 = -2.2814734e-9
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ llc = -1.18e-13
+ lln = 0.7
+ phin = 0.15
+ lu0 = -1.9229995e-10
+ mjd = 0.26
+ mjs = 0.26
+ lua = 2.4416942e-17
+ lub = -3.7091512499999996e-26
+ luc = -2.4411077e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ vfbsdoff = 0.02
+ njd = 1.02
+ njs = 1.02
+ pa0 = 0
+ nsd = 1e+20
+ kvth0we = 0.00018
+ pbd = 0.52
+ pat = -3.04e-11
+ pbs = 0.52
+ pkt1 = 5.600000000000001e-17
+ pu0 = 1.8400000000000002e-18
+ prt = 0
+ fprout = 300
+ pub = 0
+ pud = 0
+ lintnoi = -1.5e-8
+ rsh = 17.5
+ xrcrg1 = 12
+ xrcrg2 = 1
+ tcj = 0.00076
+ ua1 = 6.2327283e-10
+ ub1 = -3.3242687e-19
+ uc1 = 8.5415128e-11
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ tpb = 0.0014
+ wa0 = 0
+ ute = -1
+ paramchk = 1
+ wat = 0
+ web = 6843.8
+ wec = -25529.0
+ wlc = 0
+ wln = 1
+ wu0 = -3.6000000000000005e-11
+ rbdb = 50
+ xgl = -1.09e-8
+ prwb = 0
+ pub1 = -3.2e-34
+ prwg = 0
+ xgw = 0
+ wub = 0
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ rbpb = 50
+ rbpd = 50
+ wtvoff = 0
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ rdsw = 100
+ tvfbsdoff = 0.022
+ tvoff = 0.00065504585
+ capmod = 2
+ ijthdfwd = 0.01
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ wku0we = 2e-11
+ mobmod = 0
+ rshg = 15.6
+ ku0we = -0.0007
+ beta0 = 13
+ leta0 = 1.6000000000000003e-9
+ ijthdrev = 0.01
+ nfactor = 1
+ lpdiblc2 = -1.3831831e-9
+ wvfbsdoff = 0
+ dlcig = 2.5e-9
+ lvfbsdoff = 0
+ bgidl = 2320000000.0
+ laigsd = 3.3904273e-17
+ tnom = 25
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ nigbacc = 10
+ dmcgt = 0
+ tcjsw = 0.000357
+ lkvth0we = -2e-12
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ )

.model nch_fs_6 nmos (
+ level = 54
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ vfbsdoff = 0.02
+ toxref = 3e-9
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.0069155858
+ scref = 1e-6
+ pdiblcb = -0.3
+ pigcd = 2.621
+ aigsd = 0.01077322
+ paramchk = 1
+ lvoff = -2.08041089e-9
+ ags = 2.5825299999999998
+ lvsat = 0.0010635378699999998
+ ltvoff = 1.0839662e-10
+ lvth0 = 1.7692931699999999e-9
+ bigbacc = 0.002588
+ cjd = 0.001281008
+ cit = 0.00031861111
+ cjs = 0.001281008
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ delta = 0.007595625
+ dlc = 3.26497e-9
+ k3b = 1.9326
+ laigc = -2.2427226e-11
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ keta = -0.52835722
+ rnoia = 0
+ rnoib = 0
+ ijthdfwd = 0.01
+ kvth0we = 0.00018
+ la0 = 3.0288889e-8
+ jsd = 6.11e-7
+ lintnoi = -1.5e-8
+ jss = 6.11e-7
+ lat = -0.00054029214
+ kt1 = -0.40872879
+ kt2 = -0.10088778
+ lk2 = -4.8654938e-10
+ lku0we = 2.5e-11
+ pketa = 0
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ ngate = 8e+20
+ bigbinv = 0.004953
+ llc = 0
+ lln = 1
+ lu0 = 1.1243078e-10
+ lcit = 1.4995656e-10
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ mjd = 0.26
+ mjs = 0.26
+ lua = 3.5218789e-17
+ lub = -1.9869262700000004e-26
+ luc = 2.2716666e-18
+ lud = 0
+ epsrox = 3.9
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ ngcon = 1
+ njd = 1.02
+ njs = 1.02
+ kt1l = 0
+ pa0 = 0
+ nsd = 1e+20
+ pbd = 0.52
+ pat = -3.04e-11
+ pbs = 0.52
+ pu0 = 1.8400000000000002e-18
+ prt = 0
+ pub = 0
+ puc = 0
+ pud = 0
+ rdsmod = 0
+ ijthdrev = 0.01
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ rsh = 17.5
+ jswgs = 1.28e-13
+ lint = 0
+ tcj = 0.00076
+ igbmod = 1
+ ua1 = 8.897383e-10
+ ub1 = -8.0235504e-19
+ uc1 = -6.3390556e-11
+ tpb = 0.0014
+ lkt1 = 9.3227184e-9
+ lkt2 = 7.8751111e-10
+ wa0 = 0
+ lpdiblc2 = 6.6256944e-15
+ lmax = 9e-8
+ ute = -1
+ wat = 0
+ web = 6843.8
+ pscbe1 = 1000000000.0
+ wec = -25529.0
+ pscbe2 = 1e-20
+ lmin = 5.4e-8
+ wlc = 0
+ wln = 1
+ wu0 = -3.6000000000000005e-11
+ xgl = -1.09e-8
+ xgw = 0
+ wub = 0
+ wuc = 0
+ wud = 0
+ lpe0 = 9.2e-8
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ pbswgd = 0.95
+ lpeb = 2.5e-7
+ pbswgs = 0.95
+ minv = -0.3
+ igcmod = 1
+ lua1 = -1.7361621e-17
+ lub1 = -1.05690078e-26
+ luc1 = 9.7666522e-18
+ ndep = 1e+18
+ lwlc = 0
+ moin = 5.1
+ nigc = 3.083
+ tvfbsdoff = 0.022
+ nfactor = 1
+ lkvth0we = -2e-12
+ tvoff = -0.00034012981
+ wtvfbsdoff = 0
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ acnqsmod = 0
+ ltvfbsdoff = 0
+ permod = 1
+ ntox = 1.0
+ pcit = -1.2000000000000001e-17
+ ku0we = -0.0007
+ pclm = 1.2209944
+ beta0 = 13
+ rbodymod = 0
+ leta0 = 4.628888900000001e-9
+ nigbacc = 10
+ letab = -2.2684433e-8
+ phin = 0.15
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ pkt1 = 5.600000000000001e-17
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ voffcv = -0.16942
+ wpemod = 1
+ nigbinv = 10
+ ptvfbsdoff = 0
+ rbdb = 50
+ prwb = 0
+ pub1 = -3.2e-34
+ prwg = 0
+ dmcgt = 0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ tcjsw = 0.000357
+ rdsw = 100
+ fnoimod = 1
+ eigbinv = 1.1
+ bigsd = 0.00125
+ tpbswg = 0.0009
+ wvoff = 0
+ rshg = 15.6
+ wkvth0we = 2e-12
+ wvsat = 0.0
+ wvth0 = -3.2000000000000005e-9
+ ptvoff = 0
+ trnqsmod = 0
+ cigbacc = 0.32875
+ diomod = 1
+ lketa = 2.9484719e-8
+ xpart = 1
+ pditsd = 0
+ pditsl = 0
+ tnoimod = 0
+ cjswgd = 2.66208e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.66208e-10
+ tnom = 25
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ egidl = 0.29734
+ a0 = -0.02222221999999996
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ rgatemod = 0
+ at = 64556.761
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = -0.036807015
+ k3 = -1.8419
+ em = 1000000.0
+ cigbinv = 0.006
+ ll = 0
+ lw = 0
+ u0 = 0.0077650556
+ tnjtsswg = 1
+ w0 = 0
+ ua = -2.404272e-9
+ ub = 1.906573466e-18
+ uc = -4.166667e-12
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ mjswgd = 0.85
+ mjswgs = 0.85
+ tcjswg = 0.001
+ version = 4.5
+ wags = -8e-9
+ tempmod = 0
+ wcit = 4.0000000000000004e-11
+ voff = -0.138884931
+ acde = 0.4
+ aigbacc = 0.02
+ vsat = 89839.86
+ wint = 0
+ vth0 = 0.299621916
+ pvoff = 0
+ wkt1 = -2.5600000000000003e-9
+ wmax = 0.00090001
+ aigc = 0.011713991
+ wmin = 8.9974e-6
+ cdscb = 0
+ cdscd = 0
+ pvsat = -2.24e-11
+ wk2we = 5e-12
+ pvth0 = -1.2e-16
+ fprout = 300
+ drout = 0.56
+ xrcrg1 = 12
+ xrcrg2 = 1
+ aigbinv = 0.0163
+ voffl = 0
+ bigc = 0.001442
+ wwlc = 0
+ wtvoff = 0
+ weta0 = 0
+ lpclm = -1.1373478e-8
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ cgidl = 0.22
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ capmod = 2
+ wku0we = 2e-11
+ ijthsfwd = 0.01
+ poxedge = 1
+ mobmod = 0
+ pbswd = 0.8
+ pvfbsdoff = 0
+ pbsws = 0.8
+ binunit = 2
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ ijthsrev = 0.01
+ pdits = 0
+ cigsd = 0.069865
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ k2we = 5e-5
+ dsub = 0.75
+ dtox = 2.7e-10
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ eta0 = 0.26777778
+ etab = -0.0086762422
+ tnoia = 0
+ peta0 = 0.0
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ wketa = 0
+ tpbsw = 0.0019
+ cjswd = 7.7408e-11
+ cjsws = 7.7408e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ pkvth0we = -1.3e-19
+ njtsswg = 9
+ )

.model nch_fs_7 nmos (
+ level = 54
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ ltvoff = -2.4740506e-10
+ aigbacc = 0.02
+ rdsw = 100
+ ijthsfwd = 0.01
+ lku0we = 2.5e-11
+ aigbinv = 0.0163
+ epsrox = 3.9
+ rshg = 15.6
+ rdsmod = 0
+ igbmod = 1
+ ijthsrev = 0.01
+ pvoff = 0
+ cdscb = 0
+ cdscd = 0
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ pvsat = -2.24e-11
+ wk2we = 5e-12
+ pvth0 = -1.2e-16
+ drout = 0.56
+ pbswgd = 0.95
+ pbswgs = 0.95
+ igcmod = 1
+ poxedge = 1
+ wtvfbsdoff = 0
+ voffl = 0
+ tnom = 25
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ weta0 = 0
+ binunit = 2
+ lpclm = -7.2871722e-8
+ ltvfbsdoff = 0
+ cgidl = 0.22
+ wags = -8e-9
+ wcit = 4.0000000000000004e-11
+ pvfbsdoff = 0
+ permod = 1
+ pbswd = 0.8
+ pbsws = 0.8
+ voff = -0.112415764
+ pkvth0we = -1.3e-19
+ acde = 0.4
+ ptvfbsdoff = 0
+ vsat = 73870.58200000001
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ wint = 0
+ vth0 = 0.297517597
+ wkt1 = -2.5600000000000003e-9
+ wmax = 0.00090001
+ aigc = 0.011692671
+ pdits = 0
+ wmin = 8.9974e-6
+ vfbsdoff = 0.02
+ cigsd = 0.069865
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ voffcv = -0.16942
+ wpemod = 1
+ wub1 = 0.0
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ bigc = 0.001442
+ paramchk = 1
+ wwlc = 0
+ tnoia = 0
+ cdsc = 0
+ cgbo = 0
+ njtsswg = 9
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ peta0 = 0.0
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ tpbsw = 0.0019
+ ijthdfwd = 0.01
+ tpbswg = 0.0009
+ ckappad = 0.6
+ cjswd = 7.7408e-11
+ ckappas = 0.6
+ cjsws = 7.7408e-11
+ mjswd = 0.11
+ pdiblc1 = 0
+ pdiblc2 = 0.0069157
+ mjsws = 0.11
+ agidl = 9.41e-8
+ pdiblcb = -0.3
+ ptvoff = 0
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ ijthdrev = 0.01
+ bigbacc = 0.002588
+ diomod = 1
+ k2we = 5e-5
+ dsub = 0.75
+ scref = 1e-6
+ dtox = 2.7e-10
+ pditsd = 0
+ pditsl = 0
+ kvth0we = 0.00018
+ cjswgd = 2.66208e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.66208e-10
+ ags = 2.5825299999999998
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ pigcd = 2.621
+ aigsd = 0.01077322
+ cjd = 0.001281008
+ cit = -0.0027423847
+ cjs = 0.001281008
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ lintnoi = -1.5e-8
+ dlc = 3.26497e-9
+ bigbinv = 0.004953
+ k3b = 1.9326
+ lvoff = -3.6156221999999994e-9
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ eta0 = 0.35179556
+ etab = -1.0973583
+ lvsat = 0.0019897560999999997
+ mjswgd = 0.85
+ mjswgs = 0.85
+ lvth0 = 1.8913432999999988e-9
+ la0 = -3.1577778e-7
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = 0.0074186667
+ lkvth0we = -2e-12
+ kt1 = 0.010917511
+ kt2 = -0.10990444
+ lk2 = -1.5787889e-9
+ delta = 0.007595625
+ tcjswg = 0.001
+ llc = 0
+ laigc = -2.1190647e-11
+ lln = 1
+ lu0 = 5.565271100000001e-10
+ mjd = 0.26
+ mjs = 0.26
+ lua = 7.8730998e-17
+ lub = -4.3148946000000005e-26
+ luc = 1.578889e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 0
+ rnoia = 0
+ rnoib = 0
+ nsd = 1e+20
+ pbd = 0.52
+ pat = -3.04e-11
+ pbs = 0.52
+ pu0 = 1.8400000000000002e-18
+ prt = 0
+ pub = 0
+ puc = 0
+ pud = 0
+ acnqsmod = 0
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 3.744227e-10
+ ngate = 8e+20
+ ub1 = -1.4506222e-18
+ uc1 = -1.6722222e-10
+ tpb = 0.0014
+ ngcon = 1
+ wa0 = 0
+ ute = -1
+ wat = 0.0
+ web = 6843.8
+ wec = -25529.0
+ wlc = 0
+ wln = 1
+ wu0 = -3.6000000000000005e-11
+ xgl = -1.09e-8
+ xgw = 0
+ wub = 0
+ wuc = 0
+ wud = 0
+ rbodymod = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ a0 = 5.9444444
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = -72666.667
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = -0.017975299
+ k3 = -1.8419
+ em = 1000000.0
+ fprout = 300
+ ll = 0
+ lw = 0
+ u0 = 0.00010822221999999998
+ nfactor = 1
+ w0 = 0
+ ua = -3.1544825e-9
+ ub = 2.30794738e-18
+ uc = 7.77778e-12
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ xrcrg1 = 12
+ xrcrg2 = 1
+ wtvoff = 0
+ tvfbsdoff = 0.022
+ nigbacc = 10
+ capmod = 2
+ tvoff = 0.0057943818
+ wku0we = 2e-11
+ keta = 0.088888889
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ mobmod = 0
+ nigbinv = 10
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 3.2749431e-10
+ kt1l = 0
+ ku0we = -0.0007
+ wkvth0we = 2e-12
+ beta0 = 13
+ leta0 = -2.441421999999998e-10
+ letab = 4.0459126e-8
+ lint = 0
+ trnqsmod = 0
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ lkt1 = -1.5016767e-8
+ lkt2 = 1.3104778e-9
+ lmax = 5.4e-8
+ lmin = 4.5e-8
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ lpe0 = 9.2e-8
+ fnoimod = 1
+ lpeb = 2.5e-7
+ eigbinv = 1.1
+ minv = -0.3
+ lua1 = 1.2526683e-17
+ lub1 = 2.7030489e-26
+ luc1 = 1.5788889e-17
+ ndep = 1e+18
+ dmcgt = 0
+ rgatemod = 0
+ lwlc = 0
+ tcjsw = 0.000357
+ moin = 5.1
+ tnjtsswg = 1
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ nigc = 3.083
+ bigsd = 0.00125
+ noff = 2.7195
+ cigbacc = 0.32875
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ wvoff = 0
+ tnoimod = 0
+ ntox = 1.0
+ pcit = -1.2000000000000001e-17
+ pclm = 2.281309
+ wvsat = 0.0
+ wvth0 = -3.2000000000000005e-9
+ cigbinv = 0.006
+ phin = 0.15
+ toxref = 3e-9
+ pkt1 = 5.600000000000001e-17
+ lketa = -6.3155556e-9
+ version = 4.5
+ xpart = 1
+ tempmod = 0
+ egidl = 0.29734
+ rbdb = 50
+ prwb = 0
+ pub1 = -3.2e-34
+ prwg = 0
+ )

.model nch_fs_8 nmos (
+ level = 54
+ ngate = 8e+20
+ ngcon = 1
+ wpclm = 0
+ rdsmod = 0
+ wkvth0we = 2e-12
+ wtvfbsdoff = 0
+ igbmod = 1
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ trnqsmod = 0
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ nigbacc = 10
+ ltvfbsdoff = 0
+ pbswgd = 0.95
+ pbswgs = 0.95
+ k2we = 5e-5
+ igcmod = 1
+ dsub = 0.75
+ dtox = 2.7e-10
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ nigbinv = 10
+ rgatemod = 0
+ eta0 = -0.001232
+ etab = -0.88502038
+ tnjtsswg = 1
+ tvfbsdoff = 0.022
+ ptvfbsdoff = 0
+ tvoff = 0.0030235155
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ fnoimod = 1
+ permod = 1
+ eigbinv = 1.1
+ ku0we = -0.0007
+ beta0 = 13
+ leta0 = 1.7054208000000002e-8
+ letab = 3.0054568e-8
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ ppclm = 0
+ voffcv = -0.16942
+ wpemod = 1
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ cigbacc = 0.32875
+ dmcgt = 0
+ tnoimod = 0
+ tcjsw = 0.000357
+ cigbinv = 0.006
+ tpbswg = 0.0009
+ keta = 0.44888889
+ ijthsfwd = 0.01
+ bigsd = 0.00125
+ version = 4.5
+ wvoff = 0
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 4.4836639e-10
+ tempmod = 0
+ kt1l = 0
+ ptvoff = 0
+ wvsat = 0.0
+ wvth0 = -3.2000000000000005e-9
+ ijthsrev = 0.01
+ lint = 0
+ aigbacc = 0.02
+ lkt1 = -4.3888498e-9
+ lkt2 = 1.6072e-9
+ diomod = 1
+ lmax = 4.5e-8
+ lmin = 3.6e-8
+ lpe0 = 9.2e-8
+ pditsd = 0
+ pditsl = 0
+ lketa = -2.3955556e-8
+ lpeb = 2.5e-7
+ cjswgd = 2.66208e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.66208e-10
+ xpart = 1
+ minv = -0.3
+ aigbinv = 0.0163
+ lua1 = 7.1708778e-18
+ lub1 = -2.6342999000000003e-26
+ luc1 = -1.63268e-17
+ egidl = 0.29734
+ ndep = 1e+18
+ lwlc = 0
+ mjswgd = 0.85
+ mjswgs = 0.85
+ moin = 5.1
+ nigc = 3.083
+ tcjswg = 0.001
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ poxedge = 1
+ pkvth0we = -1.3e-19
+ ntox = 1.0
+ pcit = -1.2000000000000001e-17
+ pclm = 2.10165423
+ binunit = 2
+ pvoff = 0
+ fprout = 300
+ phin = 0.15
+ cdscb = 0
+ cdscd = 0
+ vfbsdoff = 0.02
+ pvsat = -2.24e-11
+ xrcrg1 = 12
+ xrcrg2 = 1
+ wk2we = 5e-12
+ pvth0 = -1.2e-16
+ drout = 0.56
+ pkt1 = 5.600000000000001e-17
+ voffl = 0
+ wtvoff = 0
+ paramchk = 1
+ weta0 = 0
+ rbdb = 50
+ prwb = 0
+ pub1 = -3.2e-34
+ prwg = 0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ lpclm = -6.406864000000001e-8
+ rdsw = 100
+ capmod = 2
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ cgidl = 0.22
+ wku0we = 2e-11
+ mobmod = 0
+ ijthdfwd = 0.01
+ a0 = 3.6555556
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 123237.73
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.022556861
+ k3 = -1.8419
+ em = 1000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.0030922232999999995
+ pvfbsdoff = 0
+ w0 = 0
+ ua = -2.2580401200000003e-9
+ ub = 1.5627388499999998e-18
+ uc = 2.4e-10
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ pbswd = 0.8
+ pbsws = 0.8
+ rshg = 15.6
+ ijthdrev = 0.01
+ pdits = 0
+ njtsswg = 9
+ cigsd = 0.069865
+ laigsd = -2.1777778e-17
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ ckappad = 0.6
+ ckappas = 0.6
+ pk2we = -1e-19
+ tnom = 25
+ pdiblc1 = 0
+ pdiblc2 = 0.0069157
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ pdiblcb = -0.3
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ tnoia = 0
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ peta0 = 0.0
+ lkvth0we = -2e-12
+ bigbacc = 0.002588
+ tpbsw = 0.0019
+ wags = -8e-9
+ cjswd = 7.7408e-11
+ cjsws = 7.7408e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ wcit = 4.0000000000000004e-11
+ kvth0we = 0.00018
+ acnqsmod = 0
+ voff = -0.039834349000000005
+ acde = 0.4
+ lintnoi = -1.5e-8
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ vsat = 85481.92200000002
+ rbodymod = 0
+ vtsswgs = 4.2
+ wint = 0
+ vth0 = 0.34578350300000005
+ toxref = 3e-9
+ wkt1 = -2.5600000000000003e-9
+ ags = 2.5825299999999998
+ wmax = 0.00090001
+ aigc = 0.011387162
+ wmin = 8.9974e-6
+ cjd = 0.001281008
+ cit = -0.0052091698
+ cjs = 0.001281008
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 3.26497e-9
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ scref = 1e-6
+ wub1 = 0.0
+ pigcd = 2.621
+ aigsd = 0.010773221
+ la0 = -2.0362223e-7
+ bigc = 0.001442
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.0021806488
+ kt1 = -0.20597876
+ kt2 = -0.11596
+ lk2 = -3.5648647e-9
+ wwlc = 0
+ llc = 0
+ lvoff = -7.1721119000000006e-9
+ lln = 1
+ lu0 = 4.1031107e-10
+ mjd = 0.26
+ mjs = 0.26
+ lua = 3.4805321000000004e-17
+ lub = -6.633731000000002e-27
+ luc = -9.7999999e-18
+ lud = 0
+ ltvoff = -1.1163261e-10
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 0
+ nsd = 1e+20
+ pbd = 0.52
+ pat = -3.04e-11
+ pbs = 0.52
+ pk2 = 0
+ lvsat = 0.00142080039
+ cdsc = 0
+ pu0 = 1.8400000000000002e-18
+ lvth0 = -4.736881199999997e-10
+ prt = 0
+ cgbo = 0
+ pua = 0
+ pub = 0
+ puc = 0
+ pud = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ delta = 0.007595625
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 4.8372486e-10
+ ub1 = -3.6136738e-19
+ cigc = 0.000625
+ laigc = -6.2207351e-12
+ uc1 = 4.882e-10
+ tpb = 0.0014
+ wa0 = 0
+ rnoia = 0
+ rnoib = 0
+ nfactor = 1
+ ute = -1
+ wat = 0.0
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 0
+ wlc = 0
+ lku0we = 2.5e-11
+ wln = 1
+ wu0 = -3.6000000000000005e-11
+ xgl = -1.09e-8
+ xgw = 0
+ wua = 0
+ wub = 0
+ wuc = 0
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ epsrox = 3.9
+ )

.model nch_fs_9 nmos (
+ level = 54
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ ptvfbsdoff = 0
+ voffl = 0
+ minv = -0.3
+ lub1 = -2.4000000000000004e-27
+ weta0 = 0
+ ndep = 1e+18
+ wetab = -1.0073378e-8
+ lwlc = 0
+ moin = 5.1
+ nigc = 3.083
+ cgidl = 0.22
+ lkvth0we = -2e-12
+ njtsswg = 9
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ pvfbsdoff = 0
+ noic = 45200000.0
+ permod = 1
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ acnqsmod = 0
+ pbswd = 0.8
+ pbsws = 0.8
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.018557155
+ pdiblcb = -0.3
+ ntox = 1.0
+ pcit = -1.2000000000000001e-17
+ pclm = 1.4152454
+ rbodymod = 0
+ phin = 0.15
+ voffcv = -0.16942
+ wpemod = 1
+ pdits = 0
+ cigsd = 0.069865
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ pkt1 = 5.600000000000001e-17
+ bigbacc = 0.002588
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ kvth0we = 0.00018
+ rbdb = 50
+ prwb = 0
+ pub1 = -3.2e-34
+ prwg = 0
+ wpdiblc2 = -1.7177628e-11
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ lintnoi = -1.5e-8
+ tnoia = 0
+ bigbinv = 0.004953
+ rdsw = 100
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ peta0 = 0.0
+ tpbswg = 0.0009
+ wketa = 3.3422159e-8
+ tpbsw = 0.0019
+ cjswd = 7.7408e-11
+ cjsws = 7.7408e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ ags = 0.7968331399999999
+ ptvoff = 0
+ cjd = 0.001281008
+ cit = 4.8708935e-5
+ cjs = 0.001281008
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ wkvth0we = 2e-12
+ bvs = 8.7
+ rshg = 15.6
+ waigsd = 3.0716751e-12
+ dlc = 9.8024918e-9
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ trnqsmod = 0
+ diomod = 1
+ la0 = 0
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.00016
+ kt1 = -0.19515831
+ kt2 = -0.052853133
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 2.66208e-10
+ llc = 0
+ pku0we = -1.5e-18
+ lln = 1
+ cjswgs = 2.66208e-10
+ lu0 = 9.600000000000001e-12
+ mjd = 0.26
+ mjs = 0.26
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ scref = 1e-6
+ njd = 1.02
+ njs = 1.02
+ pa0 = 0
+ nfactor = 1
+ nsd = 1e+20
+ pbd = 0.52
+ pat = -3.04e-11
+ pbs = 0.52
+ pigcd = 2.621
+ aigsd = 0.010772879
+ pu0 = 1.8400000000000002e-18
+ prt = 0
+ pud = 0
+ tnom = 25
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 1.311952e-9
+ toxe = 2.43e-9
+ ub1 = -8.0649865e-19
+ toxm = 2.43e-9
+ lvoff = -1.6e-11
+ uc1 = 3.0375074e-11
+ mjswgd = 0.85
+ mjswgs = 0.85
+ tpb = 0.0014
+ rgatemod = 0
+ wa0 = -2.5183444e-7
+ ute = -0.96248296
+ wat = 0
+ tnjtsswg = 1
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -3.7920026e-9
+ lvsat = -0.0002
+ wlc = 0
+ tcjswg = 0.001
+ wln = 1
+ wu0 = -2.9790781999999996e-10
+ xgl = -1.09e-8
+ xgw = 0
+ lvth0 = -4.8e-10
+ wua = -4.0765791e-17
+ wub = 4.0599742e-26
+ wuc = -7.8572347e-18
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ delta = 0.007595625
+ nigbacc = 10
+ rnoia = 0
+ rnoib = 0
+ wags = -9.2054279e-8
+ wcit = 5.0192733e-10
+ ngate = 8e+20
+ voff = -0.11308442
+ ngcon = 1
+ wpclm = -1.3730014e-7
+ acde = 0.4
+ nigbinv = 10
+ vsat = 103058.98
+ wint = 0
+ gbmin = 1e-12
+ vth0 = 0.32314845
+ fprout = 300
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ wkt1 = -4.8199654e-8
+ wkt2 = -3.5741805e-9
+ wmax = 8.9974e-6
+ xrcrg1 = 12
+ xrcrg2 = 1
+ aigc = 0.011766468
+ wmin = 8.974e-7
+ wtvoff = -8.3463378e-10
+ wua1 = -7.3834184e-16
+ wub1 = 7.3798399e-25
+ wuc1 = -8.5623711e-19
+ fnoimod = 1
+ bigc = 0.001442
+ wute = -4.0092044e-7
+ eigbinv = 1.1
+ wwlc = 0
+ tvfbsdoff = 0.022
+ capmod = 2
+ cdsc = 0
+ cgbo = 0
+ wku0we = 2e-11
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ tvoff = 0.0020036382
+ cigc = 0.000625
+ mobmod = 0
+ xjbvd = 1
+ ijthsfwd = 0.01
+ xjbvs = 1
+ lk2we = -1.5e-12
+ cigbacc = 0.32875
+ ku0we = -0.0007
+ beta0 = 13
+ leta0 = 1.6000000000000003e-9
+ tnoimod = 0
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ ijthsrev = 0.01
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ cigbinv = 0.006
+ dlcig = 2.5e-9
+ k2we = 5e-5
+ bgidl = 2320000000.0
+ dsub = 0.75
+ dtox = 2.7e-10
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ a0 = 3.277963
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ version = 4.5
+ at = 72000
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.023422307
+ k3 = -1.8419
+ em = 1000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.015419081999999999
+ dmcgt = 0
+ w0 = 0
+ tempmod = 0
+ ua = -1.8192461e-9
+ ub = 2.0991879e-18
+ uc = 7.4172444e-11
+ ud = 0
+ eta0 = 0.3
+ tcjsw = 0.000357
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ alpha0 = 2e-10
+ ww = 0
+ alpha1 = 3.6
+ xw = 8.600000000000001e-9
+ etab = -0.24888148
+ aigbacc = 0.02
+ bigsd = 0.00125
+ wvoff = 2.3777201e-9
+ pkvth0we = -1.3e-19
+ aigbinv = 0.0163
+ wvsat = -0.0017920539
+ wvth0 = -1.4345485000000001e-8
+ toxref = 3e-9
+ waigc = 2.6350949e-11
+ vfbsdoff = 0.02
+ xpart = 1
+ paramchk = 1
+ ltvoff = 0
+ egidl = 0.29734
+ poxedge = 1
+ binunit = 2
+ wtvfbsdoff = 0
+ keta = -0.063711099
+ lku0we = 2.5e-11
+ ijthdfwd = 0.01
+ epsrox = 3.9
+ ltvfbsdoff = 0
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = -8e-12
+ rdsmod = 0
+ kt1l = 0
+ igbmod = 1
+ ijthdrev = 0.01
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ pvoff = 0
+ lint = 6.5375218e-9
+ pbswgd = 0.95
+ cdscb = 0
+ cdscd = 0
+ pbswgs = 0.95
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ lkt1 = -4.8e-10
+ pvsat = -2.24e-11
+ lmax = 2.001e-5
+ wk2we = 5e-12
+ pvth0 = -1.2e-16
+ lmin = 8.9991e-6
+ drout = 0.56
+ igcmod = 1
+ )

.model nch_fs_10 nmos (
+ level = 54
+ xrcrg1 = 12
+ xrcrg2 = 1
+ cgidl = 0.22
+ vfbsdoff = 0.02
+ wtvoff = -8.9580408e-10
+ nfactor = 1
+ pbswd = 0.8
+ pbsws = 0.8
+ paramchk = 1
+ capmod = 2
+ wku0we = 2e-11
+ mobmod = 0
+ pdits = 0
+ cigsd = 0.069865
+ nigbacc = 10
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ ijthdfwd = 0.01
+ keta = -0.064075044
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ nigbinv = 10
+ lags = -6.3328546e-8
+ wtvfbsdoff = 0
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 1.1257416e-9
+ tnoia = 0
+ laigsd = 1.1048614e-17
+ ijthdrev = 0.01
+ kt1l = 0
+ peta0 = 0.0
+ ltvfbsdoff = 0
+ lpdiblc2 = -6.1589259e-10
+ wketa = 3.7630763e-8
+ lint = 6.5375218e-9
+ tpbsw = 0.0019
+ lkt1 = -4.6017316e-8
+ lkt2 = -1.2972142e-8
+ cjswd = 7.7408e-11
+ lmax = 8.9991e-6
+ cjsws = 7.7408e-11
+ lmin = 8.9908e-7
+ fnoimod = 1
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ lpe0 = 9.2e-8
+ eigbinv = 1.1
+ lpeb = 2.5e-7
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ minv = -0.3
+ lua1 = -4.3996966e-16
+ lub1 = 2.5820002e-25
+ luc1 = 3.9191378e-17
+ ndep = 1e+18
+ lute = -3.7058959e-8
+ lwlc = 0
+ ptvfbsdoff = 0
+ moin = 5.1
+ lkvth0we = -2e-12
+ nigc = 3.083
+ scref = 1e-6
+ pigcd = 2.621
+ aigsd = 0.010772879
+ cigbacc = 0.32875
+ acnqsmod = 0
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ lvoff = -1.4258682e-8
+ toxref = 3e-9
+ tnoimod = 0
+ pags = 2.8299487e-13
+ rbodymod = 0
+ lvsat = -0.0002
+ lvth0 = 5.0775324e-8
+ ntox = 1.0
+ pcit = -1.966418e-16
+ pclm = 1.4152454
+ cigbinv = 0.006
+ delta = 0.007595625
+ laigc = -1.4938914e-10
+ tvfbsdoff = 0.022
+ rnoia = 0
+ rnoib = 0
+ phin = 0.15
+ pkt1 = 4.9928912e-14
+ pkt2 = 1.3351872e-15
+ pketa = -3.7835355e-14
+ version = 4.5
+ ngate = 8e+20
+ ltvoff = -2.0733557e-10
+ ngcon = 1
+ tempmod = 0
+ wpclm = -1.3730014e-7
+ wpdiblc2 = -4.8108443e-11
+ gbmin = 1e-12
+ rbdb = 50
+ pua1 = 6.0905252e-22
+ prwb = 0
+ prwg = 0
+ pub1 = -5.9770157999999995e-31
+ jswgd = 1.28e-13
+ puc1 = 1.7562426e-23
+ jswgs = 1.28e-13
+ rbpb = 50
+ rbpd = 50
+ aigbacc = 0.02
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ pute = 3.9602525e-13
+ lku0we = 2.5e-11
+ rdsw = 100
+ wvfbsdoff = 0
+ epsrox = 3.9
+ lvfbsdoff = 0
+ rdsmod = 0
+ aigbinv = 0.0163
+ igbmod = 1
+ wkvth0we = 2e-12
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ pbswgd = 0.95
+ pbswgs = 0.95
+ rshg = 15.6
+ trnqsmod = 0
+ tvoff = 0.0020267011
+ igcmod = 1
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ poxedge = 1
+ ku0we = -0.0007
+ beta0 = 13
+ tnom = 25
+ rgatemod = 0
+ leta0 = 1.6000000000000003e-9
+ binunit = 2
+ tnjtsswg = 1
+ toxe = 2.43e-9
+ paigsd = -9.9503825e-23
+ toxm = 2.43e-9
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ permod = 1
+ wags = -1.2353313e-7
+ wcit = 5.224659099999999e-10
+ dmcgt = 0
+ tcjsw = 0.000357
+ voff = -0.11150014
+ acde = 0.4
+ voffcv = -0.16942
+ wpemod = 1
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ vsat = 103058.98
+ wint = 0
+ vth0 = 0.31744708
+ wkt1 = -5.3747252999999996e-8
+ wkt2 = -3.7226997e-9
+ wmax = 8.9974e-6
+ aigc = 0.011783086
+ bigsd = 0.00125
+ wmin = 8.974e-7
+ wvoff = 2.6904676e-9
+ wua1 = -8.0608962e-16
+ wub1 = 8.0443355e-25
+ wuc1 = -2.8097884e-18
+ wvsat = -0.0017920539
+ wvth0 = -1.4728173e-8
+ bigc = 0.001442
+ wute = -4.4497219e-7
+ wwlc = 0
+ waigc = 2.7413515e-11
+ tpbswg = 0.0009
+ njtsswg = 9
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ lketa = 3.2718606e-9
+ xtsswgd = 0.18
+ cgsl = 3.31989e-12
+ ijthsfwd = 0.01
+ cgso = 4.90562e-11
+ xtsswgs = 0.18
+ cigc = 0.000625
+ xpart = 1
+ ckappad = 0.6
+ ckappas = 0.6
+ ptvoff = 5.4992103e-16
+ pdiblc1 = 0
+ pdiblc2 = 0.018625664
+ pdiblcb = -0.3
+ waigsd = 3.0716862e-12
+ egidl = 0.29734
+ diomod = 1
+ ijthsrev = 0.01
+ pditsd = 0
+ pditsl = 0
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ cjswgd = 2.66208e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.66208e-10
+ ags = 0.80387747
+ bigbacc = 0.002588
+ cjd = 0.001281008
+ cit = -7.7402473e-5
+ cjs = 0.001281008
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 9.8024918e-9
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ k2we = 5e-5
+ kvth0we = 0.00018
+ dsub = 0.75
+ dtox = 2.7e-10
+ mjswgd = 0.85
+ mjswgs = 0.85
+ pvfbsdoff = 0
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ la0 = -2.0592205e-6
+ lintnoi = -1.5e-8
+ ppdiblc2 = 2.7806803e-16
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = 0.09432272500000001
+ tcjswg = 0.001
+ kt1 = -0.19009298
+ lk2 = -1.3154073e-8
+ kt2 = -0.051410181
+ bigbinv = 0.004953
+ llc = 0
+ vtsswgd = 4.2
+ lln = 1
+ vtsswgs = 4.2
+ lu0 = -1.9868409e-9
+ mjd = 0.26
+ lua = -2.2049077e-16
+ mjs = 0.26
+ lub = -1.5408759e-27
+ luc = 1.1211784e-18
+ lud = 0
+ pvoff = -2.8116001e-15
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 3.0846188e-13
+ eta0 = 0.3
+ nsd = 1e+20
+ pbd = 0.52
+ pat = -8.3091187e-9
+ pbs = 0.52
+ pk2 = -1.9754424e-15
+ cdscb = 0
+ cdscd = 0
+ etab = -0.24888148
+ pu0 = 1.1790383100000001e-17
+ pvsat = -2.24e-11
+ prt = 0
+ pua = 2.7693259e-23
+ pub = -6.3482817e-32
+ puc = -1.7214163e-23
+ pud = 0
+ wk2we = 5e-12
+ pvth0 = 3.3203639e-15
+ drout = 0.56
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 1.3608919e-9
+ ub1 = -8.3548641e-19
+ uc1 = 2.6015633e-11
+ paigc = -9.5524673e-18
+ tpb = 0.0014
+ wa0 = -2.8614611e-7
+ ute = -0.95836072
+ wat = 0.00092088084
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -3.5722648e-9
+ voffl = 0
+ wlc = 0
+ wln = 1
+ wu0 = -2.9901465e-10
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -4.3846243e-17
+ wub = 4.7661234e-26
+ wuc = -5.9424224e-18
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ a0 = 3.5070197
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ weta0 = 0
+ pkvth0we = -1.3e-19
+ at = 61490.242
+ cf = 8.15e-11
+ wetab = -1.0073378e-8
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.024885497
+ k3 = -1.8419
+ em = 1000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.015641155
+ fprout = 300
+ w0 = 0
+ ua = -1.7947198e-9
+ ub = 2.0993593e-18
+ uc = 7.4047731e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ )

.model nch_fs_11 nmos (
+ level = 54
+ ku0we = -0.0007
+ beta0 = 13
+ wku0we = 2e-11
+ leta0 = 1.6000000000000003e-9
+ rbdb = 50
+ mobmod = 0
+ pua1 = 9.7840116e-23
+ prwb = 0
+ prwg = 0
+ pub1 = -1.2272721e-31
+ puc1 = -3.5940917e-24
+ a0 = 1.2386098
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ wtvfbsdoff = 0
+ at = 220073.87
+ cf = 8.15e-11
+ rbpb = 50
+ rbpd = 50
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.024132723
+ k3 = -1.8419
+ rbps = 50
+ em = 1000000.0
+ rbsb = 50
+ pvag = 1.2
+ ll = 0
+ lw = 0
+ u0 = 0.015141687999999999
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ w0 = 0
+ ua = -1.9419497e-9
+ ub = 2.1613601e-18
+ uc = 9.7509556e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ rdsw = 100
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ ijthsfwd = 0.01
+ ltvfbsdoff = 0
+ dmcgt = 0
+ tcjsw = 0.000357
+ laigsd = -9.7335958e-18
+ ijthsrev = 0.01
+ rshg = 15.6
+ njtsswg = 9
+ bigsd = 0.00125
+ ptvfbsdoff = 0
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ wvoff = -7.7864574e-9
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.014827337
+ pdiblcb = -0.3
+ wvsat = -0.0017920539
+ ppdiblc2 = 2.4623293e-15
+ tnom = 25
+ wvth0 = -4.4261894e-9
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ waigc = -9.5733062e-12
+ lketa = -3.0044615e-8
+ bigbacc = 0.002588
+ xpart = 1
+ wags = 1.2380313e-6
+ kvth0we = 0.00018
+ toxref = 3e-9
+ egidl = 0.29734
+ pkvth0we = -1.3e-19
+ wcit = 1.9976376999999998e-10
+ ags = 0.15741391999999998
+ cjd = 0.001281008
+ cit = 0.0013334381
+ voff = -0.11121991
+ lintnoi = -1.5e-8
+ cjs = 0.001281008
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ acde = 0.4
+ dlc = 9.8024918e-9
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ k3b = 1.9326
+ vtsswgs = 4.2
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ vsat = 103058.98
+ wint = 0
+ vfbsdoff = 0.02
+ vth0 = 0.36599507
+ wkt1 = 1.5268642999999998e-8
+ wkt2 = -3.7425887e-9
+ wmax = 8.9974e-6
+ la0 = -4.0335612e-8
+ aigc = 0.011680759
+ wmin = 8.974e-7
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.0468167
+ kt1 = -0.22273968
+ lk2 = -1.2484105e-8
+ kt2 = -0.052902736
+ llc = 0
+ lln = 1
+ lu0 = -1.5423156e-9
+ mjd = 0.26
+ ltvoff = -6.7137092e-10
+ lua = -8.9456155e-17
+ mjs = 0.26
+ lub = -5.6721601e-26
+ luc = -1.9759846e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = -3.420874e-13
+ nsd = 1e+20
+ pbd = 0.52
+ pat = -3.6770881e-9
+ pbs = 0.52
+ pk2 = 6.3553328e-16
+ pvfbsdoff = 0
+ paramchk = 1
+ pu0 = 2.8138232e-17
+ wua1 = -2.3169366e-16
+ wub1 = 2.7075449e-25
+ prt = 0
+ wuc1 = 2.096158e-17
+ pua = -3.3732216e-24
+ pub = 1.7089792e-32
+ puc = 7.8894695e-24
+ pud = 0
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 9.9427719e-10
+ bigc = 0.001442
+ ub1 = -5.7879508e-19
+ uc1 = 6.536871e-11
+ pvoff = 6.5128631e-15
+ tpb = 0.0014
+ wwlc = 0
+ wa0 = 4.4480813e-7
+ ute = -1
+ wat = -0.0042836479
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -6.5059453e-9
+ cdscb = 0
+ cdscd = 0
+ lku0we = 2.5e-11
+ wlc = 0
+ wln = 1
+ wu0 = -3.1738302e-10
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -8.9400845e-18
+ wub = -4.2869787e-26
+ pvsat = -2.24e-11
+ wuc = -3.4148751e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ epsrox = 3.9
+ cdsc = 0
+ wk2we = 5e-12
+ pvth0 = -5.8484018000000006e-15
+ drout = 0.56
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ ijthdfwd = 0.01
+ cgsl = 3.31989e-12
+ paigc = 2.3365803e-17
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ rdsmod = 0
+ nfactor = 1
+ voffl = 0
+ igbmod = 1
+ weta0 = 0
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ wetab = -1.0073378e-8
+ pbswgd = 0.95
+ pbswgs = 0.95
+ ijthdrev = 0.01
+ igcmod = 1
+ cgidl = 0.22
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ lpdiblc2 = 2.7646188e-9
+ nigbacc = 10
+ k2we = 5e-5
+ pbswd = 0.8
+ pbsws = 0.8
+ dsub = 0.75
+ dtox = 2.7e-10
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ nigbinv = 10
+ paigsd = 8.7660773e-23
+ eta0 = 0.3
+ pdits = 0
+ etab = -0.24888148
+ cigsd = 0.069865
+ lkvth0we = -2e-12
+ permod = 1
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ pk2we = -1e-19
+ fnoimod = 1
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ acnqsmod = 0
+ eigbinv = 1.1
+ voffcv = -0.16942
+ wpemod = 1
+ tnoia = 0
+ rbodymod = 0
+ peta0 = 0.0
+ wketa = -4.0591301e-8
+ tpbsw = 0.0019
+ cjswd = 7.7408e-11
+ cjsws = 7.7408e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ cigbacc = 0.32875
+ wpdiblc2 = -2.5023346e-9
+ tnoimod = 0
+ tpbswg = 0.0009
+ cigbinv = 0.006
+ scref = 1e-6
+ ptvoff = 2.4706364e-16
+ pigcd = 2.621
+ keta = -0.026640801
+ aigsd = 0.010772879
+ waigsd = 3.0714759e-12
+ version = 4.5
+ lvoff = -1.4508081e-8
+ lags = 5.1202402e-7
+ wkvth0we = 2e-12
+ tempmod = 0
+ jswd = 1.28e-13
+ diomod = 1
+ jsws = 1.28e-13
+ lcit = -1.2990653e-10
+ lvsat = -0.0002
+ kt1l = 0
+ lvth0 = 7.5676154e-9
+ pditsd = 0
+ pditsl = 0
+ trnqsmod = 0
+ cjswgd = 2.66208e-10
+ tvfbsdoff = 0.022
+ pku0we = -1.5e-18
+ cjswgs = 2.66208e-10
+ delta = 0.007595625
+ laigc = -5.8318716e-11
+ aigbacc = 0.02
+ lint = 6.5375218e-9
+ rnoia = 0
+ rnoib = 0
+ lkt1 = -1.6961753e-8
+ lkt2 = -1.1643768e-8
+ lmax = 8.9908e-7
+ lmin = 4.4908e-7
+ pketa = 3.1782283e-14
+ mjswgd = 0.85
+ lpe0 = 9.2e-8
+ ngate = 8e+20
+ mjswgs = 0.85
+ lpeb = 2.5e-7
+ ngcon = 1
+ wpclm = -1.3730014e-7
+ aigbinv = 0.0163
+ tcjswg = 0.001
+ minv = -0.3
+ rgatemod = 0
+ lua1 = -1.1368255e-16
+ lub1 = 2.9744732e-26
+ luc1 = 4.1671397e-18
+ gbmin = 1e-12
+ tnjtsswg = 1
+ ndep = 1e+18
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ lwlc = 0
+ moin = 5.1
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ nigc = 3.083
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ poxedge = 1
+ fprout = 300
+ xrcrg1 = 12
+ xrcrg2 = 1
+ pags = -9.2879744e-13
+ ntox = 1.0
+ pcit = 9.056310000000001e-17
+ binunit = 2
+ pclm = 1.4152454
+ tvoff = 0.0025480892
+ wtvoff = -5.5551488e-10
+ xjbvd = 1
+ phin = 0.15
+ xjbvs = 1
+ lk2we = -1.5e-12
+ pkt1 = -1.1495235000000001e-14
+ pkt2 = 1.3528884e-15
+ capmod = 2
+ )

.model nch_fs_12 nmos (
+ level = 54
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ ptvfbsdoff = 0
+ cigbacc = 0.32875
+ laigsd = -9.015225e-17
+ wkvth0we = 2e-12
+ tnoia = 0
+ tnoimod = 0
+ trnqsmod = 0
+ peta0 = 0.0
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ wketa = 1.7936379e-8
+ tpbsw = 0.0019
+ a0 = 1.7327189
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ cigbinv = 0.006
+ at = 153009.14
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.017641707
+ k3 = -1.8419
+ em = 1000000.0
+ cjswd = 7.7408e-11
+ ll = -1.18e-13
+ cjsws = 7.7408e-11
+ lw = 0
+ u0 = 0.013035620999999999
+ w0 = 0
+ mjswd = 0.11
+ ua = -2.1226101e-9
+ ub = 2.1428106e-18
+ uc = 6.8443458e-11
+ ud = 0
+ mjsws = 0.11
+ agidl = 9.41e-8
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ k2we = 5e-5
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ dsub = 0.75
+ dtox = 2.7e-10
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ version = 4.5
+ rgatemod = 0
+ tnjtsswg = 1
+ tempmod = 0
+ eta0 = 0.3
+ etab = -0.24888148
+ aigbacc = 0.02
+ scref = 1e-6
+ pigcd = 2.621
+ aigsd = 0.010772879
+ toxref = 3e-9
+ lvoff = -6.1071145e-9
+ aigbinv = 0.0163
+ lvsat = -0.0002
+ lvth0 = -5.421492e-9
+ tvfbsdoff = 0.022
+ delta = 0.007595625
+ laigc = -1.9233809e-11
+ rnoia = 0
+ rnoib = 0
+ ltvoff = -1.0250882e-10
+ pketa = 6.0301037e-15
+ ngate = 8e+20
+ ngcon = 1
+ wpclm = -2.8227848e-7
+ poxedge = 1
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ lku0we = 2.5e-11
+ wvfbsdoff = 0
+ epsrox = 3.9
+ lvfbsdoff = 0
+ binunit = 2
+ rdsmod = 0
+ ijthsfwd = 0.01
+ igbmod = 1
+ keta = -0.041938217
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ lags = 4.5664516e-7
+ pbswgd = 0.95
+ pbswgs = 0.95
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 1.6114929e-10
+ ijthsrev = 0.01
+ igcmod = 1
+ kt1l = 0
+ tvoff = 0.0012552207
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ lint = 9.7879675e-9
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ lkt1 = -1.00758544e-8
+ lkt2 = -3.7159363e-9
+ lmax = 4.4908e-7
+ lmin = 2.1577e-7
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ ku0we = -0.0007
+ paigsd = 8.167794e-23
+ ppdiblc2 = -2.773275e-15
+ beta0 = 13
+ minv = -0.3
+ lua1 = -3.2594611e-17
+ lub1 = -2.980043e-26
+ leta0 = 1.6000000000000003e-9
+ luc1 = -3.5163101e-18
+ ndep = 1e+18
+ ppclm = 6.379047e-14
+ lwlc = 0
+ permod = 1
+ moin = 5.1
+ dlcig = 2.5e-9
+ nigc = 3.083
+ bgidl = 2320000000.0
+ njtsswg = 9
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ pkvth0we = -1.3e-19
+ dmcgt = 0
+ voffcv = -0.16942
+ ckappad = 0.6
+ wpemod = 1
+ ckappas = 0.6
+ tcjsw = 0.000357
+ pdiblc1 = 0
+ pdiblc2 = 0.026288388
+ pags = 8.4375107e-13
+ pdiblcb = -0.3
+ ntox = 1.0
+ pcit = -7.489201199999999e-17
+ pclm = 1.5752657
+ vfbsdoff = 0.02
+ phin = 0.15
+ bigsd = 0.00125
+ pkt1 = -4.2148923e-16
+ pkt2 = -1.2933793e-15
+ bigbacc = 0.002588
+ wvoff = 1.1733398e-8
+ paramchk = 1
+ wvsat = -0.0017920539
+ kvth0we = 0.00018
+ wvth0 = -2.2574896000000002e-8
+ tpbswg = 0.0009
+ rbdb = 50
+ pua1 = 1.9082335e-23
+ prwb = 0
+ prwg = 0
+ pub1 = -2.3478905e-32
+ puc1 = -7.9472634e-24
+ waigc = 5.7897385e-11
+ lintnoi = -1.5e-8
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ rdsw = 100
+ ags = 0.28327496999999996
+ lketa = -2.3313752e-8
+ ijthdfwd = 0.01
+ ptvoff = -1.6297696e-16
+ xpart = 1
+ cjd = 0.001281008
+ cit = 0.00067194759
+ cjs = 0.001281008
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ waigsd = 3.0714895e-12
+ dlc = 1.30529375e-8
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ egidl = 0.29734
+ diomod = 1
+ la0 = -2.5774361e-7
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.017308219
+ pditsd = 0
+ pditsl = 0
+ kt1 = -0.23838945
+ ijthdrev = 0.01
+ lk2 = -9.6280577e-9
+ kt2 = -0.070920535
+ cjswgd = 2.66208e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.66208e-10
+ llc = -1.18e-13
+ lln = 0.7
+ rshg = 15.6
+ lu0 = -6.1564579e-10
+ mjd = 0.26
+ lua = -9.9655811e-18
+ mjs = 0.26
+ lub = -4.8559819e-26
+ luc = -6.9707629e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 9.4027643e-14
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 2.5179517e-9
+ lpdiblc2 = -2.2782436e-9
+ pbs = 0.52
+ pk2 = 9.5548939e-17
+ pu0 = 1.0007793799999999e-17
+ prt = 0
+ pua = -7.1355685e-24
+ pub = 6.4921301e-33
+ puc = 2.8995668e-24
+ pud = 0
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 8.0998641e-10
+ ub1 = -4.4346517e-19
+ uc1 = 8.2831095e-11
+ mjswgd = 0.85
+ mjswgs = 0.85
+ tpb = 0.0014
+ wa0 = -5.4636242e-7
+ nfactor = 1
+ pvfbsdoff = 0
+ ute = -1
+ wat = -0.018363284
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -5.2787082e-9
+ tcjswg = 0.001
+ wlc = 0
+ wln = 1
+ wu0 = -2.7617748e-10
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -3.8929611e-19
+ wub = -1.8784192e-26
+ wuc = -2.2808063e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ tnom = 25
+ pvoff = -2.0758734e-15
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ cdscb = 0
+ cdscd = 0
+ lkvth0we = -2e-12
+ pvsat = -2.24e-11
+ wk2we = 5e-12
+ pvth0 = 2.1370293e-15
+ drout = 0.56
+ paigc = -6.3213007e-18
+ nigbacc = 10
+ voffl = 0
+ acnqsmod = 0
+ wags = -2.7904881000000002e-6
+ fprout = 300
+ weta0 = 0
+ wetab = -1.0073378e-8
+ wcit = 5.7579813e-10
+ xrcrg1 = 12
+ xrcrg2 = 1
+ lpclm = -7.0408907e-8
+ voff = -0.13031302
+ rbodymod = 0
+ nigbinv = 10
+ acde = 0.4
+ cgidl = 0.22
+ vsat = 103058.98
+ wtvoff = 3.7639557e-10
+ wint = 0
+ vth0 = 0.39551577
+ wkt1 = -9.8989616e-9
+ wkt2 = 2.2716562e-9
+ wmax = 8.9974e-6
+ wtvfbsdoff = 0
+ aigc = 0.01159193
+ wmin = 8.974e-7
+ capmod = 2
+ pbswd = 0.8
+ pbsws = 0.8
+ ltvfbsdoff = 0
+ fnoimod = 1
+ wua1 = -5.2698704e-17
+ wub1 = 4.5190152e-26
+ wku0we = 2e-11
+ wuc1 = 3.0855152e-17
+ eigbinv = 1.1
+ wpdiblc2 = 9.3967661e-9
+ bigc = 0.001442
+ mobmod = 0
+ wwlc = 0
+ pdits = 0
+ cigsd = 0.069865
+ cdsc = 0
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ )

.model nch_fs_13 nmos (
+ level = 54
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ lint = 9.7879675e-9
+ bigsd = 0.00125
+ lkt1 = -4.101126e-9
+ lkt2 = -5.6046527e-10
+ lmax = 2.1577e-7
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ lmin = 9e-8
+ wvoff = -2.233608000000001e-9
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ wvsat = -0.00035982647999999954
+ minv = -0.3
+ wvth0 = -9.062617000000002e-9
+ lua1 = 8.0644671e-18
+ lub1 = -5.5160301e-26
+ luc1 = -4.6427809e-18
+ ags = 2.4474682
+ ndep = 1e+18
+ waigc = 3.6164887e-11
+ cjd = 0.001281008
+ cit = 0.0010410649
+ cjs = 0.001281008
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ lwlc = 0
+ dlc = 1.30529375e-8
+ k3b = 1.9326
+ moin = 5.1
+ lkvth0we = -2e-12
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ nigc = 3.083
+ lketa = -1.0074554e-8
+ xpart = 1
+ la0 = -3.95931149e-8
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.0020360989
+ toxref = 3e-9
+ kt1 = -0.26670569
+ lk2 = -2.2996724e-9
+ kt2 = -0.085875374
+ llc = -1.18e-13
+ lln = 0.7
+ a0 = 0.69883298
+ a1 = 0
+ a2 = 1
+ lu0 = -1.8979706e-10
+ b0 = 0
+ b1 = 0
+ acnqsmod = 0
+ mjd = 0.26
+ lua = 2.3685126e-17
+ mjs = 0.26
+ lub = -3.581049857e-26
+ luc = -1.971816e-18
+ lud = 0
+ at = 80629.42
+ cf = 8.15e-11
+ lwc = 0
+ noff = 2.7195
+ lwl = 0
+ lwn = 1
+ ef = 1.0
+ k1 = 0.274
+ k2 = -0.017089977
+ k3 = -1.8419
+ em = 1000000.0
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ njd = 1.02
+ njs = 1.02
+ nfactor = 1
+ pa0 = 5.1229998e-14
+ egidl = 0.29734
+ ll = -1.18e-13
+ lw = 0
+ u0 = 0.011017379999999998
+ w0 = 0
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 7.9117566e-10
+ pbs = 0.52
+ ua = -2.2820921e-9
+ ub = 2.0823870489000003e-18
+ uc = 4.4751766e-11
+ ud = 0
+ pk2 = 1.6389978e-16
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ pu0 = -2.0701017e-17
+ prt = 0
+ pua = 6.5907354e-24
+ pub = -1.1536808500000001e-32
+ puc = -4.2264406e-24
+ pud = 0
+ pags = -3.4153056e-19
+ rbodymod = 0
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 6.1728936e-10
+ ub1 = -3.2327621e-19
+ uc1 = 8.8169819e-11
+ ntox = 1.0
+ pcit = -7.2109378e-17
+ pclm = 1.3619854
+ tpb = 0.0014
+ wa0 = -3.4353242e-7
+ ute = -1
+ wat = -0.010179511
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -5.6026458e-9
+ wlc = 0
+ wln = 1
+ wu0 = -1.30638093e-10
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -6.5442869e-17
+ wub = 6.6660889e-26
+ wuc = 1.0964484e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ ltvoff = 4.8985213e-12
+ phin = 0.15
+ pvfbsdoff = 0
+ nigbacc = 10
+ pkt1 = 2.8803122e-15
+ pkt2 = -3.7226831e-16
+ wpdiblc2 = -7.3538749e-9
+ lku0we = 2.5e-11
+ pvoff = 8.711494700000001e-16
+ rbdb = 50
+ pua1 = -3.4072796e-24
+ prwb = 0
+ prwg = 0
+ pub1 = 3.4449133e-33
+ epsrox = 3.9
+ puc1 = 3.7978198e-24
+ cdscb = 0
+ cdscd = 0
+ rbpb = 50
+ rbpd = 50
+ nigbinv = 10
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ pvsat = -3.2459949e-10
+ wk2we = 5e-12
+ pvth0 = -7.140435999999998e-16
+ rdsw = 100
+ drout = 0.56
+ rdsmod = 0
+ igbmod = 1
+ paigc = -1.7357437e-18
+ voffl = 0
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ pbswgd = 0.95
+ pbswgs = 0.95
+ weta0 = 0
+ wetab = -1.0073378e-8
+ wkvth0we = 2e-12
+ fnoimod = 1
+ lpclm = -2.540677e-8
+ igcmod = 1
+ eigbinv = 1.1
+ rshg = 15.6
+ trnqsmod = 0
+ cgidl = 0.22
+ pbswd = 0.8
+ pbsws = 0.8
+ paigsd = -5.1229584e-23
+ rgatemod = 0
+ tnom = 25
+ cigbacc = 0.32875
+ tnjtsswg = 1
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ permod = 1
+ pdits = 0
+ cigsd = 0.069865
+ tnoimod = 0
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ cigbinv = 0.006
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ wags = 1.2083338e-6
+ voffcv = -0.16942
+ wpemod = 1
+ wcit = 5.6261028e-10
+ tnoia = 0
+ voff = -0.1572150866
+ version = 4.5
+ acde = 0.4
+ tempmod = 0
+ peta0 = 0.0
+ vsat = 102561.23895
+ wint = 0
+ vth0 = 0.4100123399
+ wketa = 1.0437078e-7
+ wkt1 = -2.554731e-8
+ wkt2 = -2.0937989e-9
+ tpbsw = 0.0019
+ wmax = 8.9974e-6
+ aigc = 0.011522737
+ wmin = 8.974e-7
+ cjswd = 7.7408e-11
+ aigbacc = 0.02
+ cjsws = 7.7408e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ wua1 = 5.3887147e-17
+ wub1 = -8.2410881e-26
+ wuc1 = -2.4808749e-17
+ tpbswg = 0.0009
+ bigc = 0.001442
+ wwlc = 0
+ aigbinv = 0.0163
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ ptvoff = 8.9623963e-17
+ ijthsfwd = 0.01
+ scref = 1e-6
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ waigsd = 3.0721194e-12
+ pigcd = 2.621
+ aigsd = 0.010772879
+ diomod = 1
+ lvoff = -4.3079245999999997e-10
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 2.66208e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.66208e-10
+ lvsat = -9.496033999999993e-5
+ tvfbsdoff = 0.022
+ ijthsrev = 0.01
+ lvth0 = -8.480254980000001e-9
+ poxedge = 1
+ delta = 0.007595625
+ laigc = -4.6341008e-12
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ binunit = 2
+ rnoia = 0
+ rnoib = 0
+ mjswgd = 0.85
+ mjswgs = 0.85
+ k2we = 5e-5
+ pketa = -1.2207451e-14
+ tcjswg = 0.001
+ ngate = 8e+20
+ dsub = 0.75
+ ngcon = 1
+ dtox = 2.7e-10
+ wpclm = -2.3899735e-8
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ ppdiblc2 = 7.6111026e-16
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ eta0 = 0.3
+ etab = -0.24888148
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ fprout = 300
+ wtvfbsdoff = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ pkvth0we = -1.3e-19
+ ltvfbsdoff = 0
+ wtvoff = -8.2076521e-10
+ tvoff = 0.00074618122
+ vfbsdoff = 0.02
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ capmod = 2
+ njtsswg = 9
+ wku0we = 2e-11
+ paramchk = 1
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ ku0we = -0.0007
+ mobmod = 0
+ beta0 = 13
+ leta0 = 1.6000000000000003e-9
+ ckappad = 0.6
+ ptvfbsdoff = 0
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.022446923
+ pdiblcb = -0.3
+ ppclm = 9.2725546e-15
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ ijthdfwd = 0.01
+ keta = -0.10468292
+ bigbacc = 0.002588
+ laigsd = 3.9592657e-17
+ lags = 3.7696529e-13
+ dmcgt = 0
+ tcjsw = 0.000357
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 8.3265533e-11
+ kvth0we = 0.00018
+ ijthdrev = 0.01
+ kt1l = 0
+ lintnoi = -1.5e-8
+ lpdiblc2 = -1.4676946e-9
+ bigbinv = 0.004953
+ )

.model nch_fs_14 nmos (
+ level = 54
+ poxedge = 1
+ binunit = 2
+ scref = 1e-6
+ toxref = 3e-9
+ pigcd = 2.621
+ aigsd = 0.010772879
+ wags = 1.2083302e-6
+ lvoff = -2.0678068800000007e-9
+ pkvth0we = -1.3e-19
+ wcit = 1.9125736e-10
+ tvfbsdoff = 0.022
+ voff = -0.13980004150000003
+ lvsat = 0.00098775289
+ lvth0 = 1.7575669099999996e-9
+ acde = 0.4
+ delta = 0.007595625
+ vsat = 91042.9961
+ laigc = -2.2637509e-11
+ wint = 0
+ vfbsdoff = 0.02
+ vth0 = 0.3010993353
+ ltvoff = 1.2509019e-10
+ wkt1 = 8.1270806e-8
+ wkt2 = 1.6147625e-8
+ rnoia = 0
+ rnoib = 0
+ wmax = 8.9974e-6
+ aigc = 0.011714263
+ wmin = 8.974e-7
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ pketa = 8.4378567e-15
+ ngate = 8e+20
+ paramchk = 1
+ ngcon = 1
+ wpclm = 3.4675908e-7
+ wua1 = -1.154179e-16
+ wub1 = 3.1505286e-27
+ wuc1 = 9.7519251e-17
+ lku0we = 2.5e-11
+ a0 = -0.035582299999999956
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ bigc = 0.001442
+ gbmin = 1e-12
+ epsrox = 3.9
+ at = 65883.509
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = -0.036187969
+ k3 = -1.8419
+ wvfbsdoff = 0
+ em = 1000000.0
+ wwlc = 0
+ jswgd = 1.28e-13
+ lvfbsdoff = 0
+ jswgs = 1.28e-13
+ ll = 0
+ lw = 0
+ u0 = 0.0075965756
+ w0 = 0
+ ua = -2.421907e-9
+ ub = 1.9130826320999997e-18
+ uc = 4.338735e-12
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ rdsmod = 0
+ cdsc = 0
+ igbmod = 1
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ ijthdfwd = 0.01
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ pbswgd = 0.95
+ pbswgs = 0.95
+ njtsswg = 9
+ igcmod = 1
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ ijthdrev = 0.01
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.006833075
+ pdiblcb = -0.3
+ tvoff = -0.00053245355
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ lpdiblc2 = 7.1362462e-15
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ k2we = 5e-5
+ paigsd = 1.5255572e-23
+ dsub = 0.75
+ dtox = 2.7e-10
+ ku0we = -0.0007
+ bigbacc = 0.002588
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ beta0 = 13
+ leta0 = 4.2128654e-9
+ letab = -2.2297043e-8
+ permod = 1
+ kvth0we = 0.00018
+ ppclm = -2.5569374e-14
+ eta0 = 0.27220356
+ etab = -0.011678893
+ lkvth0we = -2e-12
+ dlcig = 2.5e-9
+ lintnoi = -1.5e-8
+ bgidl = 2320000000.0
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ acnqsmod = 0
+ voffcv = -0.16942
+ wpemod = 1
+ dmcgt = 0
+ tcjsw = 0.000357
+ rbodymod = 0
+ bigsd = 0.00125
+ ags = 2.4474722
+ wvoff = 8.241506600000007e-9
+ cjd = 0.001281008
+ cit = 0.00030181593
+ cjs = 0.001281008
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 3.26497e-9
+ tpbswg = 0.0009
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ wvsat = -0.010835494899999996
+ nfactor = 1
+ wvth0 = -1.65057091e-8
+ wpdiblc2 = 7.4309162e-10
+ waigc = -2.4473999e-12
+ la0 = 2.94419216e-8
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.00064998333
+ kt1 = -0.41803712
+ lk2 = -5.0446112e-10
+ kt2 = -0.10268076
+ llc = 0
+ lln = 1
+ lu0 = 1.3175857e-10
+ mjd = 0.26
+ lua = 3.6827721e-17
+ mjs = 0.26
+ lub = -1.9895881809999996e-26
+ luc = 1.827009e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ ptvoff = -1.5034232e-16
+ njd = 1.02
+ njs = 1.02
+ pa0 = 7.627786000000002e-15
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 9.5747885e-10
+ pbs = 0.52
+ pk2 = 1.6131306e-16
+ waigsd = 3.0714121e-12
+ lketa = 2.8547804e-8
+ pu0 = -1.7222607e-16
+ prt = 0
+ pua = -1.4490045e-23
+ xpart = 1
+ pub = 2.3973370000000036e-34
+ puc = 4.0045874e-24
+ pud = 0
+ rsh = 17.5
+ keta = -0.51555907
+ tcj = 0.00076
+ ua1 = 9.0255397e-10
+ ub1 = -8.0270486e-19
+ uc1 = -7.4218809e-11
+ diomod = 1
+ tpb = 0.0014
+ nigbacc = 10
+ wa0 = 1.203209e-7
+ egidl = 0.29734
+ ute = -1
+ wat = -0.011948694
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -5.5751276e-9
+ pditsd = 0
+ pditsl = 0
+ wlc = 0
+ wln = 1
+ wkvth0we = 2e-12
+ wu0 = 1.4813304999999998e-9
+ cjswgd = 2.66208e-10
+ pku0we = -1.5e-18
+ xgl = -1.09e-8
+ cjswgs = 2.66208e-10
+ xgw = 0
+ wua = 1.5882075e-16
+ wub = -5.862147e-26
+ wuc = -7.6599643e-17
+ wud = 0
+ wwc = 0
+ jswd = 1.28e-13
+ wwl = 0
+ wwn = 1
+ jsws = 1.28e-13
+ lcit = 1.5275494e-10
+ kt1l = 0
+ trnqsmod = 0
+ nigbinv = 10
+ lint = 0
+ mjswgd = 0.85
+ mjswgs = 0.85
+ lkt1 = 1.0124028e-8
+ lkt2 = 1.0192413e-9
+ pvfbsdoff = 0
+ lmax = 9e-8
+ tcjswg = 0.001
+ lmin = 5.4e-8
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ minv = -0.3
+ rgatemod = 0
+ lua1 = -1.8750406e-17
+ wtvfbsdoff = 0
+ lub1 = -1.00940068e-26
+ luc1 = 1.062175e-17
+ pvoff = -1.135113399999999e-16
+ tnjtsswg = 1
+ fnoimod = 1
+ ndep = 1e+18
+ eigbinv = 1.1
+ cdscb = 0
+ cdscd = 0
+ lwlc = 0
+ moin = 5.1
+ pvsat = 6.601120199999996e-10
+ wk2we = 5e-12
+ pvth0 = -1.439292199999993e-17
+ ltvfbsdoff = 0
+ drout = 0.56
+ nigc = 3.083
+ paigc = 1.8938113e-18
+ fprout = 300
+ voffl = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ weta0 = -3.9858587e-8
+ wetab = 2.7041872e-8
+ lpclm = -8.5343289e-9
+ wtvoff = 1.7320676e-9
+ cigbacc = 0.32875
+ ntox = 1.0
+ pcit = -3.7202203e-17
+ pclm = 1.1824913
+ cgidl = 0.22
+ ptvfbsdoff = 0
+ tnoimod = 0
+ phin = 0.15
+ capmod = 2
+ pkt1 = -7.1605907e-15
+ pkt2 = -2.0869621e-15
+ wku0we = 2e-11
+ cigbinv = 0.006
+ pbswd = 0.8
+ pbsws = 0.8
+ mobmod = 0
+ rbdb = 50
+ pua1 = 1.2507395e-23
+ prwb = 0
+ prwg = 0
+ pub1 = -4.5978592e-33
+ puc1 = -7.7010123e-24
+ version = 4.5
+ pdits = 0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ cigsd = 0.069865
+ tempmod = 0
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ rdsw = 100
+ ijthsfwd = 0.01
+ aigbacc = 0.02
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ laigsd = -1.6939346e-18
+ tnoia = 0
+ ijthsrev = 0.01
+ rshg = 15.6
+ peta0 = 3.7467072e-15
+ aigbinv = 0.0163
+ petab = -3.4888335e-15
+ wketa = -1.1526014e-7
+ tpbsw = 0.0019
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ cjswd = 7.7408e-11
+ cjsws = 7.7408e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ ppdiblc2 = -4.5980291e-21
+ tnom = 25
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ )

.model nch_fs_15 nmos (
+ level = 54
+ fnoimod = 1
+ ltvoff = -2.8596488e-10
+ eigbinv = 1.1
+ pvfbsdoff = 0
+ lku0we = 2.5e-11
+ epsrox = 3.9
+ pvoff = 8.85540199999999e-16
+ cdscb = 0
+ cdscd = 0
+ rdsmod = 0
+ cigbacc = 0.32875
+ pvsat = -3.1524723e-9
+ igbmod = 1
+ wk2we = 5e-12
+ pvth0 = -8.548169999999997e-16
+ drout = 0.56
+ ijthsfwd = 0.01
+ paigc = 1.0773556e-18
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ tnoimod = 0
+ voffl = 0
+ pbswgd = 0.95
+ pbswgs = 0.95
+ keta = 0.067264197
+ cigbinv = 0.006
+ weta0 = 3.2678994e-7
+ igcmod = 1
+ wetab = -1.4667966e-7
+ lpclm = -8.0899178e-8
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 3.1911574e-10
+ ijthsrev = 0.01
+ kt1l = 0
+ cgidl = 0.22
+ version = 4.5
+ a0 = 5.6809619
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = -88751.793
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = -0.016551152
+ k3 = -1.8419
+ em = 1000000.0
+ ll = 0
+ tempmod = 0
+ lw = 0
+ lint = 0
+ u0 = 0.00011525645999999995
+ w0 = 0
+ ua = -3.0786989e-9
+ ub = 2.197681248e-18
+ uc = -5.08518e-12
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ lkt1 = -1.6453162999999998e-8
+ lkt2 = 1.223943e-9
+ lmax = 5.4e-8
+ lmin = 4.5e-8
+ paigsd = -3.180948e-23
+ pbswd = 0.8
+ lpe0 = 9.2e-8
+ pbsws = 0.8
+ lpeb = 2.5e-7
+ aigbacc = 0.02
+ minv = -0.3
+ permod = 1
+ lua1 = 1.293984e-17
+ lub1 = 3.4709433900000004e-26
+ luc1 = 1.702510023e-17
+ ndep = 1e+18
+ pdits = 0
+ lwlc = 0
+ cigsd = 0.069865
+ moin = 5.1
+ aigbinv = 0.0163
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ nigc = 3.083
+ voffcv = -0.16942
+ wpemod = 1
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ pkvth0we = -1.3e-19
+ tnoia = 0
+ ntox = 1.0
+ pcit = 6.3457403e-17
+ pclm = 2.4301611
+ peta0 = -1.7518907e-14
+ petab = 6.5870154e-15
+ vfbsdoff = 0.02
+ wketa = 1.9475197e-7
+ poxedge = 1
+ tpbsw = 0.0019
+ phin = 0.15
+ cjswd = 7.7408e-11
+ cjsws = 7.7408e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ binunit = 2
+ pkt1 = 1.2992179999999999e-14
+ pkt2 = 7.7933247e-16
+ tpbswg = 0.0009
+ paramchk = 1
+ rbdb = 50
+ pua1 = -3.7208869e-24
+ prwb = 0
+ prwg = 0
+ pub1 = -6.9476579e-32
+ puc1 = -1.1133321e-23
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ ptvoff = 3.472697e-16
+ waigsd = 3.0722235e-12
+ rdsw = 100
+ ijthdfwd = 0.01
+ scref = 1e-6
+ diomod = 1
+ pigcd = 2.621
+ aigsd = 0.010772879
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ pditsd = 0
+ pditsl = 0
+ lvoff = -3.7139500800000003e-9
+ cjswgd = 2.66208e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.66208e-10
+ tvfbsdoff = 0.022
+ lvsat = 0.00233730979
+ ijthdrev = 0.01
+ lvth0 = 1.9729352399999987e-9
+ rshg = 15.6
+ delta = 0.007595625
+ laigc = -2.1310273e-11
+ wtvfbsdoff = 0
+ mjswgd = 0.85
+ mjswgs = 0.85
+ rnoia = 0
+ rnoib = 0
+ tcjswg = 0.001
+ ltvfbsdoff = 0
+ pketa = -9.5428465e-15
+ ngate = 8e+20
+ ngcon = 1
+ wpclm = -1.3405624e-6
+ njtsswg = 9
+ tnom = 25
+ wvfbsdoff = 0
+ gbmin = 1e-12
+ lvfbsdoff = 0
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ jswgd = 1.28e-13
+ toxe = 2.43e-9
+ jswgs = 1.28e-13
+ toxm = 2.43e-9
+ ckappad = 0.6
+ lkvth0we = -2e-12
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.0068331981
+ pdiblcb = -0.3
+ fprout = 300
+ ptvfbsdoff = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ acnqsmod = 0
+ wags = 1.2083302e-6
+ wcit = -1.5442530999999999e-9
+ wtvoff = -6.84745e-9
+ bigbacc = 0.002588
+ rbodymod = 0
+ voff = -0.111418263
+ acde = 0.4
+ vsat = 67774.80940000001
+ tvoff = 0.0065547027
+ kvth0we = 0.00018
+ wint = 0
+ vth0 = 0.297386088
+ wkt1 = -2.6619076e-7
+ wkt2 = -3.3271248e-8
+ xjbvd = 1
+ xjbvs = 1
+ wmax = 8.9974e-6
+ lk2we = -1.5e-12
+ capmod = 2
+ aigc = 0.011691379
+ wmin = 8.974e-7
+ lintnoi = -1.5e-8
+ bigbinv = 0.004953
+ wku0we = 2e-11
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ mobmod = 0
+ ku0we = -0.0007
+ wua1 = 1.6438006e-16
+ wub1 = 1.12174916e-24
+ wuc1 = 1.56696984e-16
+ beta0 = 13
+ wpdiblc2 = 7.4301235e-10
+ leta0 = 1.7011061900000003e-9
+ letab = 3.9727723e-8
+ bigc = 0.001442
+ wwlc = 0
+ ppclm = 7.229527e-14
+ cdsc = 0
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ laigsd = 3.532034e-18
+ dmcgt = 0
+ wkvth0we = 2e-12
+ tcjsw = 0.000357
+ nfactor = 1
+ ags = 2.4474722
+ trnqsmod = 0
+ cjd = 0.001281008
+ cit = -0.0025664738
+ cjs = 0.001281008
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ dlc = 3.26497e-9
+ k3b = 1.9326
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ bigsd = 0.00125
+ k2we = 5e-5
+ wvoff = -8.983524000000003e-9
+ la0 = -3.0211764e-7
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = 0.0083188642
+ dsub = 0.75
+ kt1 = 0.040190302
+ lk2 = -1.6433965e-9
+ kt2 = -0.1062101
+ dtox = 2.7e-10
+ llc = 0
+ lln = 1
+ lu0 = 5.656750800000001e-10
+ mjd = 0.26
+ nigbacc = 10
+ lua = 7.492165e-17
+ mjs = 0.26
+ lub = -3.6402602300000003e-26
+ luc = 2.373596e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ wvsat = 0.054898772
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ njd = 1.02
+ njs = 1.02
+ pa0 = -1.230232e-13
+ rgatemod = 0
+ wvth0 = -2.015631999999998e-9
+ nsd = 1e+20
+ pbd = 0.52
+ pat = -8.1375789e-9
+ pbs = 0.52
+ pk2 = 5.8185614e-16
+ tnjtsswg = 1
+ pu0 = -8.0546575e-17
+ prt = 0
+ pua = 3.4306982e-23
+ pub = -6.0757564e-32
+ puc = -7.1571349e-24
+ pud = 0
+ waigc = 1.1629424e-11
+ eta0 = 0.31550975
+ rsh = 17.5
+ etab = -1.0810714
+ tcj = 0.00076
+ ua1 = 3.5617042e-10
+ ub1 = -1.575178019e-18
+ uc1 = -1.8462139999999999e-10
+ tpb = 0.0014
+ wa0 = 2.372924e-6
+ ute = -1
+ wat = 0.14486265
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -1.282587e-8
+ nigbinv = 10
+ lketa = -5.2559457e-9
+ toxref = 3e-9
+ wlc = 0
+ wln = 1
+ wu0 = -9.935035400000001e-11
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -6.825073e-16
+ wub = 9.9305604e-25
+ wuc = 1.1584384e-16
+ wud = 0
+ wwc = 0
+ xpart = 1
+ wwl = 0
+ wwn = 1
+ egidl = 0.29734
+ )

.model nch_fs_16 nmos (
+ level = 54
+ pketa = 8.7750313e-15
+ pkt1 = -8.788479599999999e-16
+ pkt2 = 1.5926682e-15
+ ngate = 8e+20
+ lku0we = 2.5e-11
+ ngcon = 1
+ wpclm = -1.03603352e-6
+ epsrox = 3.9
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ wpdiblc2 = 7.4301235e-10
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ rdsmod = 0
+ bigbacc = 0.002588
+ rbdb = 50
+ pua1 = -1.9060214e-23
+ prwb = 0
+ prwg = 0
+ pub1 = 4.8168331000000005e-32
+ puc1 = 1.47310838e-23
+ igbmod = 1
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ rdsw = 100
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ kvth0we = 0.00018
+ pbswgd = 0.95
+ pbswgs = 0.95
+ lintnoi = -1.5e-8
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ igcmod = 1
+ wkvth0we = 2e-12
+ rshg = 15.6
+ trnqsmod = 0
+ tvoff = 0.002919136
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ paigsd = 4.3875156e-23
+ ku0we = -0.0007
+ permod = 1
+ beta0 = 13
+ rgatemod = 0
+ leta0 = 1.7343207e-8
+ tnom = 25
+ letab = 3.0329695e-8
+ tnjtsswg = 1
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ nfactor = 1
+ ppclm = 5.7373356e-14
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ voffcv = -0.16942
+ wpemod = 1
+ a0 = 3.2177147
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 125884.31
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.023415951
+ k3 = -1.8419
+ em = 1000000.0
+ ll = 0
+ lw = 0
+ ags = 2.4474722
+ u0 = 0.0032670623
+ w0 = 0
+ ua = -2.19661343e-9
+ ub = 1.4860819409999996e-18
+ uc = 2.2595638e-10
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ wags = 1.2083302e-6
+ xl = 4e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ cjd = 0.001281008
+ cit = -0.0057789249
+ cjs = 0.001281008
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dmcgt = 0
+ dlc = 3.26497e-9
+ wcit = 5.1712463999999996e-9
+ tcjsw = 0.000357
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ nigbacc = 10
+ voff = -0.04075972859999999
+ acde = 0.4
+ la0 = -1.8141853e-7
+ vsat = 81047.60070000001
+ wint = 0
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.0021983049
+ vth0 = 0.35253306059999995
+ kt1 = -0.20813859
+ lk2 = -3.6017846e-9
+ kt2 = -0.11042259
+ llc = 0
+ lln = 1
+ lu0 = 4.1123683e-10
+ wkt1 = 1.6891446e-8
+ wkt2 = -4.9869936e-8
+ mjd = 0.26
+ bigsd = 0.00125
+ lua = 3.1699464000000005e-17
+ mjs = 0.26
+ lub = -1.5342368999999952e-27
+ luc = -8.94744e-18
+ lud = 0
+ wmax = 8.9974e-6
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ aigc = 0.011397597
+ wmin = 8.974e-7
+ njs = 1.02
+ pa0 = -1.9996651e-13
+ nsd = 1e+20
+ nigbinv = 10
+ pbd = 0.52
+ pat = 1.2861010000000001e-10
+ pbs = 0.52
+ pk2 = 3.3250012e-16
+ tpbswg = 0.0009
+ pu0 = -6.496246999999995e-18
+ prt = 0
+ pua = 2.7971342e-23
+ pub = -4.5926045000000006e-32
+ puc = -7.6781524e-24
+ pud = 0
+ wvoff = 8.333983999999995e-9
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 4.3071269e-10
+ ub1 = -2.19332361e-19
+ uc1 = 5.294111900000001e-10
+ wua1 = 4.7742754e-16
+ tpb = 0.0014
+ wub1 = -1.27916739e-24
+ wuc1 = -3.71148e-16
+ wvsat = 0.039935568
+ wa0 = 3.9431957e-6
+ wvth0 = -6.398649699999998e-8
+ ute = -1
+ wat = -0.023835087
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -7.7369724e-9
+ bigc = 0.001442
+ wlc = 0
+ wln = 1
+ wu0 = -1.6105853600000001e-9
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -5.5320853e-16
+ wub = 6.903720200000001e-25
+ wuc = 1.2647685e-16
+ wud = 0
+ wwlc = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ waigc = -9.3979847e-11
+ ptvoff = -3.4317401e-17
+ waigsd = 3.0706789e-12
+ fnoimod = 1
+ cdsc = 0
+ eigbinv = 1.1
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ lketa = -2.4929909e-8
+ xtis = 3
+ ijthsfwd = 0.01
+ diomod = 1
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ xpart = 1
+ wtvfbsdoff = 0
+ cigc = 0.000625
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 2.66208e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.66208e-10
+ egidl = 0.29734
+ ltvfbsdoff = 0
+ ijthsrev = 0.01
+ mjswgd = 0.85
+ mjswgs = 0.85
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ cigbacc = 0.32875
+ pvfbsdoff = 0
+ tcjswg = 0.001
+ tnoimod = 0
+ k2we = 5e-5
+ dsub = 0.75
+ dtox = 2.7e-10
+ ptvfbsdoff = 0
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ cigbinv = 0.006
+ pvoff = 3.698261999999959e-17
+ cdscb = 0
+ cdscd = 0
+ eta0 = -0.003716791
+ etab = -0.88927493
+ pvsat = -2.4192770499999994e-9
+ wk2we = 5e-12
+ pvth0 = 2.1817551599999995e-15
+ drout = 0.56
+ version = 4.5
+ fprout = 300
+ paigc = 6.2522098e-18
+ tempmod = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ voffl = 0
+ weta0 = 2.2378028e-8
+ pkvth0we = -1.3e-19
+ wetab = 3.831648e-8
+ aigbacc = 0.02
+ wtvoff = 9.4004181e-10
+ lpclm = -7.043921000000001e-8
+ cgidl = 0.22
+ vfbsdoff = 0.02
+ capmod = 2
+ aigbinv = 0.0163
+ wku0we = 2e-11
+ mobmod = 0
+ pbswd = 0.8
+ pbsws = 0.8
+ paramchk = 1
+ pdits = 0
+ cigsd = 0.069865
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ poxedge = 1
+ ijthdfwd = 0.01
+ laigsd = -2.6649547e-17
+ pk2we = -1e-19
+ keta = 0.46877367
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ binunit = 2
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ tnoia = 0
+ lcit = 4.7652643e-10
+ ijthdrev = 0.01
+ kt1l = 0
+ peta0 = -2.6027237e-15
+ petab = -2.4777955e-15
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ wketa = -1.7908228e-7
+ tpbsw = 0.0019
+ lint = 0
+ cjswd = 7.7408e-11
+ cjsws = 7.7408e-11
+ lkt1 = -4.285047e-9
+ lkt2 = 1.4303548e-9
+ mjswd = 0.11
+ lmax = 4.5e-8
+ mjsws = 0.11
+ agidl = 9.41e-8
+ lmin = 3.6e-8
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ minv = -0.3
+ lua1 = 9.2872684e-18
+ lub1 = -3.17270018e-26
+ luc1 = -1.796249619e-17
+ ndep = 1e+18
+ lwlc = 0
+ lkvth0we = -2e-12
+ moin = 5.1
+ toxref = 3e-9
+ nigc = 3.083
+ scref = 1e-6
+ pigcd = 2.621
+ aigsd = 0.01077288
+ acnqsmod = 0
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ lvoff = -7.17621828e-9
+ tvfbsdoff = 0.022
+ njtsswg = 9
+ rbodymod = 0
+ lvsat = 0.001686942813
+ lvth0 = -7.292639699999997e-10
+ ntox = 1.0
+ ltvoff = -1.0782211e-10
+ pcit = -2.6560201e-16
+ pclm = 2.21669238
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ delta = 0.007595625
+ laigc = -6.9149623e-12
+ ckappad = 0.6
+ ckappas = 0.6
+ rnoia = 0
+ rnoib = 0
+ pdiblc1 = 0
+ pdiblc2 = 0.0068331981
+ phin = 0.15
+ pdiblcb = -0.3
+ )

.model nch_fs_17 nmos (
+ level = 54
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ pbswgd = 0.95
+ xtis = 3
+ pbswgs = 0.95
+ ijthdfwd = 0.01
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ aigbinv = 0.0163
+ cigc = 0.000625
+ voffl = 0
+ igcmod = 1
+ weta0 = -1.09928e-7
+ wetab = 2.7482e-8
+ ijthdrev = 0.01
+ cgidl = 0.22
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ poxedge = 1
+ k2we = 5e-5
+ pbswd = 0.8
+ pbsws = 0.8
+ dsub = 0.75
+ permod = 1
+ dtox = 2.7e-10
+ binunit = 2
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ pdits = 0
+ eta0 = 0.42133333
+ cigsd = 0.069865
+ etab = -0.29033333
+ lkvth0we = -2e-12
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ voffcv = -0.16942
+ wpemod = 1
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ acnqsmod = 0
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ tnoia = 0
+ rbodymod = 0
+ peta0 = 0.0
+ wketa = -3.7974654e-8
+ tpbsw = 0.0019
+ cjswd = 7.7408e-11
+ tpbswg = 0.0009
+ cjsws = 7.7408e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ wtvfbsdoff = 0
+ a0 = 2.2098167
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 72000
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.015086228
+ k3 = -1.8419
+ em = 1000000.0
+ wpdiblc2 = -6.449088e-9
+ ll = 0
+ lw = 0
+ u0 = 0.015266499999999999
+ w0 = 0
+ ua = -1.7855187e-9
+ ub = 2.0636167e-18
+ uc = 7.8391667e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ptvoff = 0
+ ww = 0
+ xw = 8.600000000000001e-9
+ njtsswg = 9
+ ltvfbsdoff = 0
+ waigsd = 3.0876027e-12
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ diomod = 1
+ scref = 1e-6
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.025656394
+ pigcd = 2.621
+ pdiblcb = -0.3
+ pditsd = 0
+ pditsl = 0
+ aigsd = 0.010772862
+ cjswgd = 2.66208e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.66208e-10
+ keta = 0.015093331
+ tvfbsdoff = 0.022
+ lvoff = -1.6e-11
+ wkvth0we = 2e-12
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lvsat = -0.0002
+ lcit = -8e-12
+ lvth0 = -4.8e-10
+ ptvfbsdoff = 0
+ kt1l = 0
+ mjswgd = 0.85
+ mjswgs = 0.85
+ trnqsmod = 0
+ delta = 0.007595625
+ bigbacc = 0.002588
+ tcjswg = 0.001
+ rnoia = 0
+ rnoib = 0
+ lint = 6.5375218e-9
+ kvth0we = 0.00018
+ lkt1 = -4.8e-10
+ lmax = 2.001e-5
+ lmin = 8.9991e-6
+ ngate = 8e+20
+ lintnoi = -1.5e-8
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ ngcon = 1
+ bigbinv = 0.004953
+ wpclm = 5.7423639e-7
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ rgatemod = 0
+ minv = -0.3
+ lub1 = -2.4000000000000004e-27
+ gbmin = 1e-12
+ tnjtsswg = 1
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ ndep = 1e+18
+ lwlc = 0
+ moin = 5.1
+ fprout = 300
+ nigc = 3.083
+ xrcrg1 = 12
+ xrcrg2 = 1
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ wtvoff = 9.3503662e-10
+ ntox = 1.0
+ pcit = -1.2000000000000001e-17
+ pclm = 0.629885
+ tvoff = 5.0359625e-5
+ capmod = 2
+ nfactor = 1
+ wku0we = 2e-11
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ phin = 0.15
+ mobmod = 0
+ pkt1 = 5.600000000000001e-17
+ ku0we = -0.0007
+ beta0 = 13
+ leta0 = 1.6000000000000003e-9
+ nigbacc = 10
+ rbdb = 50
+ prwb = 0
+ prwg = 0
+ pub1 = -3.2e-34
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ ags = 0.57720097
+ dlcig = 2.5e-9
+ rdsw = 100
+ bgidl = 2320000000.0
+ cjd = 0.001281008
+ cit = 6.2896875e-5
+ cjs = 0.001281008
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 9.8024918e-9
+ ijthsfwd = 0.01
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ nigbinv = 10
+ la0 = 0
+ jsd = 6.11e-7
+ dmcgt = 0
+ jss = 6.11e-7
+ lat = -0.00016
+ kt1 = -0.28314411
+ kt2 = -0.074391698
+ tcjsw = 0.000357
+ llc = 0
+ lln = 1
+ lu0 = 9.600000000000001e-12
+ mjd = 0.26
+ mjs = 0.26
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 0
+ ijthsrev = 0.01
+ nsd = 1e+20
+ pbd = 0.52
+ pat = -3.04e-11
+ pbs = 0.52
+ rshg = 15.6
+ pu0 = 1.8400000000000002e-18
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ prt = 0
+ pud = 0
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = -6.8749055e-10
+ ub1 = 1.0341951e-18
+ uc1 = 4.5339833e-11
+ fnoimod = 1
+ bigsd = 0.00125
+ tpb = 0.0014
+ wa0 = 7.159061e-7
+ eigbinv = 1.1
+ ute = -2.01925
+ wat = 0
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 3.760485e-9
+ wlc = 0
+ wln = 1
+ wu0 = -1.59669e-10
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -7.132277e-17
+ wub = 7.28273e-26
+ wuc = -1.167985e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ wvoff = 1.0181215e-9
+ wvsat = -0.0045771271
+ wvth0 = -1.19727395e-8
+ tnom = 25
+ toxe = 2.43e-9
+ waigc = 5.0140497e-11
+ toxm = 2.43e-9
+ toxref = 3e-9
+ cigbacc = 0.32875
+ xpart = 1
+ tnoimod = 0
+ wags = 1.0693246999999999e-7
+ egidl = 0.29734
+ pkvth0we = -1.3e-19
+ wcit = 4.8907306e-10
+ cigbinv = 0.006
+ voff = -0.11158375
+ ltvoff = 0
+ acde = 0.4
+ vsat = 106133.02
+ vfbsdoff = 0.02
+ wint = 0
+ pvfbsdoff = 0
+ vth0 = 0.32052953
+ wkt1 = 3.1515481e-8
+ wkt2 = 1.5939759e-8
+ wmax = 8.974e-7
+ aigc = 0.011740211
+ wmin = 5.374e-7
+ version = 4.5
+ tempmod = 0
+ lku0we = 2.5e-11
+ epsrox = 3.9
+ paramchk = 1
+ wua1 = 1.0731531e-15
+ wub1 = -9.2968455e-25
+ wuc1 = -1.4414309e-17
+ aigbacc = 0.02
+ rdsmod = 0
+ bigc = 0.001442
+ pvoff = 0
+ wute = 5.565105e-7
+ wwlc = 0
+ igbmod = 1
+ cdscb = 0
+ cdscd = 0
+ pvsat = -2.24e-11
+ wk2we = 5e-12
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ pvth0 = -1.2e-16
+ cdsc = 0
+ drout = 0.56
+ )

.model nch_fs_18 nmos (
+ level = 54
+ kt1l = 0
+ nigbacc = 10
+ tvoff = -0.0002433276
+ paigsd = 1.3573222e-22
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ lint = 6.5375218e-9
+ lkt1 = 8.5766405e-8
+ lkt2 = 5.1456509e-9
+ lmax = 8.9991e-6
+ lmin = 8.9908e-7
+ permod = 1
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ nigbinv = 10
+ ags = 0.5316128899999999
+ ku0we = -0.0007
+ ppdiblc2 = 1.9760389e-14
+ beta0 = 13
+ cjd = 0.001281008
+ leta0 = 1.6000000000000003e-9
+ cit = -0.00011782923
+ cjs = 0.001281008
+ minv = -0.3
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ lua1 = 1.38467e-15
+ lub1 = -1.4916591e-24
+ luc1 = 1.0686128e-16
+ dlc = 9.8024918e-9
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ ndep = 1e+18
+ lute = 1.0068051e-6
+ lwlc = 0
+ moin = 5.1
+ dlcig = 2.5e-9
+ voffcv = -0.16942
+ wpemod = 1
+ bgidl = 2320000000.0
+ la0 = -1.1479603e-6
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ nigc = 3.083
+ lat = 0.085185067
+ kt1 = -0.2927377
+ lk2 = -1.3507419e-8
+ kt2 = -0.074964073
+ llc = 0
+ lln = 1
+ lu0 = -1.9908396e-9
+ fnoimod = 1
+ mjd = 0.26
+ lua = -1.5028094e-16
+ mjs = 0.26
+ lub = -1.4426347e-25
+ luc = -5.2935673e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = -5.1713984e-13
+ eigbinv = 1.1
+ nsd = 1e+20
+ pbd = 0.52
+ pat = -3.04e-11
+ pbs = 0.52
+ pk2 = -1.6553107e-15
+ pu0 = 1.5413224e-17
+ prt = 0
+ noff = 2.7195
+ pua = -3.5916841e-23
+ pub = 6.5823852e-32
+ puc = 3.1761344e-23
+ pud = 0
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ pkvth0we = -1.3e-19
+ dmcgt = 0
+ rsh = 17.5
+ tcjsw = 0.000357
+ tcj = 0.00076
+ ua1 = -8.4151391e-10
+ ub1 = 1.1998524e-18
+ uc1 = 3.3453151e-11
+ tpb = 0.0014
+ wa0 = 7.7343e-7
+ pags = -1.4569295e-13
+ ute = -2.1312417
+ wtvfbsdoff = 0
+ wat = 0
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 3.944613e-9
+ wlc = 0
+ wln = 1
+ ntox = 1.0
+ wu0 = -1.6117881e-10
+ pcit = -6.4147523e-16
+ xgl = -1.09e-8
+ pclm = 0.629885
+ xgw = 0
+ wua = -6.7327571e-17
+ wub = 6.5505403e-26
+ wuc = -1.5212814e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ vfbsdoff = 0.02
+ tpbswg = 0.0009
+ bigsd = 0.00125
+ ltvfbsdoff = 0
+ phin = 0.15
+ cigbacc = 0.32875
+ wvoff = 8.2208115e-10
+ pkt1 = -6.946714e-14
+ pkt2 = -1.5079533e-14
+ paramchk = 1
+ tnoimod = 0
+ wvsat = -0.0045771271
+ wvth0 = -1.22760901e-8
+ ptvoff = -2.0299898e-15
+ waigsd = 3.0875876e-12
+ waigc = 5.030718e-11
+ rbdb = 50
+ pua1 = -1.044071e-21
+ prwb = 0
+ prwg = 0
+ pub1 = 9.8767081e-31
+ cigbinv = 0.006
+ puc1 = -4.3746501e-23
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ pute = -5.4971558e-13
+ diomod = 1
+ rdsw = 100
+ ptvfbsdoff = 0
+ lketa = -1.3350472e-7
+ ijthdfwd = 0.01
+ pditsd = 0
+ xpart = 1
+ pditsl = 0
+ cjswgd = 2.66208e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.66208e-10
+ version = 4.5
+ tempmod = 0
+ egidl = 0.29734
+ mjswgd = 0.85
+ mjswgs = 0.85
+ ijthdrev = 0.01
+ aigbacc = 0.02
+ a0 = 2.3375097
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ rshg = 15.6
+ at = 62506.667
+ cf = 8.15e-11
+ tcjswg = 0.001
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.016588722
+ k3 = -1.8419
+ em = 1000000.0
+ pvfbsdoff = 0
+ ll = 0
+ lw = 0
+ u0 = 0.015489017999999998
+ lpdiblc2 = -2.2119558e-8
+ w0 = 0
+ ua = -1.7688022e-9
+ ub = 2.0796638e-18
+ uc = 8.4279951e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ aigbinv = 0.0163
+ tnom = 25
+ pvoff = 1.7624031e-15
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ cdscb = 0
+ cdscd = 0
+ fprout = 300
+ pvsat = -2.24e-11
+ lkvth0we = -2e-12
+ wk2we = 5e-12
+ pvth0 = 2.6071227e-15
+ drout = 0.56
+ xrcrg1 = 12
+ xrcrg2 = 1
+ paigc = -1.4984839e-18
+ voffl = 0
+ poxedge = 1
+ acnqsmod = 0
+ wtvoff = 1.1608419e-9
+ wags = 1.2313859e-7
+ weta0 = -1.09928e-7
+ wetab = 2.7482e-8
+ wcit = 5.5909255e-10
+ binunit = 2
+ rbodymod = 0
+ voff = -0.1094379
+ acde = 0.4
+ capmod = 2
+ cgidl = 0.22
+ vsat = 106133.02
+ wint = 0
+ wku0we = 2e-11
+ vth0 = 0.31474059
+ wkt1 = 3.9248867000000004e-8
+ wkt2 = 1.7617127e-8
+ wmax = 8.974e-7
+ mobmod = 0
+ aigc = 0.011757817
+ wmin = 5.374e-7
+ pbswd = 0.8
+ pbsws = 0.8
+ wua1 = 1.1892901e-15
+ wub1 = -1.0395834e-24
+ wuc1 = -9.5481798e-18
+ wpdiblc2 = -8.647129e-9
+ bigc = 0.001442
+ wute = 6.1765795e-7
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ wwlc = 0
+ pdits = 0
+ cigsd = 0.069865
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ laigsd = -2.4859383e-16
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ wkvth0we = 2e-12
+ tnoia = 0
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ trnqsmod = 0
+ peta0 = 0.0
+ njtsswg = 9
+ wketa = -4.7550208e-8
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ tpbsw = 0.0019
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ cjswd = 7.7408e-11
+ cjsws = 7.7408e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.028116857
+ k2we = 5e-5
+ pdiblcb = -0.3
+ dsub = 0.75
+ dtox = 2.7e-10
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ rgatemod = 0
+ tnjtsswg = 1
+ toxref = 3e-9
+ eta0 = 0.42133333
+ etab = -0.29033333
+ bigbacc = 0.002588
+ scref = 1e-6
+ pigcd = 2.621
+ aigsd = 0.010772862
+ kvth0we = 0.00018
+ tvfbsdoff = 0.022
+ lvoff = -1.9307251000000003e-8
+ lintnoi = -1.5e-8
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ ltvoff = 2.6402481e-9
+ lvsat = -0.0002
+ lvth0 = 5.1562566e-8
+ delta = 0.007595625
+ laigc = -1.5827875e-10
+ rnoia = 0
+ rnoib = 0
+ lku0we = 2.5e-11
+ pketa = 8.6084224e-14
+ epsrox = 3.9
+ ngate = 8e+20
+ ngcon = 1
+ wvfbsdoff = 0
+ wpclm = 5.7423639e-7
+ lvfbsdoff = 0
+ rdsmod = 0
+ gbmin = 1e-12
+ igbmod = 1
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ pbswgd = 0.95
+ pbswgs = 0.95
+ nfactor = 1
+ ijthsfwd = 0.01
+ igcmod = 1
+ keta = 0.029943688
+ lags = 4.0983681e-7
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 1.6167277e-9
+ ijthsrev = 0.01
+ )

.model nch_fs_19 nmos (
+ level = 54
+ rgatemod = 0
+ tnom = 25
+ tnjtsswg = 1
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ pdits = 0
+ cigsd = 0.069865
+ voffcv = -0.16942
+ wpemod = 1
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ njtsswg = 9
+ wtvfbsdoff = 0
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ ltvfbsdoff = 0
+ ckappad = 0.6
+ ckappas = 0.6
+ wags = -7.91542e-7
+ pdiblc1 = 0
+ pdiblc2 = -0.019237439
+ pdiblcb = -0.3
+ wcit = -4.1548514e-10
+ tnoia = 0
+ voff = -0.12566406
+ acde = 0.4
+ peta0 = 0.0
+ vsat = 106133.02
+ wketa = 9.2259042e-8
+ wint = 0
+ tpbswg = 0.0009
+ vth0 = 0.37294179
+ tpbsw = 0.0019
+ wkt1 = -7.2513249e-8
+ wkt2 = 3.7202325e-9
+ wmax = 8.974e-7
+ bigbacc = 0.002588
+ cjswd = 7.7408e-11
+ aigc = 0.01160027
+ cjsws = 7.7408e-11
+ wmin = 5.374e-7
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ ptvfbsdoff = 0
+ kvth0we = 0.00018
+ ptvoff = 9.96032e-16
+ wua1 = 1.1798319e-17
+ wub1 = 1.8760115e-25
+ wuc1 = -8.2926019e-17
+ lintnoi = -1.5e-8
+ waigsd = 3.0878745e-12
+ bigbinv = 0.004953
+ bigc = 0.001442
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ wwlc = 0
+ diomod = 1
+ cdsc = 0
+ cgbo = 0
+ pditsd = 0
+ pditsl = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ cjswgd = 2.66208e-10
+ ijthsfwd = 0.01
+ scref = 1e-6
+ pku0we = -1.5e-18
+ cjswgs = 2.66208e-10
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ pigcd = 2.621
+ tvfbsdoff = 0.022
+ aigsd = 0.010772861
+ lvoff = -4.8659703e-9
+ mjswgd = 0.85
+ mjswgs = 0.85
+ lvsat = -0.0002
+ lvth0 = -2.365076e-10
+ ijthsrev = 0.01
+ tcjswg = 0.001
+ delta = 0.007595625
+ laigc = -1.8062176e-11
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ rnoia = 0
+ rnoib = 0
+ nfactor = 1
+ pketa = -3.8346008e-14
+ ngate = 8e+20
+ k2we = 5e-5
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ ngcon = 1
+ dsub = 0.75
+ wpclm = 5.7423639e-7
+ dtox = 2.7e-10
+ ppdiblc2 = -1.3176269e-14
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ fprout = 300
+ eta0 = 0.42133333
+ etab = -0.29033333
+ xrcrg1 = 12
+ xrcrg2 = 1
+ nigbacc = 10
+ a0 = 1.6362276
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 209176.65
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.013338797999999999
+ k3 = -1.8419
+ em = 1000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.014967274
+ w0 = 0
+ ua = -1.7708735e-9
+ ub = 1.8600147e-18
+ uc = 2.580063e-11
+ ud = 0
+ wtvoff = -2.2391826e-9
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ pkvth0we = -1.3e-19
+ nigbinv = 10
+ capmod = 2
+ wku0we = 2e-11
+ tvoff = 0.004406442
+ vfbsdoff = 0.02
+ mobmod = 0
+ ags = 2.397561
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ cjd = 0.001281008
+ cit = 0.0020125208
+ cjs = 0.001281008
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 9.8024918e-9
+ k3b = 1.9326
+ fnoimod = 1
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ eigbinv = 1.1
+ paramchk = 1
+ ku0we = -0.0007
+ beta0 = 13
+ la0 = -5.2381924e-7
+ leta0 = 1.6000000000000003e-9
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.04535122
+ kt1 = -0.12585017
+ lk2 = -1.0614987e-8
+ kt2 = -0.061139846
+ llc = 0
+ lln = 1
+ lu0 = -1.5264873e-9
+ mjd = 0.26
+ lua = -1.4843753e-16
+ mjs = 0.26
+ lub = 5.1224193e-26
+ luc = -8.8907704e-19
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 9.5948774e-14
+ nsd = 1e+20
+ pbd = 0.52
+ pat = -5.004813e-9
+ pbs = 0.52
+ laigsd = 2.1900591e-16
+ pk2 = -1.0578878e-15
+ pu0 = 1.3797723999999999e-17
+ dlcig = 2.5e-9
+ prt = 0
+ pua = 5.0063903e-23
+ pub = -8.0709098e-32
+ puc = -9.2074471e-24
+ pud = 0
+ bgidl = 2320000000.0
+ ijthdfwd = 0.01
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 7.2552224e-10
+ ub1 = -4.8701436e-19
+ uc1 = 1.8003493e-10
+ tpb = 0.0014
+ wa0 = 8.4566389e-8
+ ute = -1
+ wat = 0.0055892281
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 3.2733514e-9
+ keta = -0.17327473
+ cigbacc = 0.32875
+ wlc = 0
+ wln = 1
+ wu0 = -1.5936364000000001e-10
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -1.6393515e-16
+ wub = 2.3014917e-25
+ wuc = 3.0819536e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ dmcgt = 0
+ tcjsw = 0.000357
+ lags = -1.250857e-6
+ tnoimod = 0
+ jswd = 1.28e-13
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ jsws = 1.28e-13
+ lcit = -2.792838e-10
+ ijthdrev = 0.01
+ kt1l = 0
+ cigbinv = 0.006
+ lpdiblc2 = 2.0025765e-8
+ bigsd = 0.00125
+ lint = 6.5375218e-9
+ lkt1 = -6.2763496e-8
+ lkt2 = -7.1579117e-9
+ lmax = 8.9908e-7
+ lmin = 4.4908e-7
+ wvoff = 5.2999378e-9
+ lpe0 = 9.2e-8
+ version = 4.5
+ lpeb = 2.5e-7
+ tempmod = 0
+ wvsat = -0.0045771271
+ wvth0 = -1.0719922700000001e-8
+ minv = -0.3
+ lua1 = -9.9922063e-18
+ lub1 = 9.652288e-27
+ luc1 = -2.3596511e-17
+ toxref = 3e-9
+ waigc = 6.3350032e-11
+ ndep = 1e+18
+ aigbacc = 0.02
+ lwlc = 0
+ lkvth0we = -2e-12
+ moin = 5.1
+ lketa = 4.735968e-8
+ nigc = 3.083
+ xpart = 1
+ acnqsmod = 0
+ aigbinv = 0.0163
+ egidl = 0.29734
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ ltvoff = -1.4980468e-9
+ rbodymod = 0
+ pags = 6.6837277e-13
+ ntox = 1.0
+ pvfbsdoff = 0
+ pcit = 2.2589891e-16
+ pclm = 0.629885
+ phin = 0.15
+ lku0we = 2.5e-11
+ epsrox = 3.9
+ pkt1 = 3.0001144e-14
+ pkt2 = -2.7112972e-15
+ poxedge = 1
+ rdsmod = 0
+ igbmod = 1
+ wpdiblc2 = 2.8360352e-8
+ pvoff = -2.2228894e-15
+ binunit = 2
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ rbdb = 50
+ pua1 = 3.8966634e-24
+ prwb = 0
+ prwg = 0
+ pub1 = -1.0452346e-31
+ cdscb = 0
+ cdscd = 0
+ puc1 = 2.1559776e-23
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ pvsat = -2.24e-11
+ rbsb = 50
+ pvag = 1.2
+ pbswgd = 0.95
+ pbswgs = 0.95
+ wk2we = 5e-12
+ pvth0 = 1.2221337e-15
+ drout = 0.56
+ rdsw = 100
+ igcmod = 1
+ paigc = -1.3106622e-17
+ voffl = 0
+ weta0 = -1.09928e-7
+ wetab = 2.7482e-8
+ wkvth0we = 2e-12
+ trnqsmod = 0
+ cgidl = 0.22
+ rshg = 15.6
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ paigsd = -1.1957726e-22
+ permod = 1
+ pbswd = 0.8
+ pbsws = 0.8
+ )

.model nch_fs_20 nmos (
+ level = 54
+ rgatemod = 0
+ tnom = 25
+ tnjtsswg = 1
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ pdits = 0
+ cigsd = 0.069865
+ voffcv = -0.16942
+ wpemod = 1
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ njtsswg = 9
+ wtvfbsdoff = 0
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ ltvfbsdoff = 0
+ ckappad = 0.6
+ ckappas = 0.6
+ wags = 2.5066629999999997e-6
+ pdiblc1 = 0
+ pdiblc2 = 0.041730695
+ pdiblcb = -0.3
+ wcit = 1.9646632999999998e-10
+ tnoia = 0
+ voff = -0.11119538
+ acde = 0.4
+ peta0 = 0.0
+ vsat = 99029.765
+ wketa = 8.4379468e-9
+ wint = 0
+ tpbswg = 0.0009
+ vth0 = 0.38129989
+ tpbsw = 0.0019
+ wkt1 = 7.756762999999998e-9
+ wkt2 = -6.4493333e-9
+ wmax = 8.974e-7
+ bigbacc = 0.002588
+ cjswd = 7.7408e-11
+ aigc = 0.011620363
+ cjsws = 7.7408e-11
+ wmin = 5.374e-7
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ ptvfbsdoff = 0
+ kvth0we = 0.00018
+ ptvoff = -1.0913215e-16
+ wua1 = 2.6150731e-17
+ wub1 = -7.4432483e-26
+ wuc1 = -3.5091334e-17
+ lintnoi = -1.5e-8
+ waigsd = 3.0877293e-12
+ bigbinv = 0.004953
+ bigc = 0.001442
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ wwlc = 0
+ diomod = 1
+ cdsc = 0
+ cgbo = 0
+ pditsd = 0
+ pditsl = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ cjswgd = 2.66208e-10
+ ijthsfwd = 0.01
+ scref = 1e-6
+ pku0we = -1.5e-18
+ cjswgs = 2.66208e-10
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ pigcd = 2.621
+ tvfbsdoff = 0.022
+ aigsd = 0.010772861
+ lvoff = -1.123219e-8
+ mjswgd = 0.85
+ mjswgs = 0.85
+ lvsat = 0.0029254309
+ lvth0 = -3.914068e-9
+ ijthsrev = 0.01
+ tcjswg = 0.001
+ delta = 0.007595625
+ laigc = -2.6902885e-11
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ rnoia = 0
+ rnoib = 0
+ nfactor = 1
+ pketa = -1.4647263e-15
+ ngate = 8e+20
+ k2we = 5e-5
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ ngcon = 1
+ dsub = 0.75
+ wpclm = 5.7423639e-7
+ dtox = 2.7e-10
+ ppdiblc2 = 1.3236303e-15
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ fprout = 300
+ eta0 = 0.42133333
+ etab = -0.29033333
+ xrcrg1 = 12
+ xrcrg2 = 1
+ nigbacc = 10
+ a0 = -0.63009793
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 152816.98
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.012308169999999998
+ k3 = -1.8419
+ em = 1000000.0
+ ll = -1.18e-13
+ lw = 0
+ u0 = 0.012890664999999999
+ w0 = 0
+ ua = -2.0345741e-9
+ ub = 2.0265059e-18
+ uc = 2.0750138e-11
+ ud = 0
+ wtvoff = 2.7255415e-10
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ pkvth0we = -1.3e-19
+ nigbinv = 10
+ capmod = 2
+ wku0we = 2e-11
+ tvoff = 0.001369836
+ vfbsdoff = 0.02
+ mobmod = 0
+ ags = -5.5634702
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ cjd = 0.001281008
+ cit = 0.0010906361
+ cjs = 0.001281008
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 1.30529375e-8
+ k3b = 1.9326
+ fnoimod = 1
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ eigbinv = 1.1
+ paramchk = 1
+ ku0we = -0.0007
+ beta0 = 13
+ la0 = 4.73364e-7
+ leta0 = 1.6000000000000003e-9
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.020552964
+ kt1 = -0.257877
+ lk2 = -1.0161511e-8
+ kt2 = -0.061294719
+ llc = -1.18e-13
+ lln = 0.7
+ lu0 = -6.1277936e-10
+ mjd = 0.26
+ lua = -3.2409276e-17
+ mjs = 0.26
+ lub = -2.2031936e-26
+ luc = 1.3331392e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = -5.6835585e-13
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 5.4576901e-9
+ pbs = 0.52
+ laigsd = 6.148791e-17
+ pk2 = 5.7885716e-16
+ pu0 = 7.4108054e-18
+ dlcig = 2.5e-9
+ prt = 0
+ pua = 1.3198419e-23
+ pub = -1.7542132e-32
+ puc = -4.6237685e-24
+ pud = 0
+ bgidl = 2320000000.0
+ ijthdfwd = 0.01
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 7.2295613e-10
+ ub1 = -3.1143135e-19
+ uc1 = 1.5561971e-10
+ tpb = 0.0014
+ wa0 = 1.5943496e-6
+ ute = -1
+ wat = -0.018189188
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -4.4652352e-10
+ keta = -0.031454297
+ cigbacc = 0.32875
+ wlc = 0
+ wln = 1
+ wu0 = -1.4484792e-10
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -8.0149958e-17
+ wub = 8.6587882e-26
+ wuc = 2.0402085e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ dmcgt = 0
+ tcjsw = 0.000357
+ lags = 2.2519967e-6
+ tnoimod = 0
+ jswd = 1.28e-13
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ jsws = 1.28e-13
+ lcit = 1.2634545e-10
+ ijthdrev = 0.01
+ kt1l = 0
+ cigbinv = 0.006
+ lpdiblc2 = -6.8002141e-9
+ bigsd = 0.00125
+ lint = 9.7879675e-9
+ lkt1 = -4.6716909e-9
+ lkt2 = -7.0897675e-9
+ lmax = 4.4908e-7
+ lmin = 2.1577e-7
+ wvoff = -5.5871857e-9
+ lpe0 = 9.2e-8
+ version = 4.5
+ lpeb = 2.5e-7
+ tempmod = 0
+ wvsat = 0.0018584193
+ wvth0 = -9.6953081e-9
+ minv = -0.3
+ lua1 = -8.8631172e-18
+ lub1 = -6.7604234e-26
+ luc1 = -1.2853813e-17
+ toxref = 3e-9
+ waigc = 3.2137522e-11
+ ndep = 1e+18
+ aigbacc = 0.02
+ lwlc = 0
+ lkvth0we = -2e-12
+ moin = 5.1
+ lketa = -1.5041313e-8
+ nigc = 3.083
+ xpart = 1
+ acnqsmod = 0
+ aigbinv = 0.0163
+ egidl = 0.29734
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ ltvoff = -1.6194017e-10
+ rbodymod = 0
+ pags = -7.8283743e-13
+ ntox = 1.0
+ pvfbsdoff = 0
+ pcit = -4.3359735e-17
+ pclm = 0.629885
+ phin = 0.15
+ lku0we = 2.5e-11
+ epsrox = 3.9
+ pkt1 = -5.3176613e-15
+ pkt2 = 1.7633117e-15
+ poxedge = 1
+ rdsmod = 0
+ igbmod = 1
+ wpdiblc2 = -4.5939646e-9
+ pvoff = 2.567445e-15
+ binunit = 2
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ rbdb = 50
+ pua1 = -2.4183981e-24
+ prwb = 0
+ prwg = 0
+ pub1 = 1.0771342000000001e-32
+ cdscb = 0
+ cdscd = 0
+ puc1 = 5.125141e-25
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ pvsat = -2.8540404e-9
+ rbsb = 50
+ pvag = 1.2
+ pbswgd = 0.95
+ pbswgs = 0.95
+ wk2we = 5e-12
+ pvth0 = 7.713032399999999e-16
+ drout = 0.56
+ rdsw = 100
+ igcmod = 1
+ paigc = 6.2688273e-19
+ voffl = 0
+ weta0 = -1.09928e-7
+ wetab = 2.7482e-8
+ wkvth0we = 2e-12
+ trnqsmod = 0
+ cgidl = 0.22
+ rshg = 15.6
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ paigsd = -5.5708045e-23
+ permod = 1
+ pbswd = 0.8
+ pbsws = 0.8
+ )

.model nch_fs_21 nmos (
+ level = 54
+ acnqsmod = 0
+ dmcgt = 0
+ version = 4.5
+ tcjsw = 0.000357
+ ptvfbsdoff = 0
+ tempmod = 0
+ rbodymod = 0
+ tpbswg = 0.0009
+ aigbacc = 0.02
+ bigsd = 0.00125
+ wvoff = 4.2089489999999885e-10
+ ptvoff = 6.7086074e-18
+ wvsat = -0.0116031636
+ waigsd = 3.0872445e-12
+ aigbinv = 0.0163
+ wvth0 = 5.090214589999999e-9
+ wpdiblc2 = 3.4958017e-9
+ waigc = 1.7847398e-12
+ diomod = 1
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 2.66208e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.66208e-10
+ lketa = -3.6124213e-8
+ xpart = 1
+ keta = 0.068466797
+ egidl = 0.29734
+ mjswgd = 0.85
+ mjswgs = 0.85
+ wkvth0we = 2e-12
+ poxedge = 1
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ tcjswg = 0.001
+ lcit = 5.3521194000000004e-11
+ pvfbsdoff = 0
+ kt1l = 0
+ trnqsmod = 0
+ binunit = 2
+ lint = 9.7879675e-9
+ lkt1 = 2.3588251999999997e-10
+ lkt2 = 9.4878496e-10
+ lmax = 2.1577e-7
+ lmin = 9e-8
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ rgatemod = 0
+ minv = -0.3
+ lua1 = 1.428412e-17
+ pvoff = 1.2997136100000001e-15
+ lub1 = -6.5660104e-26
+ luc1 = -5.9196014e-18
+ tnjtsswg = 1
+ fprout = 300
+ ndep = 1e+18
+ cdscb = 0
+ cdscd = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ pvsat = -1.3647134000000064e-11
+ lwlc = 0
+ wk2we = 5e-12
+ pvth0 = -2.34841744e-15
+ moin = 5.1
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ drout = 0.56
+ nigc = 3.083
+ paigc = 7.0313197e-18
+ wtvoff = -2.7645419e-10
+ voffl = 0
+ noff = 2.7195
+ weta0 = -1.09928e-7
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ wetab = 2.7482e-8
+ lpclm = 5.9671804e-8
+ capmod = 2
+ wku0we = 2e-11
+ ntox = 1.0
+ cgidl = 0.22
+ pcit = -4.5161006999999997e-17
+ pclm = 0.34708024
+ mobmod = 0
+ njtsswg = 9
+ phin = 0.15
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ pkt1 = -1.0490175e-15
+ pkt2 = -1.739649e-15
+ pbswd = 0.8
+ pbsws = 0.8
+ a0 = 1.2892878
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 51380.779
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = -0.034882087
+ k3 = -1.8419
+ em = 1000000.0
+ ckappad = 0.6
+ ckappas = 0.6
+ ll = -1.18e-13
+ lw = 0
+ u0 = 0.011019764
+ w0 = 0
+ ua = -2.2703742e-9
+ ub = 2.053795462e-18
+ uc = 5.2246809e-11
+ ud = 0
+ pdiblc1 = 0
+ pdiblc2 = 0.010471563
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ pdiblcb = -0.3
+ rbdb = 50
+ pua1 = -9.0422848e-24
+ prwb = 0
+ pdits = 0
+ laigsd = -6.8373623e-17
+ prwg = 0
+ pub1 = 1.2957736e-32
+ puc1 = 4.9546192e-24
+ cigsd = 0.069865
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ rdsw = 100
+ ijthsfwd = 0.01
+ bigbacc = 0.002588
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ kvth0we = 0.00018
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ tnoia = 0
+ ijthsrev = 0.01
+ lintnoi = -1.5e-8
+ bigbinv = 0.004953
+ peta0 = 0.0
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ rshg = 15.6
+ wketa = -5.2502872e-8
+ tpbsw = 0.0019
+ cjswd = 7.7408e-11
+ cjsws = 7.7408e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ ppdiblc2 = -3.8331042e-16
+ toxref = 3e-9
+ tnom = 25
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ scref = 1e-6
+ tvfbsdoff = 0.022
+ pigcd = 2.621
+ aigsd = 0.010772862
+ nfactor = 1
+ ltvoff = 9.6416574e-11
+ wags = -1.203467e-6
+ lvoff = -9.038213999999995e-10
+ pkvth0we = -1.3e-19
+ wcit = 2.0500315999999998e-10
+ lvsat = -0.0004381747099999999
+ lvth0 = -6.676310299999999e-9
+ voff = -0.16014500000000004
+ acde = 0.4
+ delta = 0.007595625
+ laigc = -1.4310771e-11
+ vfbsdoff = 0.02
+ vsat = 114971.1026
+ wint = 0
+ vth0 = 0.39439110699999996
+ rnoia = 0
+ rnoib = 0
+ lku0we = 2.5e-11
+ wkt1 = -1.2473776800000001e-8
+ wkt2 = 1.0152376e-8
+ nigbacc = 10
+ wmax = 8.974e-7
+ epsrox = 3.9
+ aigc = 0.011560684
+ wmin = 5.374e-7
+ wvfbsdoff = 0
+ pketa = 1.139354e-14
+ lvfbsdoff = 0
+ ngate = 8e+20
+ rdsmod = 0
+ ngcon = 1
+ paramchk = 1
+ wpclm = 8.9560432e-7
+ igbmod = 1
+ wua1 = 5.7543559e-17
+ wub1 = -8.4794537e-26
+ wuc1 = -5.6143964e-17
+ gbmin = 1e-12
+ nigbinv = 10
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ bigc = 0.001442
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ wwlc = 0
+ pbswgd = 0.95
+ pbswgs = 0.95
+ cdsc = 0
+ igcmod = 1
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ ijthdfwd = 0.01
+ xtis = 3
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ fnoimod = 1
+ eigbinv = 1.1
+ ags = 5.1095
+ ijthdrev = 0.01
+ cjd = 0.001281008
+ cit = 0.0014357747
+ cjs = 0.001281008
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 1.30529375e-8
+ paigsd = 4.6587859e-23
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ tvoff = 0.00014539643
+ lpdiblc2 = -2.045371e-10
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ permod = 1
+ la0 = 6.8373618e-8
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = 0.0008500743
+ kt1 = -0.28113564
+ lk2 = -2.0436616e-10
+ kt2 = -0.099392124
+ llc = -1.18e-13
+ lln = 0.7
+ wtvfbsdoff = 0
+ lu0 = -2.1801917e-10
+ mjd = 0.26
+ lua = 1.7344554e-17
+ mjs = 0.26
+ lub = -2.7790142600000004e-26
+ luc = -5.3126584e-18
+ lud = 0
+ k2we = 5e-5
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = -4.6587862e-14
+ nsd = 1e+20
+ dsub = 0.75
+ pbd = 0.52
+ pat = -1.8236973e-9
+ pbs = 0.52
+ pk2 = -1.7344476e-15
+ cigbacc = 0.32875
+ dtox = 2.7e-10
+ ku0we = -0.0007
+ pu0 = 4.868211e-18
+ beta0 = 13
+ prt = 0
+ pua = 1.2335294e-23
+ pub = -1.88032504e-32
+ puc = -1.1996375e-24
+ pud = 0
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ leta0 = 1.6000000000000003e-9
+ ltvfbsdoff = 0
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 6.1325358e-10
+ ub1 = -3.2064524e-19
+ uc1 = 1.2275615e-10
+ tnoimod = 0
+ tpb = 0.0014
+ ppclm = -6.7808634e-14
+ wa0 = -8.7848444e-7
+ voffcv = -0.16942
+ wpemod = 1
+ ute = -1
+ wat = 0.016319757
+ eta0 = 0.42133333
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 1.0517006e-8
+ lkvth0we = -2e-12
+ etab = -0.29033333
+ wlc = 0
+ wln = 1
+ wu0 = -1.32797711e-10
+ xgl = -1.09e-8
+ xgw = 0
+ dlcig = 2.5e-9
+ wua = -7.6059319e-17
+ wub = 9.256491399999999e-26
+ wuc = 4.1739756e-18
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ bgidl = 2320000000.0
+ cigbinv = 0.006
+ )

.model nch_fs_22 nmos (
+ level = 54
+ phin = 0.15
+ cjswd = 7.7408e-11
+ cjsws = 7.7408e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ pkt1 = -2.3915509999999998e-15
+ pkt2 = 8.0276583e-16
+ ptvoff = -9.1490879e-17
+ nfactor = 1
+ paramchk = 1
+ waigsd = 3.0879615e-12
+ diomod = 1
+ rbdb = 50
+ pua1 = -1.6477593e-25
+ prwb = 0
+ prwg = 0
+ pub1 = 1.4213022e-32
+ puc1 = 1.092524e-23
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ pditsd = 0
+ pditsl = 0
+ rbsb = 50
+ pvag = 1.2
+ cjswgd = 2.66208e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.66208e-10
+ rdsw = 100
+ ijthdfwd = 0.01
+ scref = 1e-6
+ tvfbsdoff = 0.022
+ nigbacc = 10
+ pigcd = 2.621
+ aigsd = 0.010772861
+ mjswgd = 0.85
+ mjswgs = 0.85
+ lvoff = -5.128304999999991e-10
+ tcjswg = 0.001
+ lvsat = 0.0011237389840000002
+ ijthdrev = 0.01
+ lvth0 = -1.922596000000002e-10
+ nigbinv = 10
+ delta = 0.007595625
+ rshg = 15.6
+ laigc = -8.7106488e-12
+ lpdiblc2 = -4.1841324e-15
+ rnoia = 0
+ rnoib = 0
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ pketa = -2.7052976e-14
+ ngate = 8e+20
+ ngcon = 1
+ wpclm = 4.0103412e-7
+ fnoimod = 1
+ fprout = 300
+ eigbinv = 1.1
+ gbmin = 1e-12
+ tnom = 25
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ xrcrg1 = 12
+ xrcrg2 = 1
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ lkvth0we = -2e-12
+ wtvoff = 7.682212e-10
+ ags = 5.1095
+ cjd = 0.001281008
+ cit = 0.00076911293
+ cjs = 0.001281008
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ acnqsmod = 0
+ dlc = 3.26497e-9
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ wags = -1.203467e-6
+ capmod = 2
+ wcit = -2.3211370999999997e-10
+ cigbacc = 0.32875
+ rbodymod = 0
+ wku0we = 2e-11
+ la0 = -1.9182963e-7
+ voff = -0.164304478
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.0018542500800000001
+ acde = 0.4
+ kt1 = -0.33033037
+ lk2 = -1.3785596e-9
+ kt2 = -0.066210327
+ mobmod = 0
+ llc = 0
+ lln = 1
+ lu0 = -5.7555918999999996e-11
+ tnoimod = 0
+ mjd = 0.26
+ tvoff = 0.00053139469
+ lua = 2.7860169e-17
+ mjs = 0.26
+ lub = -2.7395085e-26
+ luc = 1.41139916e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ vsat = 98354.99900000001
+ njs = 1.02
+ pa0 = 2.0809981e-13
+ wint = 0
+ vth0 = 0.325411848
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 2.04854442e-9
+ pbs = 0.52
+ pk2 = 9.5324632e-16
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ wkt1 = 1.8084938999999998e-9
+ wkt2 = -1.689459e-8
+ pu0 = -7.071416999999997e-19
+ wmax = 8.974e-7
+ prt = 0
+ pua = -6.3654423e-24
+ pub = 7.034010899999999e-33
+ puc = -7.127418999999999e-24
+ pud = 0
+ cigbinv = 0.006
+ aigc = 0.011501109
+ wmin = 5.374e-7
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 8.1588744e-10
+ ub1 = -6.9089562e-19
+ uc1 = 1.6549472299999998e-10
+ tpb = 0.0014
+ wa0 = -3.5879278e-6
+ ute = -1
+ wat = -0.024874303599999998
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -1.8075483e-8
+ ku0we = -0.0007
+ wlc = 0
+ wln = 1
+ wu0 = -7.3485448e-11
+ xgl = -1.09e-8
+ xgw = 0
+ beta0 = 13
+ wua = 1.2288469e-16
+ wub = -1.8229956900000002e-25
+ wua1 = -3.6898024e-17
+ wuc = 6.7235478e-17
+ wud = 0
+ wub1 = -9.8148649e-26
+ wuc1 = -1.19661208e-16
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ leta0 = -9.226782e-9
+ wpdiblc2 = -5.8202891e-10
+ letab = -2.2164189e-8
+ version = 4.5
+ bigc = 0.001442
+ laigsd = 3.8113519e-17
+ tempmod = 0
+ wwlc = 0
+ ppclm = -2.1319035e-14
+ dlcig = 2.5e-9
+ cdsc = 0
+ bgidl = 2320000000.0
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ aigbacc = 0.02
+ xtis = 3
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ dmcgt = 0
+ tcjsw = 0.000357
+ wkvth0we = 2e-12
+ aigbinv = 0.0163
+ a0 = 4.0574074
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 80150.18699999999
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = -0.022390667
+ k3 = -1.8419
+ em = 1000000.0
+ ll = 0
+ lw = 0
+ trnqsmod = 0
+ u0 = 0.009312708
+ w0 = 0
+ ua = -2.3822425e-9
+ ub = 2.049592666e-18
+ uc = -1.5441968e-10
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ bigsd = 0.00125
+ wvoff = 3.044252900000001e-8
+ k2we = 5e-5
+ dsub = 0.75
+ dtox = 2.7e-10
+ wvsat = -0.017460162199999997
+ toxref = 3e-9
+ wvth0 = -3.853284300000001e-8
+ rgatemod = 0
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ tnjtsswg = 1
+ poxedge = 1
+ waigc = 1.9067031e-10
+ eta0 = 0.53651186
+ etab = -0.054544089
+ binunit = 2
+ lketa = 6.7720908e-8
+ xpart = 1
+ ltvoff = 6.0132739e-11
+ egidl = 0.29734
+ pvfbsdoff = 0
+ lku0we = 2.5e-11
+ epsrox = 3.9
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ rdsmod = 0
+ igbmod = 1
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ pvoff = -1.5223199999999999e-15
+ pbswgd = 0.95
+ pbswgs = 0.95
+ cdscb = 0
+ cdscd = 0
+ pvsat = 5.369107899999995e-10
+ wk2we = 5e-12
+ igcmod = 1
+ pvth0 = 1.7521499999999999e-15
+ drout = 0.56
+ paigc = -1.0723924e-17
+ ijthsfwd = 0.01
+ njtsswg = 9
+ voffl = 0
+ keta = -1.0362685
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ weta0 = -2.7932191e-7
+ wetab = 6.5877739e-8
+ wtvfbsdoff = 0
+ lpclm = -1.3225653e-8
+ ckappad = 0.6
+ ckappas = 0.6
+ jswd = 1.28e-13
+ pdiblc1 = 0
+ jsws = 1.28e-13
+ pdiblc2 = 0.0082956805
+ lcit = 1.1618741e-10
+ paigsd = -2.0809977e-23
+ pdiblcb = -0.3
+ ijthsrev = 0.01
+ kt1l = 0
+ cgidl = 0.22
+ ltvfbsdoff = 0
+ permod = 1
+ lint = 0
+ lkt1 = 4.8601869e-9
+ lkt2 = -2.1703039e-9
+ lmax = 9e-8
+ lmin = 5.4e-8
+ pbswd = 0.8
+ pbsws = 0.8
+ bigbacc = 0.002588
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ ppdiblc2 = 5.6582339e-21
+ minv = -0.3
+ kvth0we = 0.00018
+ lua1 = -4.7634626e-18
+ lub1 = -3.0856569e-26
+ luc1 = -9.937027189999999e-18
+ voffcv = -0.16942
+ wpemod = 1
+ pdits = 0
+ ndep = 1e+18
+ lintnoi = -1.5e-8
+ cigsd = 0.069865
+ ptvfbsdoff = 0
+ lwlc = 0
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ moin = 5.1
+ vtsswgs = 4.2
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ nigc = 3.083
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ pkvth0we = -1.3e-19
+ tnoia = 0
+ tpbswg = 0.0009
+ peta0 = 1.5923028e-14
+ ntox = 1.0
+ pcit = -4.072021500000001e-18
+ petab = -3.6091995e-15
+ pclm = 1.1225851
+ vfbsdoff = 0.02
+ wketa = 3.5650261e-7
+ tpbsw = 0.0019
+ )

.model nch_fs_23 nmos (
+ level = 54
+ pditsl = 0
+ cjswgd = 2.66208e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.66208e-10
+ cdsc = 0
+ lketa = -2.0578185e-8
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ ijthsfwd = 0.01
+ xtid = 3
+ xtis = 3
+ xpart = 1
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ mjswgd = 0.85
+ mjswgs = 0.85
+ egidl = 0.29734
+ tcjswg = 0.001
+ pvfbsdoff = 0
+ ijthsrev = 0.01
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ njtsswg = 9
+ k2we = 5e-5
+ dsub = 0.75
+ dtox = 2.7e-10
+ fprout = 300
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ xrcrg1 = 12
+ xrcrg2 = 1
+ pvoff = -3.925098540000001e-15
+ ckappad = 0.6
+ ckappas = 0.6
+ cdscb = 0
+ pdiblc1 = 0
+ pdiblc2 = 0.0082956083
+ cdscd = 0
+ pdiblcb = -0.3
+ pvsat = 4.008919351e-9
+ eta0 = 0.49180426
+ etab = -1.1686036
+ wk2we = 5e-12
+ pvth0 = 4.623404900000001e-15
+ drout = 0.56
+ wtvoff = -4.625476e-9
+ paigc = -1.7630641e-18
+ voffl = 0
+ weta0 = 1.6706711e-7
+ capmod = 2
+ bigbacc = 0.002588
+ wetab = -6.7375536e-8
+ pkvth0we = -1.3e-19
+ lpclm = -4.9784452e-8
+ wku0we = 2e-11
+ mobmod = 0
+ kvth0we = 0.00018
+ cgidl = 0.22
+ vfbsdoff = 0.02
+ lintnoi = -1.5e-8
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ pbswd = 0.8
+ pbsws = 0.8
+ paramchk = 1
+ laigsd = -3.1577826e-17
+ pdits = 0
+ cigsd = 0.069865
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ ijthdfwd = 0.01
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ keta = 0.48612964
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ nfactor = 1
+ tnoia = 0
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ ijthdrev = 0.01
+ lcit = 3.7801345e-10
+ peta0 = -9.9675358e-15
+ kt1l = 0
+ petab = 4.1194905e-15
+ wketa = -1.8474011e-7
+ tpbsw = 0.0019
+ lint = 0
+ cjswd = 7.7408e-11
+ cjsws = 7.7408e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ lkt1 = -1.5354128e-8
+ lkt2 = -1.4213753e-9
+ lmax = 5.4e-8
+ lmin = 4.5e-8
+ nigbacc = 10
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ toxref = 3e-9
+ minv = -0.3
+ lua1 = 7.7308837e-17
+ lub1 = -1.6131426200000002e-25
+ luc1 = -7.236573999999998e-18
+ ndep = 1e+18
+ lkvth0we = -2e-12
+ nigbinv = 10
+ lwlc = 0
+ moin = 5.1
+ a0 = 11.080765
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 31524.241299999994
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ tvfbsdoff = 0.022
+ k2 = 0.011547898
+ k3 = -1.8419
+ em = 1000000.0
+ ll = 0
+ lw = 0
+ u0 = -0.00096107274
+ scref = 1e-6
+ nigc = 3.083
+ w0 = 0
+ ua = -5.2066121e-9
+ ub = 5.20056154e-18
+ uc = 2.7090556e-10
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ pigcd = 2.621
+ aigsd = 0.010772862
+ ltvoff = -1.4697355e-10
+ acnqsmod = 0
+ lvoff = 1.5958058999999975e-9
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ fnoimod = 1
+ lvsat = -0.00556709637
+ rbodymod = 0
+ lvth0 = -4.0736673000000004e-9
+ eigbinv = 1.1
+ ntox = 1.0
+ delta = 0.007595625
+ pcit = 1.0096077e-17
+ lku0we = 2.5e-11
+ pclm = 1.7529092
+ laigc = -1.8175152e-11
+ epsrox = 3.9
+ rnoia = 0
+ rnoib = 0
+ wvfbsdoff = 0
+ phin = 0.15
+ lvfbsdoff = 0
+ rdsmod = 0
+ pketa = 4.339103e-15
+ igbmod = 1
+ ngate = 8e+20
+ pkt1 = 1.1996454999999999e-14
+ pkt2 = 3.1759909e-15
+ ngcon = 1
+ wpclm = -7.2697212e-7
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ wpdiblc2 = -5.8193135e-10
+ pbswgd = 0.95
+ gbmin = 1e-12
+ pbswgs = 0.95
+ cigbacc = 0.32875
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ ags = 5.1095
+ rbdb = 50
+ pua1 = -6.2039198e-23
+ prwb = 0
+ prwg = 0
+ pub1 = 1.08120889e-31
+ puc1 = 1.0847755599999997e-23
+ igcmod = 1
+ wtvfbsdoff = 0
+ cjd = 0.001281008
+ cit = -0.0037451293
+ cjs = 0.001281008
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ dlc = 3.26497e-9
+ k3b = 1.9326
+ tnoimod = 0
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ rdsw = 100
+ ltvfbsdoff = 0
+ cigbinv = 0.006
+ la0 = -5.9918439e-7
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = 0.0009660548200000002
+ kt1 = 0.018192305
+ lk2 = -3.3469964e-9
+ kt2 = -0.079122889
+ llc = 0
+ lln = 1
+ lu0 = 5.3832336e-10
+ mjd = 0.26
+ lua = 1.9167361e-16
+ mjs = 0.26
+ lub = -2.101512744e-25
+ luc = -1.0554871600000002e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 1.4611928e-13
+ wkvth0we = 2e-12
+ nsd = 1e+20
+ pbd = 0.52
+ pat = -1.47593358e-9
+ pbs = 0.52
+ pk2 = 2.1253177e-15
+ paigsd = 1.0451534e-29
+ pu0 = -5.5765924e-17
+ prt = 0
+ pua = -7.1470289e-23
+ pub = 9.665873609999999e-32
+ puc = 4.556057900000002e-24
+ pud = 0
+ version = 4.5
+ rsh = 17.5
+ trnqsmod = 0
+ tcj = 0.00076
+ ua1 = -5.9915221e-10
+ ub1 = 1.5583749700000001e-18
+ uc1 = 1.1893518999999988e-10
+ rshg = 15.6
+ tempmod = 0
+ tvoff = 0.0041021928
+ tpb = 0.0014
+ wa0 = -2.5192978e-6
+ permod = 1
+ ute = -1
+ wat = 0.035892558
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -3.8283609e-8
+ xjbvd = 1
+ xjbvs = 1
+ wlc = 0
+ wln = 1
+ lk2we = -1.5e-12
+ wu0 = 8.758039e-10
+ xgl = -1.09e-8
+ xgw = 0
+ wua = 1.2453821e-15
+ wub = -1.72755342e-24
+ wuc = -1.3420376999999993e-16
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ ptvfbsdoff = 0
+ aigbacc = 0.02
+ ku0we = -0.0007
+ beta0 = 13
+ rgatemod = 0
+ leta0 = -6.633740899999999e-9
+ letab = 4.245126e-8
+ voffcv = -0.16942
+ wpemod = 1
+ tnom = 25
+ tnjtsswg = 1
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ aigbinv = 0.0163
+ ppclm = 4.4105328e-14
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ wags = -1.203467e-6
+ dmcgt = 0
+ tcjsw = 0.000357
+ wcit = -4.763912600000001e-10
+ tpbswg = 0.0009
+ voff = -0.20066027000000003
+ acde = 0.4
+ poxedge = 1
+ vsat = 213714.23399999997
+ wint = 0
+ vth0 = 0.39233267
+ bigsd = 0.00125
+ binunit = 2
+ wkt1 = -2.4626057999999997e-7
+ wkt2 = -5.7812263e-8
+ wmax = 8.974e-7
+ aigc = 0.01166429
+ wmin = 5.374e-7
+ ptvoff = 2.2134356e-16
+ wvoff = 7.186973409999998e-8
+ waigsd = 3.0876027e-12
+ wvsat = -0.07732237357
+ wua1 = 1.0299024e-15
+ wub1 = -1.71724981e-24
+ wuc1 = -1.1832528899999998e-16
+ wvth0 = -8.803723199999998e-8
+ diomod = 1
+ bigc = 0.001442
+ waigc = 3.6172725e-11
+ wwlc = 0
+ pditsd = 0
+ )

.model nch_fs_24 nmos (
+ level = 54
+ lvsat = -0.0033743501999999996
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lvth0 = 5.361552700000001e-9
+ lcit = -3.5239012000000003e-10
+ trnqsmod = 0
+ kt1l = 0
+ cigbacc = 0.32875
+ delta = 0.007595625
+ laigc = -7.4258513e-12
+ rnoia = 0
+ rnoib = 0
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ tnoimod = 0
+ lint = 0
+ lkt1 = 5.314149e-10
+ lkt2 = 6.4873536e-9
+ lmax = 4.5e-8
+ pketa = 3.05233408e-14
+ ags = 5.1095
+ ngate = 8e+20
+ lmin = 3.6e-8
+ cigbinv = 0.006
+ ngcon = 1
+ lpe0 = 9.2e-8
+ cjd = 0.001281008
+ cit = 0.011161064
+ fprout = 300
+ cjs = 0.001281008
+ clc = 1e-7
+ wpclm = 9.524622100000001e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ lpeb = 2.5e-7
+ dlc = 3.26497e-9
+ k3b = 1.9326
+ xrcrg1 = 12
+ xrcrg2 = 1
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ rgatemod = 0
+ gbmin = 1e-12
+ minv = -0.3
+ tnjtsswg = 1
+ lua1 = -6.7547343e-17
+ lub1 = 1.27409254e-25
+ luc1 = 1.834266e-17
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ ndep = 1e+18
+ la0 = -5.581062559999999e-7
+ version = 4.5
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.00183504779
+ wtvoff = -5.6534448e-10
+ lwlc = 0
+ kt1 = -0.30600245
+ lk2 = -3.4047834e-9
+ kt2 = -0.24052552
+ llc = 0
+ moin = 5.1
+ lln = 1
+ lu0 = 9.4722495e-10
+ tempmod = 0
+ mjd = 0.26
+ lua = 1.9963428e-16
+ mjs = 0.26
+ lub = -1.86515944e-25
+ luc = -1.3855022100000003e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 1.41312605e-13
+ nigc = 3.083
+ nsd = 1e+20
+ pbd = 0.52
+ pat = -2.0050081000000007e-10
+ pbs = 0.52
+ pk2 = 1.540171e-16
+ pu0 = -4.9210101e-16
+ prt = 0
+ pua = -1.24177601e-22
+ pub = 1.2166737845000001e-31
+ puc = -3.231882900000001e-24
+ pud = 0
+ aigbacc = 0.02
+ capmod = 2
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 2.3570964e-9
+ ub1 = -4.3339417e-18
+ uc1 = -4.0308999999999995e-10
+ tpb = 0.0014
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ wku0we = 2e-11
+ wa0 = -2.4212027299999997e-6
+ ute = -1
+ wat = 0.009863318999999999
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 1.947015e-9
+ wlc = 0
+ wln = 1
+ wu0 = 9.780604500000001e-9
+ xgl = -1.09e-8
+ mobmod = 0
+ xgw = 0
+ wua = 2.32104147e-15
+ wub = -2.2379339299999998e-24
+ wuc = 2.4733810000000014e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ ntox = 1.0
+ pcit = 4.85396743e-16
+ pclm = 0.021884800000000038
+ tvoff = 0.0045807103
+ aigbinv = 0.0163
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ phin = 0.15
+ pkt1 = -5.2425624e-15
+ pkt2 = -2.9889728e-15
+ ku0we = -0.0007
+ beta0 = 13
+ laigsd = 2.1777751e-17
+ leta0 = 7.6237771e-9
+ letab = 3.2196399e-8
+ ppclm = -3.8186956000000005e-14
+ rbdb = 50
+ pua1 = 5.0551945e-23
+ prwb = 0
+ prwg = 0
+ pub1 = -9.600911599999999e-32
+ puc1 = -1.81613879e-23
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ poxedge = 1
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ rdsw = 100
+ ijthsfwd = 0.01
+ binunit = 2
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ dmcgt = 0
+ tcjsw = 0.000357
+ ijthsrev = 0.01
+ rshg = 15.6
+ bigsd = 0.00125
+ wvoff = -2.5396920999999984e-8
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ toxref = 3e-9
+ wvsat = -0.03971696100000001
+ wvth0 = 7.441037299999997e-8
+ tnom = 25
+ waigc = -1.3685053e-10
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ lketa = -4.89346675e-8
+ xpart = 1
+ ltvoff = -1.7042091e-10
+ egidl = 0.29734
+ njtsswg = 9
+ wags = -1.203467e-6
+ pkvth0we = -1.3e-19
+ pvfbsdoff = 0
+ wcit = -1.01764014e-8
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ voff = -0.003529144999999956
+ lku0we = 2.5e-11
+ acde = 0.4
+ ckappad = 0.6
+ epsrox = 3.9
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.0082956083
+ vfbsdoff = 0.02
+ pdiblcb = -0.3
+ vsat = 168964.27599999998
+ wint = 0
+ vth0 = 0.19977726499999998
+ wkt1 = 1.0555611e-7
+ wkt2 = 6.8003321e-8
+ rdsmod = 0
+ wtvfbsdoff = 0
+ wmax = 8.974e-7
+ aigc = 0.011444916
+ wmin = 5.374e-7
+ igbmod = 1
+ a0 = 10.24243689
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 88689.602
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.012727223
+ k3 = -1.8419
+ em = 1000000.0
+ ll = 0
+ lw = 0
+ u0 = -0.009305995800000001
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ paramchk = 1
+ w0 = 0
+ ua = -5.369074800000001e-9
+ ub = 4.718207719999999e-18
+ uc = 3.3825556e-10
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ ltvfbsdoff = 0
+ pbswgd = 0.95
+ pbswgs = 0.95
+ wua1 = -1.2678761e-15
+ wub1 = 2.44866871e-24
+ wuc1 = 4.7369808e-16
+ bigbacc = 0.002588
+ pvoff = 8.409683299999991e-16
+ bigc = 0.001442
+ igcmod = 1
+ wwlc = 0
+ cdscb = 0
+ cdscd = 0
+ kvth0we = 0.00018
+ pvsat = 2.1662543300000005e-9
+ wk2we = 5e-12
+ pvth0 = -3.336525699999999e-15
+ drout = 0.56
+ cdsc = 0
+ lintnoi = -1.5e-8
+ paigc = 6.7150752e-18
+ cgbo = 0
+ ijthdfwd = 0.01
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ voffl = 0
+ cigc = 0.000625
+ ptvfbsdoff = 0
+ weta0 = -1.6294544599999998e-7
+ wetab = 1.0177792e-7
+ paigsd = 4.9710031e-30
+ lpclm = 3.5035747999999996e-8
+ ijthdrev = 0.01
+ cgidl = 0.22
+ permod = 1
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ pbswd = 0.8
+ pbsws = 0.8
+ k2we = 5e-5
+ dsub = 0.75
+ dtox = 2.7e-10
+ voffcv = -0.16942
+ wpemod = 1
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ nfactor = 1
+ pdits = 0
+ cigsd = 0.069865
+ eta0 = 0.20083450200000003
+ lkvth0we = -2e-12
+ etab = -0.95932067
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ acnqsmod = 0
+ nigbacc = 10
+ tpbswg = 0.0009
+ tnoia = 0
+ rbodymod = 0
+ peta0 = 6.20307972e-15
+ petab = -4.1690291e-15
+ wketa = -7.1911233e-7
+ tpbsw = 0.0019
+ nigbinv = 10
+ cjswd = 7.7408e-11
+ cjsws = 7.7408e-11
+ ptvoff = 2.2397114e-17
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ waigsd = 3.0876027e-12
+ diomod = 1
+ wpdiblc2 = -5.8193135e-10
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 2.66208e-10
+ pku0we = -1.5e-18
+ fnoimod = 1
+ cjswgs = 2.66208e-10
+ eigbinv = 1.1
+ tvfbsdoff = 0.022
+ scref = 1e-6
+ pigcd = 2.621
+ mjswgd = 0.85
+ aigsd = 0.010772861
+ mjswgs = 0.85
+ keta = 1.06483334
+ tcjswg = 0.001
+ lvoff = -8.06362e-9
+ wkvth0we = 2e-12
+ )

.model nch_fs_25 nmos (
+ level = 54
+ fprout = 300
+ xrcrg1 = 12
+ xrcrg2 = 1
+ pvoff = 0
+ tnom = 25
+ cdscb = 0
+ cdscd = 0
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ wtvoff = 0
+ pvsat = -2.24e-11
+ lkvth0we = -2e-12
+ wk2we = 5e-12
+ pvth0 = -1.2e-16
+ drout = 0.56
+ voffl = 0
+ capmod = 2
+ acnqsmod = 0
+ wku0we = 2e-11
+ weta0 = -1.1162667e-8
+ wags = -7.346904000000001e-8
+ wetab = 2.2325333e-8
+ mobmod = 0
+ wcit = 3.3636880000000003e-10
+ rbodymod = 0
+ nfactor = 1
+ voff = -0.13478422
+ acde = 0.4
+ cgidl = 0.22
+ vsat = 102889.02
+ wint = 0
+ vth0 = 0.33700512
+ wkt1 = -2.6570593870000003e-9
+ wkt2 = -5.3296152e-9
+ wmax = 5.374e-7
+ aigc = 0.011779434
+ wmin = 2.674e-7
+ pbswd = 0.8
+ pbsws = 0.8
+ wua1 = -1.874362e-16
+ nigbacc = 10
+ wub1 = 1.1464267e-25
+ wuc1 = -2.7527136e-17
+ wpdiblc2 = 4.9914968e-9
+ bigc = 0.001442
+ pdits = 0
+ wwlc = 0
+ cigsd = 0.069865
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ nigbinv = 10
+ xtis = 3
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ wkvth0we = 2e-12
+ tnoia = 0
+ trnqsmod = 0
+ peta0 = 0.0
+ fnoimod = 1
+ wketa = 1.6322115e-8
+ eigbinv = 1.1
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ tpbsw = 0.0019
+ dmdg = 0
+ cjswd = 7.7408e-11
+ cjsws = 7.7408e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ toxref = 3e-9
+ k2we = 5e-5
+ dsub = 0.75
+ dtox = 2.7e-10
+ rgatemod = 0
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ tnjtsswg = 1
+ tvfbsdoff = 0.022
+ eta0 = 0.24044444
+ etab = -0.28088889
+ cigbacc = 0.32875
+ ltvoff = 0
+ scref = 1e-6
+ pigcd = 2.621
+ tnoimod = 0
+ aigsd = 0.010772818
+ wtvfbsdoff = 0
+ lvoff = -1.6e-11
+ cigbinv = 0.006
+ lvsat = -0.0002
+ lku0we = 2.5e-11
+ lvth0 = -4.8e-10
+ ltvfbsdoff = 0
+ epsrox = 3.9
+ delta = 0.007595625
+ ags = 0.9076066700000001
+ wvfbsdoff = 0
+ cjd = 0.001281008
+ cit = 0.000342575
+ version = 4.5
+ cjs = 0.001281008
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ lvfbsdoff = 0
+ rnoia = 0
+ rnoib = 0
+ rdsmod = 0
+ dlc = 9.8024918e-9
+ k3b = 1.9326
+ tempmod = 0
+ igbmod = 1
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ ngate = 8e+20
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ ngcon = 1
+ la0 = 0
+ wpclm = 9.3989653e-8
+ pbswgd = 0.95
+ jsd = 6.11e-7
+ pbswgs = 0.95
+ jss = 6.11e-7
+ lat = -0.00016
+ aigbacc = 0.02
+ kt1 = -0.22055704
+ kt2 = -0.0354368
+ llc = 0
+ lln = 1
+ lu0 = 9.600000000000001e-12
+ mjd = 0.26
+ mjs = 0.26
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ gbmin = 1e-12
+ njs = 1.02
+ pa0 = 0
+ igcmod = 1
+ nsd = 1e+20
+ pbd = 0.52
+ pat = -3.04e-11
+ jswgd = 1.28e-13
+ ptvfbsdoff = 0
+ pbs = 0.52
+ jswgs = 1.28e-13
+ pu0 = 1.8400000000000002e-18
+ prt = 0
+ pud = 0
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 1.6212811e-9
+ ub1 = -8.7849211e-19
+ uc1 = 6.9356e-11
+ tpb = 0.0014
+ aigbinv = 0.0163
+ wa0 = -1.17208e-8
+ ijthsfwd = 0.01
+ ute = -1
+ wat = 0.071441067
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 1.8596306e-9
+ wlc = 0
+ wln = 1
+ wu0 = -1.3197067000000002e-9
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -1.3097991e-16
+ wub = 9.54408e-26
+ wuc = -2.4557867e-18
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ keta = -0.084351302
+ a0 = 3.5424667
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = -58844.444
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.018567646
+ k3 = -1.8419
+ em = 1000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.017391111
+ jswd = 1.28e-13
+ w0 = 0
+ jsws = 1.28e-13
+ ijthsrev = 0.01
+ ua = -1.6762565e-9
+ ub = 2.0222e-18
+ uc = 6.1497778e-11
+ ud = 0
+ lcit = -8e-12
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ permod = 1
+ kt1l = 0
+ tvoff = 0.0017628809
+ xjbvd = 1
+ xjbvs = 1
+ poxedge = 1
+ lk2we = -1.5e-12
+ lint = 6.5375218e-9
+ lkt1 = -4.8e-10
+ lmax = 2.001e-5
+ binunit = 2
+ lmin = 8.9991e-6
+ lpe0 = 9.2e-8
+ voffcv = -0.16942
+ wpemod = 1
+ lpeb = 2.5e-7
+ ku0we = -0.0007
+ beta0 = 13
+ leta0 = 1.6000000000000003e-9
+ minv = -0.3
+ lub1 = -2.4000000000000004e-27
+ ndep = 1e+18
+ lwlc = 0
+ dlcig = 2.5e-9
+ moin = 5.1
+ bgidl = 2320000000.0
+ nigc = 3.083
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ noff = 2.7195
+ dmcgt = 0
+ noia = 3.11e+42
+ noib = 1.22e+22
+ pkvth0we = -1.3e-19
+ noic = 45200000.0
+ tpbswg = 0.0009
+ tcjsw = 0.000357
+ ntox = 1.0
+ pcit = -1.2000000000000001e-17
+ pclm = 1.5094578
+ vfbsdoff = 0.02
+ bigsd = 0.00125
+ ptvoff = 0
+ phin = 0.15
+ waigsd = 3.1112026e-12
+ wvoff = 1.3685577e-8
+ pkt1 = 5.600000000000001e-17
+ paramchk = 1
+ diomod = 1
+ wvsat = -0.0028059037
+ wvth0 = -2.0968414e-8
+ njtsswg = 9
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 2.66208e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.66208e-10
+ waigc = 2.8724444e-11
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ rbdb = 50
+ prwb = 0
+ prwg = 0
+ pub1 = -3.2e-34
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.0047029422
+ rdsw = 100
+ pdiblcb = -0.3
+ ijthdfwd = 0.01
+ mjswgd = 0.85
+ xpart = 1
+ mjswgs = 0.85
+ tcjswg = 0.001
+ egidl = 0.29734
+ pvfbsdoff = 0
+ bigbacc = 0.002588
+ ijthdrev = 0.01
+ rshg = 15.6
+ kvth0we = 0.00018
+ lintnoi = -1.5e-8
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ )

.model nch_fs_26 nmos (
+ level = 54
+ poxedge = 1
+ capmod = 2
+ wku0we = 2e-11
+ binunit = 2
+ mobmod = 0
+ pkvth0we = -1.3e-19
+ tvoff = 0.0019388906
+ vfbsdoff = 0.02
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ laigsd = -2.019482e-16
+ paramchk = 1
+ ku0we = -0.0007
+ beta0 = 13
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ leta0 = 1.6000000000000003e-9
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ ijthdfwd = 0.01
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ keta = -0.091670067
+ dmcgt = 0
+ tcjsw = 0.000357
+ lags = -1.7808411e-7
+ njtsswg = 9
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ ijthdrev = 0.01
+ lcit = 6.5978289e-10
+ kt1l = 0
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ lpdiblc2 = 2.6261368e-8
+ bigsd = 0.00125
+ ckappad = 0.6
+ ckappas = 0.6
+ lint = 6.5375218e-9
+ pdiblc1 = 0
+ pdiblc2 = 0.0017817666
+ toxref = 3e-9
+ pdiblcb = -0.3
+ lkt1 = 8.5772759e-9
+ lkt2 = -2.1662043e-8
+ lmax = 8.9991e-6
+ wvoff = 1.395365e-8
+ lmin = 8.9908e-7
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ wvsat = -0.0028059037
+ wvth0 = -2.1316317000000002e-8
+ minv = -0.3
+ wtvfbsdoff = 0
+ lua1 = -8.9279603e-16
+ lub1 = 6.8304226e-25
+ luc1 = -5.9256432e-18
+ waigc = 2.989874e-11
+ bigbacc = 0.002588
+ ndep = 1e+18
+ lkvth0we = -2e-12
+ lwlc = 0
+ moin = 5.1
+ ltvoff = -1.582327e-9
+ ltvfbsdoff = 0
+ lketa = 6.5795695e-8
+ kvth0we = 0.00018
+ nigc = 3.083
+ xpart = 1
+ lintnoi = -1.5e-8
+ acnqsmod = 0
+ pvfbsdoff = 0
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ egidl = 0.29734
+ vtsswgs = 4.2
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ lku0we = 2.5e-11
+ rbodymod = 0
+ epsrox = 3.9
+ pags = 1.7531187e-13
+ ntox = 1.0
+ pcit = -1.1898337e-16
+ pclm = 1.5094578
+ rdsmod = 0
+ ptvfbsdoff = 0
+ igbmod = 1
+ phin = 0.15
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ pbswgd = 0.95
+ pkt1 = -2.7321875e-14
+ pkt2 = -4.4253241e-16
+ pbswgs = 0.95
+ igcmod = 1
+ wpdiblc2 = 5.7318301e-9
+ pvoff = -2.4099793e-15
+ cdscb = 0
+ cdscd = 0
+ rbdb = 50
+ pua1 = 1.9942546e-22
+ prwb = 0
+ prwg = 0
+ pub1 = -1.9971615000000003e-31
+ puc1 = 1.7835157e-23
+ nfactor = 1
+ pvsat = -2.24e-11
+ rbpb = 50
+ rbpd = 50
+ wk2we = 5e-12
+ rbps = 50
+ pvth0 = 3.0076502e-15
+ rbsb = 50
+ pvag = 1.2
+ drout = 0.56
+ rdsw = 100
+ paigc = -1.0556924e-17
+ voffl = 0
+ paigsd = 1.1026372e-22
+ weta0 = -1.1162667e-8
+ wetab = 2.2325333e-8
+ wkvth0we = 2e-12
+ nigbacc = 10
+ permod = 1
+ trnqsmod = 0
+ cgidl = 0.22
+ rshg = 15.6
+ nigbinv = 10
+ pbswd = 0.8
+ pbsws = 0.8
+ voffcv = -0.16942
+ wpemod = 1
+ rgatemod = 0
+ tnjtsswg = 1
+ tnom = 25
+ pdits = 0
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ a0 = 3.8452644
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ cigsd = 0.069865
+ b1 = 0
+ at = -81312.781
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.020123392
+ k3 = -1.8419
+ em = 1000000.0
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ ll = 0
+ lw = 0
+ u0 = 0.01764456
+ w0 = 0
+ fnoimod = 1
+ ua = -1.6436128e-9
+ ub = 2.0158412e-18
+ uc = 5.8736458e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ eigbinv = 1.1
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ tpbswg = 0.0009
+ wags = -9.296980400000001e-8
+ wcit = 3.4826906000000003e-10
+ tnoia = 0
+ voff = -0.13348839
+ peta0 = 0.0
+ acde = 0.4
+ wketa = 1.8850903e-8
+ vsat = 102889.02
+ ptvoff = 2.7553621e-16
+ wint = 0
+ tpbsw = 0.0019
+ vth0 = 0.33129778
+ cigbacc = 0.32875
+ waigsd = 3.1111904e-12
+ wkt1 = 3.883104999999996e-10
+ wkt2 = -5.2803902e-9
+ cjswd = 7.7408e-11
+ cjsws = 7.7408e-11
+ wmax = 5.374e-7
+ mjswd = 0.11
+ aigc = 0.011795195
+ mjsws = 0.11
+ wmin = 2.674e-7
+ agidl = 9.41e-8
+ diomod = 1
+ tnoimod = 0
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 2.66208e-10
+ pku0we = -1.5e-18
+ wua1 = -2.0961923e-16
+ wub1 = 1.3682244e-25
+ cjswgs = 2.66208e-10
+ wuc1 = -2.9511024e-17
+ cigbinv = 0.006
+ bigc = 0.001442
+ wwlc = 0
+ tvfbsdoff = 0.022
+ cdsc = 0
+ mjswgd = 0.85
+ mjswgs = 0.85
+ scref = 1e-6
+ version = 4.5
+ ijthsfwd = 0.01
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ pigcd = 2.621
+ cgsl = 3.31989e-12
+ tcjswg = 0.001
+ cgso = 4.90562e-11
+ tempmod = 0
+ aigsd = 0.010772818
+ cigc = 0.000625
+ ags = 0.9274157999999999
+ lvoff = -1.1665524999999999e-8
+ cjd = 0.001281008
+ cit = 0.00026829437
+ cjs = 0.001281008
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ aigbacc = 0.02
+ dlc = 9.8024918e-9
+ lvsat = -0.0002
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ lvth0 = 5.0828999e-8
+ ijthsrev = 0.01
+ delta = 0.007595625
+ laigc = -1.416882e-10
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ la0 = -2.722152e-6
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ rnoia = 0
+ rnoib = 0
+ dmdg = 0
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = 0.20183035000000002
+ kt1 = -0.22156452
+ lk2 = -1.3986155e-8
+ kt2 = -0.033027229
+ llc = 0
+ lln = 1
+ lu0 = -2.2689026e-9
+ mjd = 0.26
+ aigbinv = 0.0163
+ lua = -2.9346741e-16
+ mjs = 0.26
+ lub = 5.7165214e-26
+ luc = 2.4824263e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 3.4236885e-13
+ fprout = 300
+ nsd = 1e+20
+ pbd = 0.52
+ pat = -6.371872400000001e-8
+ pbs = 0.52
+ pketa = -2.2733801e-14
+ pk2 = -1.3939214e-15
+ ngate = 8e+20
+ pu0 = 1.6723558e-16
+ xrcrg1 = 12
+ xrcrg2 = 1
+ k2we = 5e-5
+ prt = 0
+ pua = 4.226297e-23
+ pub = -4.4156209e-32
+ puc = -1.0695581e-23
+ pud = 0
+ ngcon = 1
+ wpclm = 9.3989653e-8
+ dsub = 0.75
+ rsh = 17.5
+ tcj = 0.00076
+ dtox = 2.7e-10
+ ua1 = 1.720591e-9
+ ub1 = -9.5473708e-19
+ uc1 = 7.0015137e-11
+ ppdiblc2 = -6.6555967e-15
+ tpb = 0.0014
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ wa0 = -4.9804098e-8
+ gbmin = 1e-12
+ ute = -1
+ wat = 0.078525419
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 2.0146831e-9
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ wtvoff = -3.0649189e-11
+ wlc = 0
+ wln = 1
+ wu0 = -1.3381044000000001e-9
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -1.3568102e-16
+ wub = 1.003525e-25
+ wuc = -1.2660669e-18
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ eta0 = 0.24044444
+ etab = -0.28088889
+ )

.model nch_fs_27 nmos (
+ level = 54
+ ntox = 1.0
+ pcit = -1.2805802e-16
+ pclm = 1.5094578
+ fnoimod = 1
+ phin = 0.15
+ eigbinv = 1.1
+ pbswd = 0.8
+ pbsws = 0.8
+ pkt1 = 4.8688443000000005e-15
+ pkt2 = 2.2738921e-15
+ pdits = 0
+ rbdb = 50
+ pua1 = -2.6369043e-23
+ prwb = 0
+ prwg = 0
+ pub1 = 4.8439292000000003e-32
+ cigsd = 0.069865
+ puc1 = 6.8677984e-24
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ dvt0w = 0
+ pvag = 1.2
+ dvt1w = 0
+ dvt2w = 0
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ rdsw = 100
+ ijthsfwd = 0.01
+ cigbacc = 0.32875
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ tnoimod = 0
+ tnoia = 0
+ ijthsrev = 0.01
+ cigbinv = 0.006
+ peta0 = 0.0
+ rshg = 15.6
+ wketa = -2.2122195e-8
+ wtvfbsdoff = 0
+ tpbsw = 0.0019
+ toxref = 3e-9
+ cjswd = 7.7408e-11
+ cjsws = 7.7408e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ version = 4.5
+ ltvfbsdoff = 0
+ tempmod = 0
+ ppdiblc2 = 1.7501102e-15
+ tnom = 25
+ aigbacc = 0.02
+ tvfbsdoff = 0.022
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ ltvoff = 1.3913801e-9
+ ags = 0.25766657
+ scref = 1e-6
+ cjd = 0.001281008
+ cit = 0.00059502911
+ cjs = 0.001281008
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 9.8024918e-9
+ pigcd = 2.621
+ k3b = 1.9326
+ aigsd = 0.010772818
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ ptvfbsdoff = 0
+ aigbinv = 0.0163
+ lvoff = -5.173220300000001e-10
+ wags = 3.7684035999999996e-7
+ lku0we = 2.5e-11
+ pkvth0we = -1.3e-19
+ la0 = 3.6355951e-7
+ epsrox = 3.9
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.052898453
+ kt1 = -0.19312528
+ lk2 = -1.4722356e-8
+ kt2 = -0.039065148
+ wcit = 3.584653e-10
+ lvsat = -0.0002
+ llc = 0
+ lln = 1
+ lu0 = -1.7420993e-9
+ mjd = 0.26
+ lvth0 = -8.6958156e-9
+ lua = -1.1159069e-16
+ mjs = 0.26
+ lub = -2.3732546e-26
+ luc = -2.9405776e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ voff = -0.14601446
+ njs = 1.02
+ pa0 = -3.8856002e-13
+ nsd = 1e+20
+ delta = 0.007595625
+ acde = 0.4
+ pbd = 0.52
+ wvfbsdoff = 0
+ pat = -8.840236300000001e-10
+ pbs = 0.52
+ rdsmod = 0
+ pk2 = 1.1847359e-15
+ lvfbsdoff = 0
+ laigc = -3.3762752e-11
+ pu0 = 1.3152191e-16
+ vfbsdoff = 0.02
+ igbmod = 1
+ prt = 0
+ pua = 2.9945529e-23
+ pub = -3.9782718e-32
+ puc = 6.3626704e-24
+ pud = 0
+ vsat = 102889.02
+ wint = 0
+ rnoia = 0
+ rnoib = 0
+ vth0 = 0.39817958999999997
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 6.6639379e-10
+ ub1 = 1.1665789e-19
+ uc1 = 5.9635906e-11
+ wkt1 = -3.5781036999999996e-8
+ wkt2 = -8.3325526e-9
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ tpb = 0.0014
+ wmax = 5.374e-7
+ wa0 = 7.714643e-7
+ aigc = 0.01167393
+ wmin = 2.674e-7
+ ute = -1
+ wat = 0.0079246317
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -8.8268726e-10
+ pbswgd = 0.95
+ pketa = 1.3732256e-14
+ poxedge = 1
+ pbswgs = 0.95
+ ngate = 8e+20
+ wlc = 0
+ wln = 1
+ wu0 = -1.2979767e-9
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -1.218412e-16
+ wub = 9.5438468e-26
+ wuc = -2.0432641e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ ngcon = 1
+ paramchk = 1
+ wpclm = 9.3989653e-8
+ igcmod = 1
+ binunit = 2
+ wua1 = 4.4082452e-17
+ wub1 = -1.420039e-25
+ wuc1 = -1.718815e-17
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ bigc = 0.001442
+ wwlc = 0
+ cdsc = 0
+ ijthdfwd = 0.01
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ permod = 1
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ ijthdrev = 0.01
+ tvoff = -0.0014023534
+ lpdiblc2 = -7.3119259e-9
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ voffcv = -0.16942
+ wpemod = 1
+ k2we = 5e-5
+ ku0we = -0.0007
+ dsub = 0.75
+ dtox = 2.7e-10
+ beta0 = 13
+ leta0 = 1.6000000000000003e-9
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ njtsswg = 9
+ lkvth0we = -2e-12
+ eta0 = 0.24044444
+ etab = -0.28088889
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.039504569
+ pdiblcb = -0.3
+ tpbswg = 0.0009
+ acnqsmod = 0
+ dmcgt = 0
+ tcjsw = 0.000357
+ rbodymod = 0
+ ptvoff = -5.8159511e-16
+ bigbacc = 0.002588
+ waigsd = 3.1113143e-12
+ bigsd = 0.00125
+ a0 = 0.37817284
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 204899.36
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.020950589999999998
+ k3 = -1.8419
+ em = 1000000.0
+ kvth0we = 0.00018
+ diomod = 1
+ ll = 0
+ lw = 0
+ u0 = 0.017052646
+ w0 = 0
+ wvoff = 1.6411259e-8
+ ua = -1.8479686e-9
+ ub = 2.1067376e-18
+ uc = 1.1966909e-10
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ lintnoi = -1.5e-8
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 2.66208e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.66208e-10
+ bigbinv = 0.004953
+ wvsat = -0.0028059037
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ wvth0 = -2.4499761e-8
+ wpdiblc2 = -3.7127843e-9
+ waigc = 2.313153e-11
+ mjswgd = 0.85
+ mjswgs = 0.85
+ lketa = -4.8021757e-8
+ tcjswg = 0.001
+ xpart = 1
+ pvfbsdoff = 0
+ keta = 0.03621471
+ egidl = 0.29734
+ wkvth0we = 2e-12
+ lags = 4.1799271e-7
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 3.6898897e-10
+ trnqsmod = 0
+ kt1l = 0
+ nfactor = 1
+ lint = 6.5375218e-9
+ fprout = 300
+ lkt1 = -1.6733642999999998e-8
+ lkt2 = -1.6288295e-8
+ xrcrg1 = 12
+ xrcrg2 = 1
+ lmax = 8.9908e-7
+ lmin = 4.4908e-7
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ rgatemod = 0
+ wtvoff = 9.3241971e-10
+ pvoff = -4.5972513e-15
+ minv = -0.3
+ tnjtsswg = 1
+ lua1 = 4.5439491e-17
+ lub1 = -2.7049927e-25
+ luc1 = 3.3118724e-18
+ cdscb = 0
+ cdscd = 0
+ nigbacc = 10
+ ndep = 1e+18
+ pvsat = -2.24e-11
+ wk2we = 5e-12
+ pvth0 = 5.8409157999999994e-15
+ lwlc = 0
+ drout = 0.56
+ moin = 5.1
+ capmod = 2
+ paigc = -4.5341069e-18
+ nigc = 3.083
+ voffl = 0
+ wku0we = 2e-11
+ nigbinv = 10
+ mobmod = 0
+ weta0 = -1.1162667e-8
+ wetab = 2.2325333e-8
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ pags = -2.4281917e-13
+ cgidl = 0.22
+ )

.model nch_fs_28 nmos (
+ level = 54
+ wuc1 = -1.3268706e-17
+ bigc = 0.001442
+ ppclm = -7.9196439e-14
+ wwlc = 0
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ cdsc = 0
+ bigbacc = 0.002588
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ wtvfbsdoff = 0
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ kvth0we = 0.00018
+ dmcgt = 0
+ tcjsw = 0.000357
+ wkvth0we = 2e-12
+ lintnoi = -1.5e-8
+ ltvfbsdoff = 0
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ trnqsmod = 0
+ toxref = 3e-9
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ bigsd = 0.00125
+ wvoff = 5.1767953e-9
+ k2we = 5e-5
+ dsub = 0.75
+ wvsat = -0.0054199005
+ dtox = 2.7e-10
+ ptvfbsdoff = 0
+ wvth0 = -6.886954300000001e-9
+ rgatemod = 0
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ tnjtsswg = 1
+ waigc = -1.6608588e-12
+ ltvoff = -7.6859018e-11
+ eta0 = 0.24044444
+ etab = -0.28088889
+ lketa = -5.7215427e-9
+ nfactor = 1
+ xpart = 1
+ pvfbsdoff = 0
+ lku0we = 2.5e-11
+ egidl = 0.29734
+ epsrox = 3.9
+ rdsmod = 0
+ igbmod = 1
+ nigbacc = 10
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ pbswgd = 0.95
+ pbswgs = 0.95
+ igcmod = 1
+ nigbinv = 10
+ pvoff = 3.4591262e-16
+ cdscb = 0
+ cdscd = 0
+ pvsat = 1.1277586e-9
+ wk2we = 5e-12
+ pvth0 = -1.9087192e-15
+ drout = 0.56
+ paigc = 6.374544e-18
+ ijthsfwd = 0.01
+ paigsd = 2.2627557e-23
+ voffl = 0
+ fnoimod = 1
+ eigbinv = 1.1
+ keta = -0.05992214
+ weta0 = -1.1162667e-8
+ wetab = 2.2325333e-8
+ permod = 1
+ lpclm = 1.4504842e-7
+ lags = 5.906061e-7
+ jswd = 1.28e-13
+ ijthsrev = 0.01
+ jsws = 1.28e-13
+ lcit = 8.536557100000001e-11
+ cgidl = 0.22
+ kt1l = 0
+ lint = 9.7879675e-9
+ voffcv = -0.16942
+ wpemod = 1
+ lkt1 = 8.3803069e-9
+ lkt2 = -2.5638367e-9
+ lmax = 4.4908e-7
+ cigbacc = 0.32875
+ pbswd = 0.8
+ pbsws = 0.8
+ lmin = 2.1577e-7
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ ppdiblc2 = -5.242001e-17
+ tnoimod = 0
+ minv = -0.3
+ lua1 = -4.6794128e-17
+ lub1 = -3.5289654e-26
+ luc1 = -2.1335001e-17
+ pdits = 0
+ ndep = 1e+18
+ cigsd = 0.069865
+ cigbinv = 0.006
+ dvt0w = 0
+ lwlc = 0
+ dvt1w = 0
+ dvt2w = 0
+ moin = 5.1
+ nigc = 3.083
+ tpbswg = 0.0009
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ version = 4.5
+ tempmod = 0
+ pkvth0we = -1.3e-19
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ tnoia = 0
+ pags = 1.2428184e-13
+ peta0 = 0.0
+ ptvoff = -1.5558646e-16
+ aigbacc = 0.02
+ ntox = 1.0
+ pcit = -2.09847229e-17
+ pclm = 1.1798023
+ waigsd = 3.1112628e-12
+ wketa = 2.3981389e-8
+ vfbsdoff = 0.02
+ tpbsw = 0.0019
+ cjswd = 7.7408e-11
+ cjsws = 7.7408e-11
+ diomod = 1
+ mjswd = 0.11
+ phin = 0.15
+ mjsws = 0.11
+ agidl = 9.41e-8
+ pditsd = 0
+ pditsl = 0
+ aigbinv = 0.0163
+ pkt1 = -1.2444052000000001e-14
+ pkt2 = -7.0784646e-16
+ cjswgd = 2.66208e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.66208e-10
+ paramchk = 1
+ ags = -0.134636584
+ cjd = 0.001281008
+ tvfbsdoff = 0.022
+ cit = 0.0012396277
+ cjs = 0.001281008
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 1.30529375e-8
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ rbdb = 50
+ pua1 = 1.8291934e-23
+ prwb = 0
+ prwg = 0
+ pub1 = -6.872418799999999e-33
+ puc1 = 5.143243e-24
+ mjswgd = 0.85
+ mjswgs = 0.85
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ tcjswg = 0.001
+ rdsw = 100
+ scref = 1e-6
+ ijthdfwd = 0.01
+ la0 = -6.0902319e-7
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.015196938
+ kt1 = -0.25020244
+ lk2 = -1.0681005e-8
+ kt2 = -0.070257098
+ pigcd = 2.621
+ llc = -1.18e-13
+ lln = 0.7
+ aigsd = 0.010772818
+ lu0 = -6.9623626e-10
+ mjd = 0.26
+ lua = -1.8564943e-17
+ mjs = 0.26
+ lub = -5.2748233e-26
+ luc = -4.2757753e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 2.2627554e-14
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 2.5333001000000004e-9
+ poxedge = 1
+ pbs = 0.52
+ pk2 = 8.6250113e-16
+ lvoff = -7.1634494e-9
+ a0 = 2.5885881
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ pu0 = 5.2978272000000005e-17
+ at = 119214.09
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.011765692
+ k3 = -1.8419
+ em = 1000000.0
+ prt = 0
+ pua = 5.6394132e-24
+ pub = -7.710339e-34
+ puc = -1.5613012e-24
+ pud = 0
+ ll = -1.18e-13
+ lw = 0
+ u0 = 0.014675684
+ w0 = 0
+ ua = -2.0593908e-9
+ ub = 2.1726824e-18
+ uc = 6.2555449e-11
+ ud = 0
+ wl = 0
+ rsh = 17.5
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ tcj = 0.00076
+ ua1 = 8.7601565e-10
+ lvsat = -0.0043672412
+ ub1 = -4.1790941e-19
+ uc1 = 1.1565153e-10
+ binunit = 2
+ lvth0 = 9.94398e-10
+ ijthdrev = 0.01
+ tpb = 0.0014
+ wvfbsdoff = 0
+ wa0 = -1.6305293e-7
+ lvfbsdoff = 0
+ ute = -1
+ wat = 0.00015798693
+ delta = 0.007595625
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -1.5033038e-10
+ laigc = -3.7429738e-11
+ wlc = 0
+ wln = 1
+ rshg = 15.6
+ wu0 = -1.1194684000000002e-9
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -6.6600022e-17
+ wub = 6.7755498e-27
+ wuc = -2.4236148e-18
+ wud = 0
+ lpdiblc2 = -4.2799755e-9
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ rnoia = 0
+ rnoib = 0
+ fprout = 300
+ xrcrg1 = 12
+ xrcrg2 = 1
+ pketa = -6.5533207e-15
+ ngate = 8e+20
+ ngcon = 1
+ wpclm = 2.7398156e-7
+ wtvoff = -3.5781771e-11
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ tnom = 25
+ jswgs = 1.28e-13
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ lkvth0we = -2e-12
+ capmod = 2
+ wku0we = 2e-11
+ mobmod = 0
+ acnqsmod = 0
+ wags = -4.5748013000000004e-7
+ wcit = 1.1511689100000001e-10
+ rbodymod = 0
+ voff = -0.13090963
+ acde = 0.4
+ tvoff = 0.0019345538
+ njtsswg = 9
+ vsat = 112360.02
+ wint = 0
+ xjbvd = 1
+ xjbvs = 1
+ vth0 = 0.37615638
+ lk2we = -1.5e-12
+ wkt1 = 3.5664547999999997e-9
+ wkt2 = -1.5558741e-9
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ wmax = 5.374e-7
+ laigsd = -8.1983894e-17
+ aigc = 0.011682264
+ wmin = 2.674e-7
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.032613772
+ pdiblcb = -0.3
+ ku0we = -0.0007
+ beta0 = 13
+ leta0 = 1.6000000000000003e-9
+ wua1 = -5.7419768e-17
+ wpdiblc2 = 3.8387521e-10
+ wub1 = -1.6295463e-26
+ )

.model nch_fs_29 nmos (
+ level = 54
+ keta = 0.0092481698
+ aigbinv = 0.0163
+ tnoia = 0
+ ijthdrev = 0.01
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = -2.1537106e-11
+ peta0 = 0.0
+ ptvfbsdoff = 0
+ kt1l = 0
+ wketa = -2.0169501e-8
+ toxref = 3e-9
+ lpdiblc2 = -9.0824285e-10
+ tpbsw = 0.0019
+ ags = 2.6644444
+ cjswd = 7.7408e-11
+ cjsws = 7.7408e-11
+ lint = 9.7879675e-9
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ cjd = 0.001281008
+ cit = 0.0017462755
+ cjs = 0.001281008
+ clc = 1e-7
+ cle = 0.6
+ lkt1 = -3.0062126e-9
+ bvd = 8.7
+ lkt2 = -3.9513595e-9
+ bvs = 8.7
+ lmax = 2.1577e-7
+ dlc = 1.30529375e-8
+ lmin = 9e-8
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ poxedge = 1
+ tvfbsdoff = 0.022
+ la0 = -2.075695e-7
+ minv = -0.3
+ jsd = 6.11e-7
+ ltvoff = 5.8839234e-11
+ jss = 6.11e-7
+ lat = -0.0017537311
+ lua1 = -5.8912951e-18
+ lub1 = -3.1777439e-26
+ luc1 = 1.0640856e-17
+ kt1 = -0.1962379
+ lk2 = -3.2022951e-9
+ kt2 = -0.063681161
+ llc = -1.18e-13
+ binunit = 2
+ lln = 0.7
+ lu0 = -2.4591767000000003e-10
+ mjd = 0.26
+ lua = 5.2959027e-17
+ mjs = 0.26
+ lub = -7.97606935e-26
+ luc = -8.8267893e-18
+ lud = 0
+ lwc = 0
+ ndep = 1e+18
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ lkvth0we = -2e-12
+ njs = 1.02
+ pa0 = 1.0407708e-13
+ nsd = 1e+20
+ lwlc = 0
+ pbd = 0.52
+ pat = -4.0201951e-10
+ pbs = 0.52
+ pk2 = -9.7578421e-17
+ moin = 5.1
+ pu0 = 2.0100797e-17
+ prt = 0
+ pua = -7.1102082e-24
+ pub = 9.57267e-33
+ puc = 7.19078e-25
+ pud = 0
+ scref = 1e-6
+ nigc = 3.083
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 6.8216336e-10
+ pigcd = 2.621
+ ub1 = -4.3455498e-19
+ uc1 = -3.5892821e-11
+ aigsd = 0.010772818
+ tpb = 0.0014
+ lku0we = 2.5e-11
+ wa0 = -5.4906963e-7
+ acnqsmod = 0
+ ute = -1
+ wat = 0.014069454
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 4.3998097e-9
+ epsrox = 3.9
+ lvoff = 2.31636653e-9
+ wlc = 0
+ wln = 1
+ wu0 = -9.6365099e-10
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -6.1752756e-18
+ wub = -4.2246744000000004e-26
+ wuc = -1.3231099e-17
+ wud = 0
+ wwc = 0
+ noff = 2.7195
+ wwl = 0
+ wwn = 1
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ lvsat = -0.0006573482700000001
+ rbodymod = 0
+ rdsmod = 0
+ wvfbsdoff = 0
+ lvth0 = -1.26749906e-8
+ lvfbsdoff = 0
+ igbmod = 1
+ delta = 0.007595625
+ laigc = 2.6175146e-12
+ ntox = 1.0
+ pcit = -4.179175200000001e-18
+ jtsswgd = 2.3e-7
+ pclm = 2.3689724
+ jtsswgs = 2.3e-7
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ rnoia = 0
+ rnoib = 0
+ pbswgd = 0.95
+ pbswgs = 0.95
+ phin = 0.15
+ pketa = 2.762517e-15
+ ngate = 8e+20
+ igcmod = 1
+ ngcon = 1
+ pkt1 = 7.2116645e-16
+ pkt2 = 9.3582987e-16
+ wpclm = -2.0834879e-7
+ wpdiblc2 = 1.3111248e-10
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ rbdb = 50
+ pua1 = 1.9734917e-24
+ prwb = 0
+ prwg = 0
+ pub1 = -5.5422001e-33
+ puc1 = -4.0873907e-24
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ njtsswg = 9
+ paigsd = -9.4615512e-24
+ rdsw = 100
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ permod = 1
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.016633997
+ pdiblcb = -0.3
+ wkvth0we = 2e-12
+ trnqsmod = 0
+ tvoff = 0.0012914341
+ rshg = 15.6
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ voffcv = -0.16942
+ wpemod = 1
+ bigbacc = 0.002588
+ ku0we = -0.0007
+ kvth0we = 0.00018
+ beta0 = 13
+ leta0 = 1.6000000000000003e-9
+ rgatemod = 0
+ lintnoi = -1.5e-8
+ tnjtsswg = 1
+ tnom = 25
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ ppclm = 2.2575265e-14
+ vtsswgs = 4.2
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ tpbswg = 0.0009
+ dmcgt = 0
+ wags = 1.3153333e-7
+ tcjsw = 0.000357
+ wcit = 3.5469746200000003e-11
+ ptvoff = 2.7225835e-17
+ voff = -0.175837897
+ waigsd = 3.1114149e-12
+ acde = 0.4
+ vsat = 94777.65030000001
+ wint = 0
+ bigsd = 0.00125
+ vth0 = 0.440940454
+ diomod = 1
+ wkt1 = -5.8827946e-8
+ wkt2 = -9.3458092e-9
+ wmax = 5.374e-7
+ aigc = 0.011492467
+ wmin = 2.674e-7
+ nfactor = 1
+ pditsd = 0
+ pditsl = 0
+ wvoff = 8.989216699999998e-9
+ cjswgd = 2.66208e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.66208e-10
+ wvsat = -0.0005775380999999999
+ wvth0 = -2.0325728e-8
+ wua1 = 1.991882e-17
+ wub1 = -2.2599817e-26
+ wuc1 = 3.0478373e-17
+ waigc = 3.9031408e-11
+ bigc = 0.001442
+ mjswgd = 0.85
+ mjswgs = 0.85
+ wwlc = 0
+ tcjswg = 0.001
+ nigbacc = 10
+ lketa = -2.0316478e-8
+ cdsc = 0
+ ijthsfwd = 0.01
+ cgbo = 0
+ xpart = 1
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ pvfbsdoff = 0
+ xtid = 3
+ xtis = 3
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ egidl = 0.29734
+ nigbinv = 10
+ ijthsrev = 0.01
+ fprout = 300
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ fnoimod = 1
+ k2we = 5e-5
+ wtvoff = -9.0219076e-10
+ eigbinv = 1.1
+ dsub = 0.75
+ dtox = 2.7e-10
+ ppdiblc2 = 9.1292629e-19
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ pvoff = -4.585090499999998e-16
+ a0 = 0.68596391
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 55502.213
+ cf = 8.15e-11
+ cdscb = 0
+ cdscd = 0
+ ef = 1.0
+ k1 = 0.274
+ k2 = -0.02367843
+ k3 = -1.8419
+ em = 1000000.0
+ ll = -1.18e-13
+ lw = 0
+ u0 = 0.012541473
+ pvsat = 1.0602156000000003e-10
+ w0 = 0
+ ua = -2.398367e-9
+ ub = 2.300703286e-18
+ uc = 8.4124236e-11
+ ud = 0
+ wk2we = 5e-12
+ capmod = 2
+ wl = 0
+ wr = 1
+ pvth0 = 9.268619999999999e-16
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ eta0 = 0.24044444
+ xw = 8.600000000000001e-9
+ drout = 0.56
+ etab = -0.28088889
+ wku0we = 2e-11
+ paigc = -2.2115244e-18
+ mobmod = 0
+ voffl = 0
+ cigbacc = 0.32875
+ weta0 = -1.1162667e-8
+ wetab = 2.2325333e-8
+ pkvth0we = -1.3e-19
+ lpclm = -1.0586647e-7
+ tnoimod = 0
+ cgidl = 0.22
+ vfbsdoff = 0.02
+ cigbinv = 0.006
+ laigsd = 3.4280989e-17
+ pbswd = 0.8
+ pbsws = 0.8
+ paramchk = 1
+ version = 4.5
+ wtvfbsdoff = 0
+ tempmod = 0
+ pdits = 0
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ cigsd = 0.069865
+ ltvfbsdoff = 0
+ dvt0w = 0
+ aigbacc = 0.02
+ dvt1w = 0
+ dvt2w = 0
+ ijthdfwd = 0.01
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ )

.model nch_fs_30 nmos (
+ level = 54
+ keta = -0.29566775
+ aigbinv = 0.0163
+ tnoia = 0
+ ijthdrev = 0.01
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 1.6634428e-10
+ peta0 = -9.3037135e-16
+ ptvfbsdoff = 0
+ petab = -1.2138265e-15
+ kt1l = 0
+ wketa = -4.7865407e-8
+ toxref = 3e-9
+ lpdiblc2 = 8.2379047e-15
+ tpbsw = 0.0019
+ ags = 2.6644444
+ cjswd = 7.7408e-11
+ cjsws = 7.7408e-11
+ lint = 0
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ cjd = 0.001281008
+ cit = -0.00025246267
+ cjs = 0.001281008
+ clc = 1e-7
+ cle = 0.6
+ lkt1 = -8.9750836e-9
+ bvd = 8.7
+ lkt2 = 3.8424987e-10
+ bvs = 8.7
+ lmax = 9e-8
+ dlc = 3.26497e-9
+ lmin = 5.4e-8
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ poxedge = 1
+ tvfbsdoff = 0.022
+ la0 = 3.9829889e-7
+ minv = -0.3
+ jsd = 6.11e-7
+ ltvoff = -2.7237524e-10
+ jss = 6.11e-7
+ lat = 0.005125604979999999
+ lua1 = -1.2736334e-17
+ lub1 = 1.3685594e-26
+ luc1 = 1.132730421e-17
+ kt1 = -0.13273927
+ lk2 = 1.0502722e-9
+ kt2 = -0.10980467
+ llc = 0
+ binunit = 2
+ lln = 1
+ lu0 = -1.9515966e-10
+ mjd = 0.26
+ lua = -7.6887484e-18
+ mjs = 0.26
+ lub = 6.3606825e-27
+ luc = -3.2720592999999998e-18
+ lud = 0
+ lwc = 0
+ ndep = 1e+18
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ lkvth0we = -2e-12
+ njs = 1.02
+ pa0 = -1.1411036e-13
+ nsd = 1e+20
+ lwlc = 0
+ pbd = 0.52
+ pat = -1.7624563e-9
+ pbs = 0.52
+ pk2 = -3.7289588e-16
+ moin = 5.1
+ pu0 = 7.4424501e-17
+ prt = 0
+ pua = 1.3044266e-23
+ pub = -1.13966382e-32
+ puc = 2.3653651e-24
+ pud = 0
+ scref = 1e-6
+ nigc = 3.083
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 7.5498293e-10
+ pigcd = 2.621
+ ub1 = -9.1820427e-19
+ uc1 = -4.319545900000001e-11
+ aigsd = 0.010772818
+ tpb = 0.0014
+ lku0we = 2.5e-11
+ wa0 = 1.7720733e-6
+ acnqsmod = 0
+ ute = -1
+ wat = 0.028542186400000003
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 7.3287188e-9
+ epsrox = 3.9
+ lvoff = -3.2671799e-9
+ wlc = 0
+ wln = 1
+ wu0 = -1.5415627e-9
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -2.2058458e-16
+ wub = 1.80830997e-25
+ wuc = -3.0744792e-17
+ wud = 0
+ wwc = 0
+ noff = 2.7195
+ wwl = 0
+ wwn = 1
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ lvsat = 0.0027394203000000008
+ rbodymod = 0
+ rdsmod = 0
+ wvfbsdoff = 0
+ lvth0 = 3.109724299999999e-9
+ lvfbsdoff = 0
+ igbmod = 1
+ delta = 0.007595625
+ laigc = -3.0244582e-11
+ ntox = 1.0
+ pcit = -3.1457676000000004e-17
+ jtsswgd = 2.3e-7
+ pclm = 1.7776553
+ jtsswgs = 2.3e-7
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ rnoia = 0
+ rnoib = 0
+ pbswgd = 0.95
+ pbswgs = 0.95
+ phin = 0.15
+ pketa = 5.3659323e-15
+ ngate = 8e+20
+ igcmod = 1
+ ngcon = 1
+ pkt1 = 5.1625068e-15
+ pkt2 = -5.9202052e-16
+ wpclm = 4.3365813e-8
+ wpdiblc2 = 1.4083642e-10
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ rbdb = 50
+ pua1 = 4.1884121e-24
+ prwb = 0
+ prwg = 0
+ pub1 = -1.01069988e-32
+ puc1 = -6.8508479999999965e-25
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ njtsswg = 9
+ rdsw = 100
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ permod = 1
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.0069717513
+ pdiblcb = -0.3
+ wkvth0we = 2e-12
+ trnqsmod = 0
+ tvoff = 0.0048149924
+ rshg = 15.6
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ voffcv = -0.16942
+ wpemod = 1
+ bigbacc = 0.002588
+ ku0we = -0.0007
+ kvth0we = 0.00018
+ beta0 = 13
+ leta0 = 2.1640249e-8
+ rgatemod = 0
+ letab = -2.6551319e-8
+ lintnoi = -1.5e-8
+ tnjtsswg = 1
+ tnom = 25
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ ppclm = -1.085908e-15
+ vtsswgs = 4.2
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ tpbswg = 0.0009
+ dmcgt = 0
+ wags = 1.3153333e-7
+ tcjsw = 0.000357
+ wcit = 3.2566656e-10
+ ptvoff = 9.0058483e-17
+ voff = -0.116438471
+ waigsd = 3.1113143e-12
+ acde = 0.4
+ vsat = 58641.813
+ wint = 0
+ bigsd = 0.00125
+ vth0 = 0.273017953
+ diomod = 1
+ wkt1 = -1.0607625000000001e-7
+ wkt2 = 6.9079183e-9
+ wmax = 5.374e-7
+ aigc = 0.011842064
+ wmin = 2.674e-7
+ nfactor = 1
+ pditsd = 0
+ pditsl = 0
+ wvoff = 4.307686799999997e-9
+ cjswgd = 2.66208e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.66208e-10
+ wvsat = 0.0042232395
+ wvth0 = -9.925777100000002e-9
+ wua1 = -3.6441631e-18
+ wub1 = 2.5961869999999995e-26
+ wuc1 = -5.7163699999999976e-18
+ waigc = 4.5087747e-12
+ bigc = 0.001442
+ mjswgd = 0.85
+ mjswgs = 0.85
+ wwlc = 0
+ tcjswg = 0.001
+ nigbacc = 10
+ lketa = 8.345618e-9
+ cdsc = 0
+ ijthsfwd = 0.01
+ cgbo = 0
+ xpart = 1
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ pvfbsdoff = 0
+ xtid = 3
+ xtis = 3
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ egidl = 0.29734
+ nigbinv = 10
+ ijthsrev = 0.01
+ fprout = 300
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ fnoimod = 1
+ k2we = 5e-5
+ wtvoff = -1.5706231e-9
+ eigbinv = 1.1
+ dsub = 0.75
+ dtox = 2.7e-10
+ ppdiblc2 = -1.1241984e-21
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ pvoff = -1.8445117999999986e-17
+ a0 = -5.7594444
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = -17682.2125
+ cf = 8.15e-11
+ cdscb = 0
+ cdscd = 0
+ ef = 1.0
+ k1 = 0.274
+ k2 = -0.068918509
+ k3 = -1.8419
+ em = 1000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.012001494
+ pvsat = -3.452516000000002e-10
+ w0 = 0
+ ua = -1.7531779e-9
+ ub = 1.3845184050000002e-18
+ uc = 2.5031363e-11
+ ud = 0
+ wk2we = 5e-12
+ capmod = 2
+ wl = 0
+ wr = 1
+ pvth0 = -5.073333999999973e-17
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ eta0 = 0.027250304
+ xw = 8.600000000000001e-9
+ drout = 0.56
+ etab = 0.001571952
+ wku0we = 2e-11
+ paigc = 1.0336032e-18
+ mobmod = 0
+ voffl = 0
+ cigbacc = 0.32875
+ weta0 = -1.2650991e-9
+ wetab = 3.5238381e-8
+ pkvth0we = -1.3e-19
+ lpclm = -5.0282662e-8
+ tnoimod = 0
+ cgidl = 0.22
+ vfbsdoff = 0.02
+ cigbinv = 0.006
+ pbswd = 0.8
+ pbsws = 0.8
+ paramchk = 1
+ version = 4.5
+ wtvfbsdoff = 0
+ tempmod = 0
+ pdits = 0
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ cigsd = 0.069865
+ ltvfbsdoff = 0
+ dvt0w = 0
+ aigbacc = 0.02
+ dvt1w = 0
+ dvt2w = 0
+ ijthdfwd = 0.01
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ )

.model nch_fs_31 nmos (
+ level = 54
+ nigbacc = 10
+ wvoff = 2.6164685300000083e-9
+ wvsat = 0.0269709042
+ wvth0 = -3.3487313000000005e-8
+ ltvoff = 2.6647905e-10
+ waigc = 1.8753243e-11
+ tnom = 25
+ nigbinv = 10
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ lketa = -2.3617222e-8
+ pvfbsdoff = 0
+ xpart = 1
+ lku0we = 2.5e-11
+ epsrox = 3.9
+ egidl = 0.29734
+ fnoimod = 1
+ pkvth0we = -1.3e-19
+ wags = 1.3153333e-7
+ rdsmod = 0
+ eigbinv = 1.1
+ wcit = 4.1128934000000004e-10
+ igbmod = 1
+ voff = -0.07382279000000001
+ acde = 0.4
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ vfbsdoff = 0.02
+ vsat = 22700.879999999997
+ pbswgd = 0.95
+ pbswgs = 0.95
+ wint = 0
+ vth0 = 0.29242439000000003
+ wkt1 = -1.9254349e-8
+ wkt2 = -2.0876247e-8
+ wmax = 5.374e-7
+ igcmod = 1
+ aigc = 0.011696193
+ wmin = 2.674e-7
+ paramchk = 1
+ cigbacc = 0.32875
+ wua1 = -1.1132499e-16
+ wub1 = 7.746802000000003e-26
+ wuc1 = 1.6593491000000002e-16
+ pvoff = 7.964544000000045e-17
+ bigc = 0.001442
+ cdscb = 0
+ cdscd = 0
+ tnoimod = 0
+ wwlc = 0
+ pvsat = -1.6646160000000002e-9
+ wk2we = 5e-12
+ pvth0 = 1.3158357999999997e-15
+ drout = 0.56
+ paigsd = 1.7624612e-23
+ cdsc = 0
+ paigc = 2.0742404e-19
+ cigbinv = 0.006
+ ijthdfwd = 0.01
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ voffl = 0
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ permod = 1
+ weta0 = -1.2005104e-7
+ wetab = 5.6750807e-8
+ lpclm = 5.458214e-8
+ version = 4.5
+ tempmod = 0
+ ijthdrev = 0.01
+ cgidl = 0.22
+ voffcv = -0.16942
+ wpemod = 1
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ aigbacc = 0.02
+ pbswd = 0.8
+ pbsws = 0.8
+ k2we = 5e-5
+ dsub = 0.75
+ dtox = 2.7e-10
+ aigbinv = 0.0163
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ pdits = 0
+ cigsd = 0.069865
+ lkvth0we = -2e-12
+ eta0 = 1.0176617
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ etab = -1.3959412
+ tpbswg = 0.0009
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ acnqsmod = 0
+ tnoia = 0
+ ptvoff = -4.401556e-18
+ poxedge = 1
+ rbodymod = 0
+ ags = 2.6644444
+ waigsd = 3.1110104e-12
+ peta0 = 5.9592132e-15
+ cjd = 0.001281008
+ cit = -0.0053709179
+ cjs = 0.001281008
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ petab = -2.4615472e-15
+ dlc = 3.26497e-9
+ binunit = 2
+ wketa = -5.877032e-8
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ diomod = 1
+ tpbsw = 0.0019
+ cjswd = 7.7408e-11
+ cjsws = 7.7408e-11
+ mjswd = 0.11
+ pditsd = 0
+ pditsl = 0
+ mjsws = 0.11
+ agidl = 9.41e-8
+ cjswgd = 2.66208e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.66208e-10
+ la0 = -1.4097724e-8
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.0008794376999999999
+ kt1 = -0.39757001
+ lk2 = 7.4338958e-10
+ kt2 = -0.14677127
+ llc = 0
+ lln = 1
+ lu0 = 5.173005800000001e-10
+ mjd = 0.26
+ lua = 6.4763643e-17
+ mjs = 0.26
+ lub = -2.3096342000000002e-26
+ luc = -1.0931136000000001e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = -1.7333804e-13
+ nsd = 1e+20
+ pbd = 0.52
+ pat = -4.6829471e-10
+ tvfbsdoff = 0.022
+ pbs = 0.52
+ pk2 = -1.0803308e-16
+ wpdiblc2 = 1.4081704e-10
+ pu0 = -4.4287482999999995e-17
+ prt = 0
+ pua = -2.1774501e-24
+ pub = -5.473259300000002e-33
+ puc = 4.761497700000001e-24
+ pud = 0
+ mjswgd = 0.85
+ mjswgs = 0.85
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 1.4910078e-9
+ ub1 = -1.7286540799999999e-18
+ uc1 = -4.0168785999999996e-10
+ tpb = 0.0014
+ tcjswg = 0.001
+ wa0 = 2.7932403e-6
+ ute = -1
+ wat = 0.006229054600000004
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 2.7621189e-9
+ wlc = 0
+ wln = 1
+ wu0 = 5.051956e-10
+ jtsswgd = 2.3e-7
+ xgl = -1.09e-8
+ jtsswgs = 2.3e-7
+ xgw = 0
+ wua = 4.1858808e-17
+ wub = 7.870378029999999e-26
+ wuc = -7.2057435e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ scref = 1e-6
+ pigcd = 2.621
+ aigsd = 0.010772819
+ keta = 0.2554158
+ lvoff = -5.7388898000000006e-9
+ wkvth0we = 2e-12
+ wvfbsdoff = 0
+ lvsat = 0.00482399457
+ lvfbsdoff = 0
+ lvth0 = 1.9841506000000015e-9
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 4.6321468999999995e-10
+ trnqsmod = 0
+ delta = 0.007595625
+ laigc = -2.1784105e-11
+ kt1l = 0
+ fprout = 300
+ xrcrg1 = 12
+ xrcrg2 = 1
+ rnoia = 0
+ rnoib = 0
+ lint = 0
+ njtsswg = 9
+ lkt1 = 6.3850994e-9
+ lkt2 = 2.528313e-9
+ pketa = 5.998417e-15
+ ngate = 8e+20
+ lmax = 5.4e-8
+ lmin = 4.5e-8
+ wtvoff = 5.799816e-11
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ ngcon = 1
+ wpclm = 2.4669208e-7
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ ckappad = 0.6
+ ckappas = 0.6
+ rgatemod = 0
+ gbmin = 1e-12
+ pdiblc1 = 0
+ pdiblc2 = 0.0069718933
+ pdiblcb = -0.3
+ tnjtsswg = 1
+ minv = -0.3
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ lua1 = -5.5425775e-17
+ lub1 = 6.069167999999999e-26
+ luc1 = 3.2119863e-17
+ capmod = 2
+ ndep = 1e+18
+ wku0we = 2e-11
+ lwlc = 0
+ moin = 5.1
+ mobmod = 0
+ nigc = 3.083
+ bigbacc = 0.002588
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ kvth0we = 0.00018
+ wtvfbsdoff = 0
+ lintnoi = -1.5e-8
+ bigbinv = 0.004953
+ tvoff = -0.0044755986
+ ntox = 1.0
+ vtsswgd = 4.2
+ pcit = -3.6423797000000005e-17
+ vtsswgs = 4.2
+ pclm = -0.030358553
+ laigsd = -6.385731e-17
+ xjbvd = 1
+ a0 = 1.350842
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ xjbvs = 1
+ lk2we = -1.5e-12
+ at = 85853.00300000001
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = -0.063627428
+ k3 = -1.8419
+ em = 1000000.0
+ ltvfbsdoff = 0
+ ll = 0
+ lw = 0
+ u0 = -0.00028230295310000003
+ w0 = 0
+ ua = -3.002357e-9
+ ub = 1.89239813e-18
+ uc = 1.5708441000000004e-10
+ ud = 0
+ phin = 0.15
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ pkt1 = 1.2683666000000002e-16
+ pkt2 = 1.019461e-15
+ ku0we = -0.0007
+ beta0 = 13
+ leta0 = -3.5803611e-8
+ letab = 5.4504443e-8
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ ppclm = -1.2878832e-14
+ rbdb = 50
+ pua1 = 1.04339e-23
+ prwb = 0
+ prwg = 0
+ pub1 = -1.3094356e-32
+ puc1 = -1.0640858600000001e-23
+ rbpb = 50
+ rbpd = 50
+ dlcig = 2.5e-9
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ bgidl = 2320000000.0
+ ptvfbsdoff = 0
+ rdsw = 100
+ ijthsfwd = 0.01
+ nfactor = 1
+ dmcgt = 0
+ tcjsw = 0.000357
+ ijthsrev = 0.01
+ toxref = 3e-9
+ rshg = 15.6
+ bigsd = 0.00125
+ )

.model nch_fs_32 nmos (
+ level = 54
+ eta0 = -0.25440451
+ etab = -0.81370191
+ scref = 1e-6
+ lku0we = 2.5e-11
+ pigcd = 2.621
+ epsrox = 3.9
+ aigsd = 0.010772817
+ njtsswg = 9
+ lvoff = -6.3427068e-9
+ rdsmod = 0
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ igbmod = 1
+ lvsat = -0.0013575165999999998
+ ckappad = 0.6
+ ckappas = 0.6
+ lvth0 = -7.221341000000012e-10
+ pdiblc1 = 0
+ pdiblc2 = 0.0069718933
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ pdiblcb = -0.3
+ delta = 0.007595625
+ laigc = 9.707156e-12
+ pbswgd = 0.95
+ pbswgs = 0.95
+ rnoia = 0
+ rnoib = 0
+ igcmod = 1
+ pketa = -6.053668000000001e-15
+ ngate = 8e+20
+ ngcon = 1
+ wpclm = 1.6305740000000013e-7
+ bigbacc = 0.002588
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ kvth0we = 0.00018
+ paigsd = -1.2154906e-23
+ lintnoi = -1.5e-8
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ ijthsfwd = 0.01
+ permod = 1
+ keta = -0.59506219
+ ijthsrev = 0.01
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 6.00154e-10
+ tvoff = 0.0034020192
+ kt1l = 0
+ voffcv = -0.16942
+ wpemod = 1
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ lint = 0
+ lkt1 = -1.9009946e-8
+ lkt2 = 1.0897551e-9
+ lmax = 4.5e-8
+ lmin = 3.6e-8
+ ku0we = -0.0007
+ nfactor = 1
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ beta0 = 13
+ leta0 = 2.6527632200000003e-8
+ letab = 2.5974719e-8
+ minv = -0.3
+ lua1 = 7.6118385e-17
+ lub1 = -1.3030425e-25
+ luc1 = -3.7246243e-17
+ ppclm = -8.780734400000002e-15
+ ndep = 1e+18
+ dlcig = 2.5e-9
+ lwlc = 0
+ tpbswg = 0.0009
+ bgidl = 2320000000.0
+ moin = 5.1
+ nigc = 3.083
+ nigbacc = 10
+ dmcgt = 0
+ pkvth0we = -1.3e-19
+ noff = 2.7195
+ tcjsw = 0.000357
+ ptvoff = -5.392468e-18
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ waigsd = 3.1116181e-12
+ nigbinv = 10
+ diomod = 1
+ ntox = 1.0
+ pcit = -3.4693290999999997e-17
+ vfbsdoff = 0.02
+ pclm = 1.46768105
+ bigsd = 0.00125
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 2.66208e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.66208e-10
+ phin = 0.15
+ wvoff = 6.255152000000001e-9
+ paramchk = 1
+ pkt1 = 5.4270205e-15
+ pkt2 = -4.1883975e-17
+ wvsat = -0.028736825999999997
+ wvth0 = -6.330829000000001e-9
+ fnoimod = 1
+ mjswgd = 0.85
+ mjswgs = 0.85
+ eigbinv = 1.1
+ waigc = 7.6854687e-11
+ tcjswg = 0.001
+ rbdb = 50
+ pua1 = -2.7889543e-23
+ prwb = 0
+ prwg = 0
+ pub1 = 4.4702459e-32
+ puc1 = 1.2190153e-23
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ pvfbsdoff = 0
+ lketa = 1.80561909e-8
+ ijthdfwd = 0.01
+ rdsw = 100
+ xpart = 1
+ egidl = 0.29734
+ cigbacc = 0.32875
+ ijthdrev = 0.01
+ fprout = 300
+ rshg = 15.6
+ xrcrg1 = 12
+ xrcrg2 = 1
+ tnoimod = 0
+ cigbinv = 0.006
+ wtvoff = 7.822084e-11
+ pvoff = -9.865003999999993e-17
+ version = 4.5
+ capmod = 2
+ tnom = 25
+ cdscb = 0
+ cdscd = 0
+ tempmod = 0
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ pvsat = 1.0650628200000002e-9
+ wku0we = 2e-11
+ lkvth0we = -2e-12
+ wk2we = 5e-12
+ pvth0 = -1.483420999999992e-17
+ drout = 0.56
+ mobmod = 0
+ wtvfbsdoff = 0
+ paigc = -2.6395467e-18
+ aigbacc = 0.02
+ voffl = 0
+ acnqsmod = 0
+ ltvfbsdoff = 0
+ weta0 = 8.5615058e-8
+ wetab = 2.2270081e-8
+ wags = 1.3153333e-7
+ lpclm = -1.8821805999999992e-8
+ wcit = 3.759659e-10
+ rbodymod = 0
+ aigbinv = 0.0163
+ voff = -0.061499972999999986
+ cgidl = 0.22
+ acde = 0.4
+ laigsd = 4.4039511e-17
+ vsat = 148854.172
+ wint = 0
+ vth0 = 0.347654671
+ wkt1 = -1.2742136999999998e-7
+ wkt2 = 7.8385579e-10
+ wmax = 5.374e-7
+ aigc = 0.011053515
+ wmin = 2.674e-7
+ pbswd = 0.8
+ pbsws = 0.8
+ ptvfbsdoff = 0
+ wpdiblc2 = 1.4081704e-10
+ wua1 = 6.7078609e-16
+ wub1 = -1.1020589000000001e-24
+ wuc1 = -3.0000411e-16
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ poxedge = 1
+ bigc = 0.001442
+ pdits = 0
+ wwlc = 0
+ cigsd = 0.069865
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ binunit = 2
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ ags = 2.6644444
+ cgsl = 3.31989e-12
+ pk2we = -1e-19
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ a0 = 10.55945905
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 101543.357
+ cf = 8.15e-11
+ cjd = 0.001281008
+ cit = -0.0081656108
+ cjs = 0.001281008
+ clc = 1e-7
+ ef = 1.0
+ k1 = 0.274
+ cle = 0.6
+ k2 = 0.037527322
+ k3 = -1.8419
+ em = 1000000.0
+ bvd = 8.7
+ bvs = 8.7
+ ll = 0
+ lw = 0
+ dlc = 3.26497e-9
+ u0 = 0.006433017400000001
+ w0 = 0
+ k3b = 1.9326
+ ua = -1.7148580999999998e-9
+ ub = 1.250859149999999e-18
+ uc = 5.4381728e-10
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ dwb = 0
+ ww = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ xw = 8.600000000000001e-9
+ wkvth0we = 2e-12
+ tnoia = 0
+ toxref = 3e-9
+ peta0 = -4.1184253e-15
+ la0 = -4.65319969e-7
+ trnqsmod = 0
+ petab = -7.719916e-16
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.0016482648800000001
+ kt1 = 0.12069622
+ lk2 = -4.2131932e-9
+ kt2 = -0.11741295
+ wketa = 1.87190595e-7
+ llc = 0
+ lln = 1
+ lu0 = 1.8825002000000003e-10
+ mjd = 0.26
+ lua = 1.6761980000000137e-18
+ mjs = 0.26
+ lub = 8.339062399999967e-27
+ luc = -2.98810456e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ tpbsw = 0.0019
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 9.065128000000001e-14
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ nsd = 1e+20
+ pbd = 0.52
+ pat = -3.0248428e-10
+ pbs = 0.52
+ pk2 = 5.9540883e-16
+ cjswd = 7.7408e-11
+ cjsws = 7.7408e-11
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ pu0 = -7.7700919e-17
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ prt = 0
+ pua = -1.6092489999999997e-23
+ pub = 1.5276544400000003e-32
+ puc = 5.518326299999999e-24
+ pud = 0
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = -1.1935669e-9
+ ub1 = 2.1692222300000005e-18
+ uc1 = 1.0139469700000001e-9
+ tpb = 0.0014
+ k2we = 5e-5
+ wa0 = -2.59429679e-6
+ tvfbsdoff = 0.022
+ ute = -1
+ wat = 0.0028451685
+ dsub = 0.75
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -1.1593839e-8
+ ltvoff = -1.1952424e-10
+ dtox = 2.7e-10
+ wlc = 0
+ wln = 1
+ rgatemod = 0
+ wu0 = 1.18710292e-9
+ xgl = -1.09e-8
+ xgw = 0
+ wua = 3.2583921000000013e-16
+ wub = -3.447615700000002e-25
+ wuc = -8.750290400000002e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ tnjtsswg = 1
+ )

.model nch_fs_33 nmos (
+ level = 54
+ rbodymod = 0
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ version = 4.5
+ pbswgd = 0.95
+ pbswgs = 0.95
+ ntox = 1.0
+ pcit = -1.2000000000000001e-17
+ pclm = 1.8851852
+ tempmod = 0
+ igcmod = 1
+ phin = 0.15
+ aigbacc = 0.02
+ pkt1 = 5.600000000000001e-17
+ wpdiblc2 = -2.9834e-10
+ pvoff = 0
+ cdscb = 0
+ cdscd = 0
+ pvsat = -2.24e-11
+ aigbinv = 0.0163
+ rbdb = 50
+ prwb = 0
+ prwg = 0
+ pub1 = -3.2e-34
+ wk2we = 5e-12
+ pvth0 = -1.2e-16
+ drout = 0.56
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ rdsw = 100
+ permod = 1
+ voffl = 0
+ weta0 = 0
+ wkvth0we = 2e-12
+ cgidl = 0.22
+ trnqsmod = 0
+ voffcv = -0.16942
+ wpemod = 1
+ poxedge = 1
+ rshg = 15.6
+ binunit = 2
+ pbswd = 0.8
+ pbsws = 0.8
+ rgatemod = 0
+ tnjtsswg = 1
+ tnom = 25
+ pdits = 0
+ ags = 0.6088259300000001
+ cigsd = 0.069865
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ tpbswg = 0.0009
+ cjd = 0.001281008
+ dvt0w = 0
+ cit = 0.002342713
+ dvt1w = 0
+ cjs = 0.001281008
+ clc = 1e-7
+ cle = 0.6
+ dvt2w = 0
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 9.8024918e-9
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ jtsswgd = 2.3e-7
+ pk2we = -1e-19
+ jtsswgs = 2.3e-7
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ la0 = 0
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.00016
+ kt1 = -0.21767878
+ kt2 = -0.055117852
+ ptvoff = 0
+ llc = 0
+ lln = 1
+ lu0 = 9.600000000000001e-12
+ wags = 8.994443999999999e-9
+ mjd = 0.26
+ mjs = 0.26
+ lub = 0
+ lud = 0
+ lwc = 0
+ waigsd = 3.1789128e-12
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 0
+ tnoia = 0
+ nsd = 1e+20
+ pbd = 0.52
+ pat = -3.04e-11
+ wcit = -2.1566928e-10
+ pbs = 0.52
+ pu0 = 1.8400000000000002e-18
+ prt = 0
+ pub = 0
+ pud = 0
+ peta0 = 0.0
+ diomod = 1
+ voff = -0.095952978
+ acde = 0.4
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 9.5347726e-10
+ wketa = -1.1490089e-9
+ ub1 = -5.3850981e-19
+ uc1 = -6.0041111e-11
+ tpb = 0.0014
+ tpbsw = 0.0019
+ pditsd = 0
+ pditsl = 0
+ vsat = 84306.193
+ wa0 = 0
+ cjswgd = 2.66208e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.66208e-10
+ wint = 0
+ ute = -1
+ wat = 0
+ vth0 = 0.28549411
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 3.0219344e-9
+ cjswd = 7.7408e-11
+ cjsws = 7.7408e-11
+ wlc = 0
+ wln = 1
+ wu0 = -1.2693333000000005e-11
+ wkt1 = -3.4514582500000003e-9
+ wkt2 = 1.0235511e-10
+ xgl = -1.09e-8
+ mjswd = 0.11
+ xgw = 0
+ mjsws = 0.11
+ wua = -1.6467997e-17
+ wub = 3.619626e-26
+ wuc = -1.4955111e-18
+ wud = 0
+ agidl = 9.41e-8
+ wmax = 2.674e-7
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ aigc = 0.01181895
+ wmin = 1.08e-7
+ tvfbsdoff = 0.022
+ njtsswg = 9
+ mjswgd = 0.85
+ mjswgs = 0.85
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ wua1 = -3.1223388e-18
+ wub1 = 2.0807554e-26
+ wuc1 = 8.1864667e-18
+ tcjswg = 0.001
+ bigc = 0.001442
+ ckappad = 0.6
+ ckappas = 0.6
+ wwlc = 0
+ pdiblc1 = 0
+ pdiblc2 = 0.023869018
+ pdiblcb = -0.3
+ scref = 1e-6
+ cdsc = 0
+ ijthsfwd = 0.01
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ pigcd = 2.621
+ aigsd = 0.010772573
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ lvoff = -1.6e-11
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ bigbacc = 0.002588
+ lvsat = -0.0002
+ lvth0 = -4.8e-10
+ fprout = 300
+ ijthsrev = 0.01
+ delta = 0.007595625
+ xrcrg1 = 12
+ xrcrg2 = 1
+ kvth0we = 0.00018
+ rnoia = 0
+ rnoib = 0
+ lintnoi = -1.5e-8
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ wtvoff = 2.5061202e-10
+ ngate = 8e+20
+ wtvfbsdoff = 0
+ ngcon = 1
+ wpclm = -9.7111111e-9
+ k2we = 5e-5
+ dsub = 0.75
+ dtox = 2.7e-10
+ gbmin = 1e-12
+ capmod = 2
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ ltvfbsdoff = 0
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ wku0we = 2e-11
+ mobmod = 0
+ eta0 = 0.2
+ etab = -0.2
+ pkvth0we = -1.3e-19
+ nfactor = 1
+ ptvfbsdoff = 0
+ tvoff = 0.00085486634
+ vfbsdoff = 0.02
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ paramchk = 1
+ nigbacc = 10
+ ku0we = -0.0007
+ beta0 = 13
+ leta0 = 1.6000000000000003e-9
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ dlcig = 2.5e-9
+ nigbinv = 10
+ bgidl = 2320000000.0
+ ijthdfwd = 0.01
+ keta = -0.021050128
+ dmcgt = 0
+ tcjsw = 0.000357
+ toxref = 3e-9
+ ijthdrev = 0.01
+ fnoimod = 1
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = -8e-12
+ eigbinv = 1.1
+ kt1l = 0
+ bigsd = 0.00125
+ lint = 6.5375218e-9
+ lkt1 = -4.8e-10
+ wvoff = 2.9681533e-9
+ lmax = 2.001e-5
+ lmin = 8.9991e-6
+ ltvoff = 0
+ lpe0 = 9.2e-8
+ wvsat = 0.002322956
+ lpeb = 2.5e-7
+ wvth0 = -6.7513739000000004e-9
+ a0 = 3.5
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 200000
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.014356400999999998
+ k3 = -1.8419
+ em = 1000000.0
+ minv = -0.3
+ waigc = 1.7818122e-11
+ ll = 0
+ lw = 0
+ u0 = 0.012655556
+ w0 = 0
+ lub1 = -2.4000000000000004e-27
+ ua = -2.0911548e-9
+ ub = 2.2368542e-18
+ uc = 5.8018519e-11
+ ud = 0
+ cigbacc = 0.32875
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ ndep = 1e+18
+ lkvth0we = -2e-12
+ pvfbsdoff = 0
+ lwlc = 0
+ moin = 5.1
+ lku0we = 2.5e-11
+ tnoimod = 0
+ epsrox = 3.9
+ xpart = 1
+ nigc = 3.083
+ cigbinv = 0.006
+ acnqsmod = 0
+ rdsmod = 0
+ egidl = 0.29734
+ igbmod = 1
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ )

.model nch_fs_34 nmos (
+ level = 54
+ paramchk = 1
+ wpclm = -9.7111111e-9
+ gbmin = 1e-12
+ wua1 = -1.7574281e-19
+ wub1 = 1.7597088e-26
+ wuc1 = 8.3134424e-18
+ jswgd = 1.28e-13
+ nfactor = 1
+ jswgs = 1.28e-13
+ paigsd = -3.8370159e-23
+ bigc = 0.001442
+ wwlc = 0
+ permod = 1
+ cdsc = 0
+ ijthdfwd = 0.01
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ nigbacc = 10
+ ijthdrev = 0.01
+ voffcv = -0.16942
+ wpemod = 1
+ tvoff = 0.00082419905
+ lpdiblc2 = -9.2950492e-9
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ nigbinv = 10
+ k2we = 5e-5
+ ku0we = -0.0007
+ beta0 = 13
+ dsub = 0.75
+ leta0 = 1.6000000000000003e-9
+ dtox = 2.7e-10
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ tpbswg = 0.0009
+ fnoimod = 1
+ lkvth0we = -2e-12
+ eigbinv = 1.1
+ dlcig = 2.5e-9
+ eta0 = 0.2
+ bgidl = 2320000000.0
+ etab = -0.2
+ acnqsmod = 0
+ ptvoff = -2.3727895e-16
+ waigsd = 3.1789171e-12
+ dmcgt = 0
+ tcjsw = 0.000357
+ rbodymod = 0
+ diomod = 1
+ cigbacc = 0.32875
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 2.66208e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.66208e-10
+ bigsd = 0.00125
+ tnoimod = 0
+ wvoff = 3.141381e-9
+ mjswgd = 0.85
+ mjswgs = 0.85
+ cigbinv = 0.006
+ wvsat = 0.002322956
+ wvth0 = -6.936365900000001e-9
+ wpdiblc2 = -6.4961636e-10
+ tcjswg = 0.001
+ waigc = 1.8291238e-11
+ pvfbsdoff = 0
+ version = 4.5
+ lketa = -2.7750915e-8
+ tempmod = 0
+ xpart = 1
+ egidl = 0.29734
+ aigbacc = 0.02
+ keta = -0.017963263
+ wkvth0we = 2e-12
+ wtvfbsdoff = 0
+ fprout = 300
+ lags = 4.3821463e-7
+ xrcrg1 = 12
+ xrcrg2 = 1
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = -1.7265105499999998e-11
+ trnqsmod = 0
+ kt1l = 0
+ ltvfbsdoff = 0
+ aigbinv = 0.0163
+ wtvoff = 2.7700567e-10
+ lint = 6.5375218e-9
+ lkt1 = -8.9298468e-8
+ lkt2 = -1.6837724e-8
+ lmax = 8.9991e-6
+ lmin = 8.9908e-7
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ capmod = 2
+ rgatemod = 0
+ pvoff = -1.5573172e-15
+ tnjtsswg = 1
+ wku0we = 2e-11
+ minv = -0.3
+ lua1 = -7.4262143e-17
+ lub1 = -1.4398035e-25
+ luc1 = 6.2830403e-17
+ cdscb = 0
+ cdscd = 0
+ mobmod = 0
+ pvsat = -2.24e-11
+ ndep = 1e+18
+ wk2we = 5e-12
+ pvth0 = 1.5430782e-15
+ ptvfbsdoff = 0
+ drout = 0.56
+ lwlc = 0
+ poxedge = 1
+ moin = 5.1
+ paigc = -4.2533129e-18
+ nigc = 3.083
+ voffl = 0
+ binunit = 2
+ weta0 = 0
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ laigsd = 3.3658034e-16
+ pags = 5.2134206e-15
+ cgidl = 0.22
+ ntox = 1.0
+ pcit = 6.7881874e-17
+ pclm = 1.8851852
+ phin = 0.15
+ pbswd = 0.8
+ pbsws = 0.8
+ ags = 0.5600812500000001
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ pkt1 = -3.0816964e-16
+ pkt2 = -1.7740443e-15
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ cjd = 0.001281008
+ cit = 0.0023437436
+ cjs = 0.001281008
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 9.8024918e-9
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ pdits = 0
+ cigsd = 0.069865
+ rbdb = 50
+ pua1 = -2.6489898e-23
+ prwb = 0
+ prwg = 0
+ pub1 = 2.854209e-32
+ puc1 = -1.1415122e-24
+ dvt0w = 0
+ la0 = -1.6207075e-6
+ dvt1w = 0
+ dvt2w = 0
+ rbpb = 50
+ rbpd = 50
+ jsd = 6.11e-7
+ rbps = 50
+ jss = 6.11e-7
+ lat = -0.043382769
+ rbsb = 50
+ pvag = 1.2
+ kt1 = -0.20779908
+ lk2 = -1.5849432e-8
+ kt2 = -0.053244913
+ llc = 0
+ lln = 1
+ lu0 = -1.6696432e-9
+ mjd = 0.26
+ lua = -1.2813977e-16
+ mjs = 0.26
+ lub = -8.5009677e-26
+ luc = -2.2547224e-17
+ lud = 0
+ ijthsfwd = 0.01
+ lwc = 0
+ lwl = 0
+ rdsw = 100
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 3.8370159e-14
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 3.9600965e-9
+ pbs = 0.52
+ pk2 = -8.7965669e-16
+ pk2we = -1e-19
+ pu0 = 1.839999999998372e-18
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ prt = 0
+ pua = -3.3674591e-24
+ pub = -4.9159389e-33
+ puc = 2.3789498e-24
+ pud = 0
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 9.6173779e-10
+ ub1 = -5.2276116e-19
+ uc1 = -6.7030033e-11
+ njtsswg = 9
+ tpb = 0.0014
+ toxref = 3e-9
+ wa0 = -4.2680933e-9
+ tnoia = 0
+ ute = -1
+ wat = -0.0004438817
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 3.1197827e-9
+ wlc = 0
+ wln = 1
+ wu0 = -1.2693333000000005e-11
+ ijthsrev = 0.01
+ xgl = -1.09e-8
+ xtsswgd = 0.18
+ xgw = 0
+ xtsswgs = 0.18
+ wua = -1.6093419e-17
+ wub = 3.6743083e-26
+ wuc = -1.7601329e-18
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ peta0 = 0.0
+ wketa = -1.4921751e-9
+ ckappad = 0.6
+ ckappas = 0.6
+ rshg = 15.6
+ pdiblc1 = 0
+ pdiblc2 = 0.02490295
+ tpbsw = 0.0019
+ pdiblcb = -0.3
+ cjswd = 7.7408e-11
+ cjsws = 7.7408e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ tvfbsdoff = 0.022
+ ltvoff = 2.7569894e-10
+ ppdiblc2 = 3.1579745e-15
+ bigbacc = 0.002588
+ tnom = 25
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ kvth0we = 0.00018
+ lku0we = 2.5e-11
+ epsrox = 3.9
+ scref = 1e-6
+ lintnoi = -1.5e-8
+ pigcd = 2.621
+ bigbinv = 0.004953
+ aigsd = 0.010772573
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ rdsmod = 0
+ wvfbsdoff = 0
+ igbmod = 1
+ lvoff = -1.4754881e-8
+ lvfbsdoff = 0
+ pkvth0we = -1.3e-19
+ wags = 8.414531e-9
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ lvsat = -0.0002
+ wcit = -2.2455490999999997e-10
+ lvth0 = 5.613542e-8
+ pbswgd = 0.95
+ pbswgs = 0.95
+ voff = -0.094313503
+ delta = 0.007595625
+ laigc = -1.6452737e-10
+ acde = 0.4
+ a0 = 3.6802789
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ vfbsdoff = 0.02
+ igcmod = 1
+ at = 204807.87
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.016119408
+ k3 = -1.8419
+ em = 1000000.0
+ rnoia = 0
+ rnoib = 0
+ ll = 0
+ lw = 0
+ vsat = 84306.193
+ u0 = 0.012842346
+ w0 = 0
+ wint = 0
+ ua = -2.0769012e-9
+ ub = 2.2463102e-18
+ uc = 6.0526552e-11
+ ud = 0
+ vth0 = 0.27919651
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ wkt1 = -3.4109499500000005e-9
+ wkt2 = 2.996904e-10
+ wmax = 2.674e-7
+ aigc = 0.011837251
+ wmin = 1.08e-7
+ pketa = 3.0850638e-15
+ ngate = 8e+20
+ ngcon = 1
+ )

.model nch_fs_35 nmos (
+ level = 54
+ a0 = 2.7573663
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ voffl = 0
+ at = 225908.74
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.009086581
+ k3 = -1.8419
+ em = 1000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.012432289999999999
+ w0 = 0
+ ua = -2.2251639e-9
+ ub = 2.3450974e-18
+ uc = 3.6825844e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ weta0 = 0
+ keta = -0.063873893
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ voffcv = -0.16942
+ wpemod = 1
+ lags = -4.2829945e-7
+ ijthsrev = 0.01
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ cgidl = 0.22
+ lcit = -6.2690204e-10
+ kt1l = 0
+ ags = 1.5336926
+ cjd = 0.001281008
+ cit = 0.0030287289
+ cjs = 0.001281008
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 9.8024918e-9
+ k3b = 1.9326
+ lint = 6.5375218e-9
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ lkt1 = 4.8571427e-8
+ lkt2 = -1.4519819e-8
+ pbswd = 0.8
+ pbsws = 0.8
+ lmax = 8.9908e-7
+ lmin = 4.4908e-7
+ lpe0 = 9.2e-8
+ la0 = -7.9931523e-7
+ lpeb = 2.5e-7
+ jsd = 6.11e-7
+ ppdiblc2 = -1.3141262e-15
+ jss = 6.11e-7
+ lat = -0.062162545
+ kt1 = -0.36270908
+ lk2 = -9.5902228e-9
+ kt2 = -0.0558493
+ llc = 0
+ lln = 1
+ lu0 = -1.3046934e-9
+ njtsswg = 9
+ mjd = 0.26
+ lua = 3.8140531e-18
+ mjs = 0.26
+ lub = -1.7293024e-25
+ luc = -1.4535934e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ tpbswg = 0.0009
+ njd = 1.02
+ minv = -0.3
+ njs = 1.02
+ pa0 = -6.7606598e-14
+ lua1 = -1.6437259e-16
+ lub1 = 2.0418042999999997e-26
+ nsd = 1e+20
+ pdits = 0
+ luc1 = 5.6450349e-17
+ pbd = 0.52
+ pat = 1.6728657e-9
+ pbs = 0.52
+ pk2 = -2.3173279e-16
+ cigsd = 0.069865
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ pu0 = 1.0797874200000001e-17
+ prt = 0
+ ndep = 1e+18
+ pua = -1.9061799e-24
+ pub = 1.3958464e-33
+ puc = -1.352132e-24
+ pud = 0
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ lwlc = 0
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 1.0629855e-9
+ ckappad = 0.6
+ ub1 = -7.0747845e-19
+ moin = 5.1
+ uc1 = -5.9861432e-11
+ ckappas = 0.6
+ tpb = 0.0014
+ pdiblc1 = 0
+ pdiblc2 = 0.01020022
+ pdiblcb = -0.3
+ wa0 = 1.1480691e-7
+ ute = -1
+ nigc = 3.083
+ wat = 0.0021260405
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 2.3917793e-9
+ wlc = 0
+ pk2we = -1e-19
+ ptvoff = -4.8469984e-16
+ wln = 1
+ wu0 = -2.2758360000000004e-11
+ xgl = -1.09e-8
+ dvtp0 = 4e-7
+ xgw = 0
+ dvtp1 = 0.01
+ wua = -1.7735306e-17
+ wub = 2.9651178e-26
+ wuc = 2.4320938e-18
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ waigsd = 3.178874e-12
+ pkvth0we = -1.3e-19
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ tnoia = 0
+ diomod = 1
+ bigbacc = 0.002588
+ peta0 = 0.0
+ pags = -9.2425378e-15
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 2.66208e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.66208e-10
+ wketa = 5.5022601e-9
+ vfbsdoff = 0.02
+ ntox = 1.0
+ pcit = 1.468079e-16
+ pclm = 1.8851852
+ tpbsw = 0.0019
+ kvth0we = 0.00018
+ cjswd = 7.7408e-11
+ cjsws = 7.7408e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ phin = 0.15
+ tvfbsdoff = 0.022
+ lintnoi = -1.5e-8
+ bigbinv = 0.004953
+ mjswgd = 0.85
+ mjswgs = 0.85
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ paramchk = 1
+ pkt1 = -1.3155355000000001e-14
+ pkt2 = 1.7857928e-15
+ tcjswg = 0.001
+ wtvfbsdoff = 0
+ rbdb = 50
+ pua1 = 3.1539092e-23
+ prwb = 0
+ prwg = 0
+ pub1 = -3.1853886e-32
+ puc1 = -7.798421e-24
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ scref = 1e-6
+ ijthdfwd = 0.01
+ rdsw = 100
+ pigcd = 2.621
+ aigsd = 0.010772573
+ ltvfbsdoff = 0
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ lvoff = -2.8472354000000002e-8
+ fprout = 300
+ lvsat = -0.0002
+ xrcrg1 = 12
+ xrcrg2 = 1
+ lvth0 = 1.8274806e-8
+ ijthdrev = 0.01
+ delta = 0.007595625
+ nfactor = 1
+ laigc = -6.1235169e-11
+ lpdiblc2 = 3.7903799e-9
+ rshg = 15.6
+ rnoia = 0
+ rnoib = 0
+ wtvoff = 5.5500668e-10
+ ptvfbsdoff = 0
+ pketa = -3.1399835e-15
+ ngate = 8e+20
+ ngcon = 1
+ wpclm = -9.7111111e-9
+ capmod = 2
+ wku0we = 2e-11
+ gbmin = 1e-12
+ nigbacc = 10
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ mobmod = 0
+ tnom = 25
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ lkvth0we = -2e-12
+ nigbinv = 10
+ acnqsmod = 0
+ wags = 2.4657181000000002e-8
+ rbodymod = 0
+ wcit = -3.1323583999999997e-10
+ voff = -0.078900611
+ tvoff = -3.4914836e-5
+ acde = 0.4
+ fnoimod = 1
+ xjbvd = 1
+ xjbvs = 1
+ vsat = 84306.193
+ lk2we = -1.5e-12
+ eigbinv = 1.1
+ wint = 0
+ vth0 = 0.32173651999999997
+ wkt1 = 1.1024089999999999e-8
+ wkt2 = -3.7001265e-9
+ wmax = 2.674e-7
+ aigc = 0.011721192
+ wmin = 1.08e-7
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ ku0we = -0.0007
+ beta0 = 13
+ leta0 = 1.6000000000000003e-9
+ wpdiblc2 = 4.3752159e-9
+ wua1 = -6.5376855e-17
+ wub1 = 8.5457734e-26
+ wuc1 = 1.5793115e-17
+ bigc = 0.001442
+ wwlc = 0
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ cigbacc = 0.32875
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ tnoimod = 0
+ cigc = 0.000625
+ toxref = 3e-9
+ dmcgt = 0
+ tcjsw = 0.000357
+ wkvth0we = 2e-12
+ cigbinv = 0.006
+ trnqsmod = 0
+ bigsd = 0.00125
+ version = 4.5
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ tempmod = 0
+ ltvoff = 1.0403103e-9
+ wvoff = -2.1121636e-9
+ k2we = 5e-5
+ wvsat = 0.002322956
+ aigbacc = 0.02
+ dsub = 0.75
+ wvth0 = -3.4014741000000007e-9
+ dtox = 2.7e-10
+ rgatemod = 0
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ tnjtsswg = 1
+ waigc = 1.00872e-11
+ pvfbsdoff = 0
+ lku0we = 2.5e-11
+ epsrox = 3.9
+ eta0 = 0.2
+ etab = -0.2
+ lketa = 1.3109546e-8
+ aigbinv = 0.0163
+ xpart = 1
+ rdsmod = 0
+ igbmod = 1
+ egidl = 0.29734
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ pbswgd = 0.95
+ pbswgs = 0.95
+ igcmod = 1
+ poxedge = 1
+ binunit = 2
+ pvoff = 3.1183375e-15
+ cdscb = 0
+ cdscd = 0
+ pvsat = -2.24e-11
+ wk2we = 5e-12
+ pvth0 = -1.6029756e-15
+ drout = 0.56
+ permod = 1
+ paigc = 3.0482801e-18
+ ijthsfwd = 0.01
+ )

.model nch_fs_36 nmos (
+ level = 54
+ rshg = 15.6
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ cigbacc = 0.32875
+ tnoimod = 0
+ ku0we = -0.0007
+ a0 = 2.8517872
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ beta0 = 13
+ at = 72186.119
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.0025801551000000002
+ k3 = -1.8419
+ em = 1000000.0
+ leta0 = 1.6000000000000003e-9
+ rgatemod = 0
+ ll = -1.18e-13
+ lw = 0
+ u0 = 0.010648434
+ tpbswg = 0.0009
+ w0 = 0
+ ua = -2.2247872e-9
+ ub = 2.0937783e-18
+ uc = 7.1203963e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ tnjtsswg = 1
+ ww = 0
+ xw = 8.600000000000001e-9
+ cigbinv = 0.006
+ tnom = 25
+ ppclm = 2.75592e-14
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ ptvoff = 2.8225911e-16
+ version = 4.5
+ waigsd = 3.178874e-12
+ tempmod = 0
+ dmcgt = 0
+ tcjsw = 0.000357
+ diomod = 1
+ wags = 2.3808180000000002e-7
+ aigbacc = 0.02
+ wcit = 2.2683634e-10
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 2.66208e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.66208e-10
+ voff = -0.13810998
+ acde = 0.4
+ bigsd = 0.00125
+ vsat = 84306.193
+ wint = 0
+ vth0 = 0.38435442
+ wtvfbsdoff = 0
+ wkt1 = -4.1130622999999995e-8
+ wkt2 = -4.3121065e-11
+ aigbinv = 0.0163
+ wmax = 2.674e-7
+ mjswgd = 0.85
+ mjswgs = 0.85
+ aigc = 0.011581706
+ wmin = 1.08e-7
+ wvoff = 7.1640927e-9
+ tcjswg = 0.001
+ wvsat = 0.002322956
+ ltvfbsdoff = 0
+ wvth0 = -9.1496131e-9
+ wua1 = 2.3276683e-17
+ wub1 = 1.5603072e-26
+ wuc1 = -5.1034561e-18
+ waigc = 2.6093343e-11
+ pvfbsdoff = 0
+ bigc = 0.001442
+ wwlc = 0
+ lketa = -3.8407777e-8
+ ijthsfwd = 0.01
+ cdsc = 0
+ xpart = 1
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ poxedge = 1
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ egidl = 0.29734
+ fprout = 300
+ ptvfbsdoff = 0
+ binunit = 2
+ xrcrg1 = 12
+ xrcrg2 = 1
+ ijthsrev = 0.01
+ wtvoff = -1.1880818e-9
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ capmod = 2
+ k2we = 5e-5
+ wku0we = 2e-11
+ ppdiblc2 = 3.3310302e-16
+ dsub = 0.75
+ dtox = 2.7e-10
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ pvoff = -9.6321526e-16
+ mobmod = 0
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ cdscb = 0
+ cdscd = 0
+ pvsat = -2.24e-11
+ wk2we = 5e-12
+ pvth0 = 9.262056000000001e-16
+ drout = 0.56
+ eta0 = 0.2
+ etab = -0.2
+ paigc = -3.9944226e-18
+ voffl = 0
+ weta0 = 0
+ pkvth0we = -1.3e-19
+ ags = -2.6547885
+ lpclm = -2.4174737e-7
+ cjd = 0.001281008
+ cit = 0.00083484714
+ cjs = 0.001281008
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 1.30529375e-8
+ k3b = 1.9326
+ njtsswg = 9
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ cgidl = 0.22
+ vfbsdoff = 0.02
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ la0 = -8.4086042e-7
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = 0.0054754098
+ kt1 = -0.088256509
+ lk2 = -6.7273888e-9
+ kt2 = -0.075738087
+ ckappad = 0.6
+ ckappas = 0.6
+ llc = -1.18e-13
+ lln = 0.7
+ lu0 = -5.197967099999999e-10
+ mjd = 0.26
+ pdiblc1 = 0
+ pdiblc2 = 0.031716534
+ lua = 3.6483177e-18
+ mjs = 0.26
+ lub = -6.2349821e-26
+ luc = -1.6579966e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ pdiblcb = -0.3
+ njd = 1.02
+ njs = 1.02
+ pa0 = 8.661463e-14
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ pbswd = 0.8
+ pbsws = 0.8
+ nsd = 1e+20
+ pbd = 0.52
+ pat = -3.1722679e-9
+ pbs = 0.52
+ pk2 = -2.2869691e-16
+ paramchk = 1
+ pu0 = 4.2809578e-18
+ prt = 0
+ pua = -4.9144669e-25
+ pub = 1.8790045e-33
+ puc = 1.8346553e-24
+ pud = 0
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 5.8363721e-10
+ ub1 = -5.3348382e-19
+ uc1 = 8.6067289e-11
+ tpb = 0.0014
+ wa0 = -2.3569588e-7
+ ute = -1
+ wat = 0.013137708
+ pdits = 0
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 2.3848778e-9
+ wlc = 0
+ wln = 1
+ cigsd = 0.069865
+ wu0 = -7.947187000000004e-12
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -2.0950609e-17
+ wub = 2.8553091e-26
+ wuc = -4.8106046e-18
+ wud = 0
+ wwc = 0
+ bigbacc = 0.002588
+ wwl = 0
+ wwn = 1
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ ijthdfwd = 0.01
+ kvth0we = 0.00018
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ toxref = 3e-9
+ lintnoi = -1.5e-8
+ keta = 0.053210932
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ tnoia = 0
+ lags = 1.4146322e-6
+ ijthdrev = 0.01
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ peta0 = 0.0
+ lcit = 3.3840592e-10
+ wketa = -7.2433388e-9
+ kt1l = 0
+ lpdiblc2 = -5.676798e-9
+ tpbsw = 0.0019
+ cjswd = 7.7408e-11
+ cjsws = 7.7408e-11
+ mjswd = 0.11
+ tvfbsdoff = 0.022
+ mjsws = 0.11
+ ltvoff = -1.663256e-9
+ agidl = 9.41e-8
+ lint = 9.7879675e-9
+ lkt1 = -7.2187703e-8
+ lkt2 = -5.7687528e-9
+ lmax = 4.4908e-7
+ lmin = 2.1577e-7
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ minv = -0.3
+ lku0we = 2.5e-11
+ lua1 = 4.6540649e-17
+ lub1 = -5.6139597e-26
+ luc1 = -7.7582888e-18
+ epsrox = 3.9
+ lkvth0we = -2e-12
+ ndep = 1e+18
+ nfactor = 1
+ lwlc = 0
+ moin = 5.1
+ scref = 1e-6
+ rdsmod = 0
+ pigcd = 2.621
+ nigc = 3.083
+ igbmod = 1
+ aigsd = 0.010772573
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ acnqsmod = 0
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ lvoff = -2.4202325e-9
+ pbswgd = 0.95
+ noff = 2.7195
+ pbswgs = 0.95
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ lvsat = -0.0002
+ rbodymod = 0
+ lvth0 = -9.2770687e-9
+ igcmod = 1
+ nigbacc = 10
+ delta = 0.007595625
+ pags = -1.0314937e-13
+ laigc = 1.3898222e-13
+ ntox = 1.0
+ pcit = -9.082386e-17
+ pclm = 2.434611
+ rnoia = 0
+ rnoib = 0
+ phin = 0.15
+ pketa = 2.46808e-15
+ ngate = 8e+20
+ nigbinv = 10
+ ngcon = 1
+ wpclm = -7.2345657e-8
+ pkt1 = 9.7927187e-15
+ pkt2 = 1.7671038e-16
+ wpdiblc2 = 6.3151306e-10
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ permod = 1
+ rbdb = 50
+ pua1 = -7.4684646e-24
+ prwb = 0
+ prwg = 0
+ pub1 = -1.1178346e-33
+ puc1 = 1.3960704e-24
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ fnoimod = 1
+ rdsw = 100
+ eigbinv = 1.1
+ wkvth0we = 2e-12
+ voffcv = -0.16942
+ wpemod = 1
+ trnqsmod = 0
+ tvoff = 0.006109554
+ )

.model nch_fs_37 nmos (
+ level = 54
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ pdits = 0
+ cigsd = 0.069865
+ lkvth0we = -2e-12
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ eta0 = 0.2
+ etab = -0.2
+ ptvoff = -1.8615536e-17
+ waigsd = 3.178874e-12
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ acnqsmod = 0
+ diomod = 1
+ wtvfbsdoff = 0
+ tnoia = 0
+ pditsd = 0
+ pditsl = 0
+ rbodymod = 0
+ cjswgd = 2.66208e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.66208e-10
+ a0 = -2.4455841
+ a1 = 0
+ a2 = 1
+ peta0 = 0.0
+ b0 = 0
+ b1 = 0
+ ltvfbsdoff = 0
+ at = 121458.51
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = -0.0069973019999999995
+ k3 = -1.8419
+ em = 1000000.0
+ ll = -1.18e-13
+ wketa = 1.5290605e-8
+ lw = 0
+ u0 = 0.009044212999999999
+ w0 = 0
+ ua = -2.2679307e-9
+ ub = 1.903479518e-18
+ uc = 2.5998306e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ tpbsw = 0.0019
+ nfactor = 1
+ tvfbsdoff = 0.022
+ cjswd = 7.7408e-11
+ cjsws = 7.7408e-11
+ mjswgd = 0.85
+ mjswd = 0.11
+ mjswgs = 0.85
+ mjsws = 0.11
+ agidl = 9.41e-8
+ tcjswg = 0.001
+ wpdiblc2 = 2.0871493e-9
+ ptvfbsdoff = 0
+ nigbacc = 10
+ scref = 1e-6
+ wvfbsdoff = 0
+ pigcd = 2.621
+ lvfbsdoff = 0
+ aigsd = 0.010772573
+ fprout = 300
+ lvoff = 4.8514199999999965e-11
+ nigbinv = 10
+ keta = -0.11923047
+ xrcrg1 = 12
+ xrcrg2 = 1
+ wkvth0we = 2e-12
+ lvsat = -0.0005892742949999998
+ lvth0 = -8.3419377e-9
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ trnqsmod = 0
+ delta = 0.007595625
+ lcit = -4.7333293e-11
+ wtvoff = 2.3786433e-10
+ laigc = -6.7426314e-12
+ kt1l = 0
+ rnoia = 0
+ rnoib = 0
+ fnoimod = 1
+ lint = 9.7879675e-9
+ pketa = -2.286582e-15
+ ngate = 8e+20
+ capmod = 2
+ eigbinv = 1.1
+ lkt1 = 7.879381000000001e-11
+ lkt2 = 1.6714521e-10
+ lmax = 2.1577e-7
+ ngcon = 1
+ lmin = 9e-8
+ wpclm = 1.5314007e-7
+ wku0we = 2e-11
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ mobmod = 0
+ rgatemod = 0
+ gbmin = 1e-12
+ tnjtsswg = 1
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ minv = -0.3
+ lua1 = -6.7367772e-18
+ lub1 = -4.0761216e-26
+ luc1 = -1.0970607e-17
+ ndep = 1e+18
+ lwlc = 0
+ moin = 5.1
+ nigc = 3.083
+ cigbacc = 0.32875
+ tnoimod = 0
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ cigbinv = 0.006
+ tvoff = -0.0028392003
+ ntox = 1.0
+ pcit = 2.9405719999999994e-18
+ pclm = 1.0592301
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ phin = 0.15
+ version = 4.5
+ tempmod = 0
+ pkt1 = -1.3029532999999997e-16
+ pkt2 = -2.0087744e-16
+ ku0we = -0.0007
+ beta0 = 13
+ leta0 = 1.6000000000000003e-9
+ ppclm = -2.0018289e-14
+ aigbacc = 0.02
+ rbdb = 50
+ pua1 = 2.2068447e-24
+ prwb = 0
+ prwg = 0
+ pub1 = -3.0626774000000002e-33
+ puc1 = 1.8773731e-24
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ ijthsfwd = 0.01
+ rdsw = 100
+ toxref = 3e-9
+ aigbinv = 0.0163
+ dmcgt = 0
+ tcjsw = 0.000357
+ ijthsrev = 0.01
+ rshg = 15.6
+ bigsd = 0.00125
+ ltvoff = 2.2493116e-10
+ wvoff = 1.8056166e-9
+ poxedge = 1
+ wvsat = 0.00180338308
+ ppdiblc2 = 2.596377e-17
+ wvth0 = -3.4848103e-9
+ binunit = 2
+ pvfbsdoff = 0
+ lku0we = 2.5e-11
+ waigc = 5.3999849e-12
+ tnom = 25
+ epsrox = 3.9
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ rdsmod = 0
+ lketa = -2.0226409e-9
+ igbmod = 1
+ xpart = 1
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ egidl = 0.29734
+ pbswgd = 0.95
+ pbswgs = 0.95
+ pkvth0we = -1.3e-19
+ wags = -2.5077778e-7
+ igcmod = 1
+ wcit = -2.1754486e-10
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ voff = -0.149810363
+ acde = 0.4
+ vfbsdoff = 0.02
+ vsat = 86151.12359999999
+ wint = 0
+ vth0 = 0.379922633
+ wkt1 = 5.8978791e-9
+ wkt2 = 1.7463947e-9
+ wmax = 2.674e-7
+ aigc = 0.01161432
+ wmin = 1.08e-7
+ paramchk = 1
+ pvoff = 1.6741822e-16
+ wua1 = -2.2577864e-17
+ wub1 = 2.4820337e-26
+ wuc1 = -7.3845115e-18
+ cdscb = 0
+ cdscd = 0
+ bigc = 0.001442
+ permod = 1
+ pvsat = 8.723312000000006e-11
+ wwlc = 0
+ njtsswg = 9
+ wk2we = 5e-12
+ pvth0 = -2.6906061999999997e-16
+ drout = 0.56
+ ags = 4.0496296
+ paigc = 3.7187593e-19
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ ijthdfwd = 0.01
+ cdsc = 0
+ cjd = 0.001281008
+ cit = 0.0026629951
+ cgbo = 0
+ cjs = 0.001281008
+ clc = 1e-7
+ cle = 0.6
+ voffl = 0
+ cgdl = 3.31989e-12
+ bvd = 8.7
+ cgdo = 4.90562e-11
+ xtid = 3
+ bvs = 8.7
+ xtis = 3
+ dlc = 1.30529375e-8
+ ckappad = 0.6
+ ckappas = 0.6
+ k3b = 1.9326
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ cigc = 0.000625
+ pdiblc1 = 0
+ pdiblc2 = 0.0095469071
+ pdiblcb = -0.3
+ weta0 = 0
+ voffcv = -0.16942
+ wpemod = 1
+ lpclm = 4.8457997e-8
+ la0 = 2.768849e-7
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.004921064100000001
+ kt1 = -0.43075175
+ lk2 = -4.7065454e-9
+ kt2 = -0.10387031
+ ijthdrev = 0.01
+ llc = -1.18e-13
+ lln = 0.7
+ lu0 = -1.8130617e-10
+ mjd = 0.26
+ mjs = 0.26
+ lua = 1.2751594e-17
+ lub = -2.21968369e-26
+ cgidl = 0.22
+ luc = -7.0415723e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = -2.9632335e-14
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 4.721644e-10
+ pbs = 0.52
+ pk2 = 3.1759465e-16
+ lpdiblc2 = -9.9900678e-10
+ pu0 = 2.26802262e-18
+ bigbacc = 0.002588
+ prt = 0
+ pua = 3.9870432e-24
+ pub = -6.31495433e-33
+ puc = 2.2635812e-25
+ pud = 0
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 8.3613685e-10
+ ub1 = -6.0636714e-19
+ uc1 = 1.0129155e-10
+ tpb = 0.0014
+ wa0 = 3.1523761e-7
+ kvth0we = 0.00018
+ pbswd = 0.8
+ pbsws = 0.8
+ ute = -1
+ wat = -0.0041344832
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -2.0418175e-10
+ wlc = 0
+ wln = 1
+ wu0 = 1.5927899999999929e-12
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -4.2175679e-17
+ wub = 6.73870221e-26
+ wuc = 2.8116572e-18
+ wud = 0
+ k2we = 5e-5
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ lintnoi = -1.5e-8
+ tpbswg = 0.0009
+ dsub = 0.75
+ bigbinv = 0.004953
+ dtox = 2.7e-10
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ )

.model nch_fs_38 nmos (
+ level = 54
+ dmcgt = 0
+ poxedge = 1
+ pkvth0we = -1.3e-19
+ tcjsw = 0.000357
+ pditsd = 0
+ pditsl = 0
+ noff = 2.7195
+ cjswgd = 2.66208e-10
+ pku0we = -1.5e-18
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ cjswgs = 2.66208e-10
+ binunit = 2
+ vfbsdoff = 0.02
+ ntox = 1.0
+ pcit = -1.3274523900000001e-17
+ pclm = 2.2357699
+ bigsd = 0.00125
+ ptvfbsdoff = 0
+ mjswgd = 0.85
+ mjswgs = 0.85
+ tcjswg = 0.001
+ phin = 0.15
+ wvoff = 4.874463324000002e-9
+ paramchk = 1
+ pkt1 = -2.3945624e-15
+ pkt2 = 3.9546557e-16
+ wvsat = 0.0029164640999999984
+ wvth0 = -1.1808433999999988e-9
+ pvfbsdoff = 0
+ waigc = -1.2918923e-11
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ rbdb = 50
+ pua1 = -4.7371604e-25
+ prwb = 0
+ pub1 = -2.954512000000003e-34
+ prwg = 0
+ puc1 = -4.218097e-24
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ lketa = 2.9224258e-8
+ a0 = 0.7744856
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ ijthdfwd = 0.01
+ at = 98374.6784
+ cf = 8.15e-11
+ xpart = 1
+ ef = 1.0
+ k1 = 0.274
+ k2 = -0.044938197
+ k3 = -1.8419
+ em = 1000000.0
+ rdsw = 100
+ ll = 0
+ lw = 0
+ u0 = 0.0048412099
+ w0 = 0
+ ua = -2.6695158e-9
+ ub = 2.0926996330000003e-18
+ uc = -9.6044814e-11
+ ud = 0
+ fprout = 300
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ xrcrg1 = 12
+ xrcrg2 = 1
+ egidl = 0.29734
+ ijthdrev = 0.01
+ wtvoff = 2.7545299e-10
+ lpdiblc2 = 4.9724259e-14
+ rshg = 15.6
+ njtsswg = 9
+ capmod = 2
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ wku0we = 2e-11
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = -0.0010813536
+ mobmod = 0
+ pdiblcb = -0.3
+ ags = 4.0496296
+ pvoff = -1.2105337000000015e-16
+ cjd = 0.001281008
+ cit = 0.001090691
+ cjs = 0.001281008
+ clc = 1e-7
+ cle = 0.6
+ cdscb = 0
+ cdscd = 0
+ bvd = 8.7
+ tnom = 25
+ bvs = 8.7
+ dlc = 3.26497e-9
+ pvsat = -1.7396500000000034e-11
+ k3b = 1.9326
+ lkvth0we = -2e-12
+ wk2we = 5e-12
+ toxe = 2.43e-9
+ dwb = 0
+ dwc = 0
+ toxm = 2.43e-9
+ dwg = 0
+ dwj = 0
+ pvth0 = -4.856335000000001e-16
+ drout = 0.56
+ paigc = 2.0938533e-18
+ bigbacc = 0.002588
+ la0 = -2.5801646e-8
+ voffl = 0
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.00275118425
+ kt1 = -0.62571779
+ kt2 = -0.068117715
+ lk2 = -1.1401013e-9
+ llc = 0
+ lln = 1
+ lu0 = 2.1377612e-10
+ mjd = 0.26
+ acnqsmod = 0
+ mjs = 0.26
+ lua = 5.0500592e-17
+ lub = -3.9983527e-26
+ luc = 4.4304811e-18
+ lud = 0
+ laigsd = 1.06572e-17
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ kvth0we = 0.00018
+ weta0 = 4.2794074e-8
+ pa0 = 2.9413877e-15
+ wetab = -1.5859302e-8
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 4.1153749e-10
+ pbs = 0.52
+ pk2 = 2.316472e-16
+ lpclm = -6.2136744e-8
+ pu0 = -3.8441774999999997e-17
+ wags = -2.5077778e-7
+ prt = 0
+ pua = -3.0159915e-24
+ pub = 1.3943639e-33
+ puc = 2.394639e-25
+ pud = 0
+ lintnoi = -1.5e-8
+ rbodymod = 0
+ wcit = -4.504383699999999e-11
+ bigbinv = 0.004953
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 7.2026227e-10
+ vtsswgd = 4.2
+ ub1 = -8.074069000000001e-19
+ vtsswgs = 4.2
+ uc1 = -2.7209866e-10
+ cgidl = 0.22
+ tpb = 0.0014
+ wa0 = -3.1291358e-8
+ voff = -0.11849200800000002
+ ute = -1
+ wat = -0.00348951596
+ acde = 0.4
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 7.1015279e-10
+ wlc = 0
+ wln = 1
+ wu0 = 4.3467574000000004e-10
+ xgl = -1.09e-8
+ xgw = 0
+ wua = 3.2324691e-17
+ wub = -1.4627000299999995e-26
+ wuc = 2.6722336e-18
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ vsat = 63376.513000000006
+ wint = 0
+ vth0 = 0.24133340800000003
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ wkt1 = 2.9985826000000005e-8
+ wkt2 = -4.5976799e-9
+ wmax = 2.674e-7
+ aigc = 0.011905208
+ wmin = 1.08e-7
+ pbswd = 0.8
+ pbsws = 0.8
+ wpdiblc2 = 2.3634934e-9
+ wua1 = 5.9387403e-18
+ wub1 = -4.618226000000001e-27
+ wuc1 = 5.7460914e-17
+ pdits = 0
+ bigc = 0.001442
+ cigsd = 0.069865
+ wwlc = 0
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ cdsc = 0
+ nfactor = 1
+ toxref = 3e-9
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ wkvth0we = 2e-12
+ tnoia = 0
+ peta0 = -4.0226429e-15
+ trnqsmod = 0
+ petab = 1.4907744e-15
+ wketa = -4.815885e-9
+ tpbsw = 0.0019
+ ltvoff = 1.3417313e-10
+ nigbacc = 10
+ tvfbsdoff = 0.022
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ cjswd = 7.7408e-11
+ cjsws = 7.7408e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ k2we = 5e-5
+ nigbinv = 10
+ dsub = 0.75
+ rgatemod = 0
+ lku0we = 2.5e-11
+ dtox = 2.7e-10
+ tnjtsswg = 1
+ epsrox = 3.9
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ rdsmod = 0
+ eta0 = -0.13238438
+ etab = 0.18670848
+ igbmod = 1
+ scref = 1e-6
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ pigcd = 2.621
+ aigsd = 0.010772573
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ fnoimod = 1
+ pbswgd = 0.95
+ pbswgs = 0.95
+ eigbinv = 1.1
+ lvoff = -2.8954111999999996e-9
+ igcmod = 1
+ lvsat = 0.0015515391499999998
+ lvth0 = 4.6854495e-9
+ delta = 0.007595625
+ laigc = -3.4086068e-11
+ rnoia = 0
+ rnoib = 0
+ pketa = -3.9657201e-16
+ ngate = 8e+20
+ paigsd = -2.9413875e-24
+ ngcon = 1
+ cigbacc = 0.32875
+ wpclm = -8.3073835e-8
+ gbmin = 1e-12
+ tnoimod = 0
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ permod = 1
+ cigbinv = 0.006
+ ijthsfwd = 0.01
+ voffcv = -0.16942
+ wpemod = 1
+ version = 4.5
+ keta = -0.45164428
+ tempmod = 0
+ ijthsrev = 0.01
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 1.004633e-10
+ tvoff = -0.0018736893
+ aigbacc = 0.02
+ kt1l = 0
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ lint = 0
+ lkt1 = 1.8405602e-8
+ lkt2 = -3.1935983e-9
+ lmax = 9e-8
+ lmin = 5.4e-8
+ tpbswg = 0.0009
+ ku0we = -0.0007
+ aigbinv = 0.0163
+ beta0 = 13
+ lpe0 = 9.2e-8
+ ppdiblc2 = -1.2574432e-20
+ lpeb = 2.5e-7
+ leta0 = 3.2844132e-8
+ letab = -3.6350598e-8
+ wtvfbsdoff = 0
+ minv = -0.3
+ ppclm = 2.1858187e-15
+ lua1 = 4.1554342e-18
+ lub1 = -2.1863483e-26
+ luc1 = 2.4128073e-17
+ ndep = 1e+18
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ ptvoff = -2.2148869e-17
+ lwlc = 0
+ moin = 5.1
+ ltvfbsdoff = 0
+ waigsd = 3.1789053e-12
+ nigc = 3.083
+ diomod = 1
+ )

.model nch_fs_39 nmos (
+ level = 54
+ wkt1 = -2.8322054999999998e-8
+ wkt2 = 1.1625249e-8
+ wmax = 2.674e-7
+ aigc = 0.011615807
+ wmin = 1.08e-7
+ fnoimod = 1
+ eigbinv = 1.1
+ wua1 = -1.0774777e-16
+ wub1 = 1.2771999e-25
+ wuc1 = 1.606153e-17
+ bigc = 0.001442
+ wwlc = 0
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ scref = 1e-6
+ ijthsfwd = 0.01
+ cdsc = 0
+ fprout = 300
+ pigcd = 2.621
+ cgbo = 0
+ aigsd = 0.010772573
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ xrcrg1 = 12
+ xrcrg2 = 1
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ lvoff = -6.504439899999998e-9
+ cigbacc = 0.32875
+ lvsat = -0.0024565101
+ wtvoff = 7.91509e-11
+ lvth0 = 7.430732700000001e-9
+ ijthsrev = 0.01
+ tnoimod = 0
+ delta = 0.007595625
+ laigc = -1.730084e-11
+ rnoia = 0
+ rnoib = 0
+ cigbinv = 0.006
+ dmcg = 3.1e-8
+ capmod = 2
+ dmci = 3.1e-8
+ dmdg = 0
+ wku0we = 2e-11
+ pketa = 1.224516e-15
+ ngate = 8e+20
+ a0 = 19.191807
+ a1 = 0
+ a2 = 1
+ ngcon = 1
+ b0 = 0
+ b1 = 0
+ mobmod = 0
+ wpclm = -5.2664346e-8
+ at = 83923.56199999999
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = -0.059313829
+ k3 = -1.8419
+ em = 1000000.0
+ k2we = 5e-5
+ ll = 0
+ lw = 0
+ u0 = 0.0018707365
+ w0 = 0
+ ua = -2.3710013e-9
+ ub = 1.4550579529999998e-18
+ uc = -1.4785261e-10
+ ud = 0
+ version = 4.5
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ dsub = 0.75
+ dtox = 2.7e-10
+ gbmin = 1e-12
+ tempmod = 0
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ eta0 = 1.1504337
+ aigbacc = 0.02
+ etab = -1.3364008
+ pkvth0we = -1.3e-19
+ aigbinv = 0.0163
+ tvoff = -0.0045522389
+ vfbsdoff = 0.02
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ paramchk = 1
+ ku0we = -0.0007
+ beta0 = 13
+ leta0 = -4.1559315e-8
+ poxedge = 1
+ letab = 5.198974e-8
+ ppclm = 4.2206835e-16
+ binunit = 2
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ ijthdfwd = 0.01
+ toxref = 3e-9
+ dmcgt = 0
+ keta = 0.16119603
+ tcjsw = 0.000357
+ ijthdrev = 0.01
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 4.5379023e-10
+ ltvoff = 2.8952901e-10
+ kt1l = 0
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ bigsd = 0.00125
+ lint = 0
+ wvoff = -2.2288246e-9
+ lkt1 = 3.267505000000001e-9
+ lkt2 = 8.1983323e-9
+ lmax = 5.4e-8
+ lmin = 4.5e-8
+ wvsat = -0.0033283578000000017
+ lku0we = 2.5e-11
+ pvfbsdoff = 0
+ lpe0 = 9.2e-8
+ wvth0 = -6.322442099999999e-9
+ lpeb = 2.5e-7
+ epsrox = 3.9
+ waigc = 4.0939876e-11
+ minv = -0.3
+ lua1 = -3.9796071e-17
+ lub1 = 4.2129051e-26
+ luc1 = 1.4911728e-19
+ rdsmod = 0
+ lkvth0we = -2e-12
+ ndep = 1e+18
+ igbmod = 1
+ lwlc = 0
+ lketa = -6.3204807e-9
+ moin = 5.1
+ njtsswg = 9
+ xpart = 1
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ nigc = 3.083
+ pbswgd = 0.95
+ pbswgs = 0.95
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ acnqsmod = 0
+ egidl = 0.29734
+ igcmod = 1
+ ckappad = 0.6
+ ckappas = 0.6
+ noff = 2.7195
+ pdiblc1 = 0
+ pdiblc2 = -0.0010804963
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ pdiblcb = -0.3
+ rbodymod = 0
+ ntox = 1.0
+ pcit = -3.3822647e-17
+ pclm = 1.0542662
+ ags = 4.0496296
+ bigbacc = 0.002588
+ phin = 0.15
+ cjd = 0.001281008
+ cit = -0.0050011527
+ cjs = 0.001281008
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 3.26497e-9
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ pkt1 = 9.872907599999998e-16
+ pkt2 = -5.454643e-16
+ dwg = 0
+ dwj = 0
+ kvth0we = 0.00018
+ wpdiblc2 = 2.3632766e-9
+ permod = 1
+ pvoff = 2.9093734999999984e-16
+ lintnoi = -1.5e-8
+ la0 = -1.0940063e-6
+ cdscb = 0
+ cdscd = 0
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.0019130205800000008
+ bigbinv = 0.004953
+ kt1 = -0.36471641
+ kt2 = -0.26453031
+ lk2 = -3.0631458e-10
+ vtsswgd = 4.2
+ pvsat = 3.4480318e-10
+ vtsswgs = 4.2
+ llc = 0
+ lln = 1
+ lu0 = 3.8606358e-10
+ wk2we = 5e-12
+ pvth0 = -1.8742074599999998e-16
+ mjd = 0.26
+ mjs = 0.26
+ lua = 3.3186753e-17
+ lub = -3.0003129999999985e-27
+ luc = 7.435334e-18
+ lud = 0
+ rbdb = 50
+ pua1 = 6.1201017e-24
+ prwb = 0
+ lwc = 0
+ pub1 = -7.9710719e-33
+ prwg = 0
+ drout = 0.56
+ lwl = 0
+ puc1 = -1.8169327e-24
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 1.2471671e-13
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ nsd = 1e+20
+ pvag = 1.2
+ pbd = 0.52
+ pat = -1.8302546000000003e-10
+ pbs = 0.52
+ pk2 = 1.8168527e-16
+ paigc = -1.0299571e-18
+ pu0 = -8.066070399999998e-18
+ prt = 0
+ pua = 6.5377716e-24
+ pub = -1.101976303e-32
+ rdsw = 100
+ puc = -3.076481e-25
+ pud = 0
+ voffl = 0
+ rsh = 17.5
+ tcj = 0.00076
+ voffcv = -0.16942
+ wpemod = 1
+ ua1 = 1.4780468e-9
+ ub1 = -1.9107259e-18
+ uc1 = 1.4133161e-10
+ tpb = 0.0014
+ wa0 = -2.130866e-6
+ weta0 = -1.5669611e-7
+ ute = -1
+ wetab = 4.0317659e-8
+ wat = 0.006761574299999999
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 1.5715655e-9
+ wlc = 0
+ wln = 1
+ wu0 = -8.904329700000001e-11
+ lpclm = 6.3904735e-9
+ xgl = -1.09e-8
+ wkvth0we = 2e-12
+ xgw = 0
+ wua = -1.3239536e-16
+ wub = 1.9940967600000001e-25
+ wuc = 1.2105201e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ cgidl = 0.22
+ trnqsmod = 0
+ rshg = 15.6
+ wtvfbsdoff = 0
+ nfactor = 1
+ pbswd = 0.8
+ pbsws = 0.8
+ tpbswg = 0.0009
+ ltvfbsdoff = 0
+ rgatemod = 0
+ tnjtsswg = 1
+ pdits = 0
+ tnom = 25
+ cigsd = 0.069865
+ toxe = 2.43e-9
+ ptvoff = -1.0763348e-17
+ toxm = 2.43e-9
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ waigsd = 3.1788545e-12
+ nigbacc = 10
+ pk2we = -1e-19
+ diomod = 1
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ ptvfbsdoff = 0
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 2.66208e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.66208e-10
+ wags = -2.5077778e-7
+ tnoia = 0
+ nigbinv = 10
+ wcit = 3.0923414e-10
+ peta0 = 7.5477876e-15
+ petab = -1.7674893e-15
+ voff = -0.056267378999999965
+ wketa = -3.2765679e-8
+ acde = 0.4
+ tvfbsdoff = 0.022
+ tpbsw = 0.0019
+ mjswgd = 0.85
+ mjswgs = 0.85
+ vsat = 132480.81299999997
+ wint = 0
+ cjswd = 7.7408e-11
+ cjsws = 7.7408e-11
+ vth0 = 0.19400093900000004
+ tcjswg = 0.001
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ )

.model nch_fs_40 nmos (
+ level = 54
+ wkt1 = 2.9249329999999966e-9
+ wkt2 = -1.1473225e-8
+ wmax = 2.674e-7
+ aigc = 0.011144932
+ wmin = 1.08e-7
+ fnoimod = 1
+ eigbinv = 1.1
+ wua1 = 1.9140234e-16
+ wub1 = -2.914296e-25
+ wuc1 = -2.3798265000000004e-17
+ bigc = 0.001442
+ wwlc = 0
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ scref = 1e-6
+ ijthsfwd = 0.01
+ cdsc = 0
+ fprout = 300
+ pigcd = 2.621
+ cgbo = 0
+ aigsd = 0.010772574
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ xrcrg1 = 12
+ xrcrg2 = 1
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ lvoff = -7.122739300000001e-9
+ cigbacc = 0.32875
+ lvsat = 0.0054477623200000005
+ wtvoff = -7.2128996e-10
+ lvth0 = -4.5987852e-9
+ ijthsrev = 0.01
+ tnoimod = 0
+ delta = 0.007595625
+ laigc = 5.7720314e-12
+ rnoia = 0
+ rnoib = 0
+ cigbinv = 0.006
+ dmcg = 3.1e-8
+ capmod = 2
+ dmci = 3.1e-8
+ dmdg = 0
+ wku0we = 2e-11
+ pketa = -8.4677334e-15
+ ngate = 8e+20
+ a0 = -5.925916599999999
+ a1 = 0
+ a2 = 1
+ ngcon = 1
+ b0 = 0
+ b1 = 0
+ mobmod = 0
+ wpclm = -7.2101286e-7
+ at = 102879.242
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.013923130999999998
+ k3 = -1.8419
+ em = 1000000.0
+ k2we = 5e-5
+ ll = 0
+ lw = 0
+ u0 = 0.012408487999999999
+ w0 = 0
+ ua = -5.589164400000002e-10
+ ub = 8.937269600000036e-20
+ uc = 2.381934e-10
+ ud = 0
+ version = 4.5
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ dsub = 0.75
+ dtox = 2.7e-10
+ gbmin = 1e-12
+ tempmod = 0
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ eta0 = -0.288265897
+ aigbacc = 0.02
+ etab = -0.74723747
+ laigsd = -1.5325105e-17
+ pkvth0we = -1.3e-19
+ aigbinv = 0.0163
+ tvoff = 0.0062987975
+ vfbsdoff = 0.02
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ paramchk = 1
+ ku0we = -0.0007
+ beta0 = 13
+ leta0 = 2.8936964e-8
+ poxedge = 1
+ letab = 2.3120738e-8
+ ppclm = 3.3171145e-14
+ binunit = 2
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ ijthdfwd = 0.01
+ toxref = 3e-9
+ dmcgt = 0
+ keta = -0.51478944
+ tcjsw = 0.000357
+ ijthdrev = 0.01
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 2.322945e-10
+ ltvoff = -2.4217179e-10
+ kt1l = 0
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ bigsd = 0.00125
+ lint = 0
+ wvoff = 1.3282831000000013e-9
+ lkt1 = 2.6234833e-9
+ lkt2 = -1.1864945e-9
+ lmax = 4.5e-8
+ lmin = 3.6e-8
+ wvsat = 0.020304221399999996
+ lku0we = 2.5e-11
+ pvfbsdoff = 0
+ lpe0 = 9.2e-8
+ wvth0 = -3.1680437e-8
+ lpeb = 2.5e-7
+ epsrox = 3.9
+ waigc = 5.1623453e-11
+ minv = -0.3
+ lua1 = 6.0050187e-18
+ lub1 = -1.38723653e-26
+ luc1 = 6.4275095e-18
+ rdsmod = 0
+ lkvth0we = -2e-12
+ ndep = 1e+18
+ igbmod = 1
+ lwlc = 0
+ lketa = 2.6802806000000003e-8
+ moin = 5.1
+ njtsswg = 9
+ xpart = 1
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ nigc = 3.083
+ pbswgd = 0.95
+ pbswgs = 0.95
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ acnqsmod = 0
+ egidl = 0.29734
+ igcmod = 1
+ ckappad = 0.6
+ ckappas = 0.6
+ noff = 2.7195
+ pdiblc1 = 0
+ pdiblc2 = -0.0010804963
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ pdiblcb = -0.3
+ rbodymod = 0
+ ntox = 1.0
+ pcit = 6.683632e-17
+ pclm = 4.6708343
+ ags = 4.0496296
+ bigbacc = 0.002588
+ phin = 0.15
+ paigsd = 4.2297301e-24
+ cjd = 0.001281008
+ cit = -0.0004808017000000001
+ cjs = 0.001281008
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 3.26497e-9
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ pkt1 = -5.438076399999999e-16
+ pkt2 = 5.863609e-16
+ dwg = 0
+ dwj = 0
+ kvth0we = 0.00018
+ wpdiblc2 = 2.3632766e-9
+ permod = 1
+ pvoff = 1.1663916e-16
+ lintnoi = -1.5e-8
+ la0 = 1.3676219000000002e-7
+ cdscb = 0
+ cdscd = 0
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.0028418533199999997
+ bigbinv = 0.004953
+ kt1 = -0.35157258
+ kt2 = -0.073003235
+ lk2 = -3.894925700000001e-9
+ vtsswgd = 4.2
+ pvsat = -8.1319336e-10
+ vtsswgs = 4.2
+ llc = 0
+ lln = 1
+ lu0 = -1.3028556e-10
+ wk2we = 5e-12
+ pvth0 = 1.05512139e-15
+ mjd = 0.26
+ mjs = 0.26
+ lua = -5.56054081e-17
+ lub = 6.391826569999999e-26
+ luc = -1.14809219e-17
+ lud = 0
+ rbdb = 50
+ pua1 = -8.5382538e-24
+ prwb = 0
+ lwc = 0
+ pub1 = 1.2567259000000002e-32
+ prwg = 0
+ drout = 0.56
+ lwl = 0
+ puc1 = 1.361972e-25
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = -7.5523402e-14
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ nsd = 1e+20
+ pvag = 1.2
+ pbd = 0.52
+ pat = 2.6945479999999945e-11
+ pbs = 0.52
+ pk2 = 5.0756697e-16
+ paigc = -1.5534524e-18
+ pu0 = 1.02148438e-17
+ prt = 0
+ pua = -2.8276596999999977e-25
+ pub = -6.331388000000253e-35
+ rdsw = 100
+ puc = 4.398917e-25
+ pud = 0
+ voffl = 0
+ rsh = 17.5
+ tcj = 0.00076
+ voffcv = -0.16942
+ wpemod = 1
+ ua1 = 5.4333072e-10
+ ub1 = -7.678405400000001e-19
+ uc1 = 1.3201149999999995e-11
+ tpb = 0.0014
+ wa0 = 1.9556670799999998e-6
+ weta0 = 9.4960797e-8
+ ute = -1
+ wetab = 3.9258957e-9
+ wat = 0.0024764724999999993
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -5.0790816e-9
+ wlc = 0
+ wln = 1
+ wu0 = -4.6212356999999993e-10
+ lpclm = -1.70821362e-7
+ xgl = -1.09e-8
+ wkvth0we = 2e-12
+ xgw = 0
+ wua = 6.799270000000015e-18
+ wub = -2.4191335000000008e-26
+ wuc = -3.150715e-18
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ cgidl = 0.22
+ trnqsmod = 0
+ rshg = 15.6
+ wtvfbsdoff = 0
+ nfactor = 1
+ pbswd = 0.8
+ pbsws = 0.8
+ tpbswg = 0.0009
+ ltvfbsdoff = 0
+ rgatemod = 0
+ tnjtsswg = 1
+ pdits = 0
+ tnom = 25
+ cigsd = 0.069865
+ toxe = 2.43e-9
+ ptvoff = 2.8458255e-17
+ toxm = 2.43e-9
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ waigsd = 3.1787682e-12
+ nigbacc = 10
+ pk2we = -1e-19
+ diomod = 1
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ ptvfbsdoff = 0
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 2.66208e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.66208e-10
+ wags = -2.5077778e-7
+ tnoia = 0
+ nigbinv = 10
+ wcit = -1.74502578e-9
+ peta0 = -4.7834008e-15
+ petab = 1.5707054e-17
+ voff = -0.043649036000000016
+ wketa = 1.65035329e-7
+ acde = 0.4
+ tvfbsdoff = 0.022
+ tpbsw = 0.0019
+ mjswgd = 0.85
+ mjswgs = 0.85
+ vsat = -28830.753999999986
+ wint = 0
+ cjswd = 7.7408e-11
+ cjsws = 7.7408e-11
+ vth0 = 0.439501247
+ tcjswg = 0.001
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ )

.model nch_sf_1 nmos (
+ level = 54
+ fprout = 300
+ xrcrg1 = 12
+ xrcrg2 = 1
+ ags = 0.9475
+ wtvoff = 0
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ tvoff = 0.0019109629
+ keta = -0.06
+ cjd = 0.001432992
+ cit = 0.0001
+ cjs = 0.001432992
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 9.8024918e-9
+ xjbvd = 1
+ k3b = 1.9326
+ xjbvs = 1
+ lk2we = -1.5e-12
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ tvfbsdoff = 0.022
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 8e-12
+ capmod = 2
+ la0 = 0
+ kt1l = 0
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = 8e-5
+ kt1 = -0.200226
+ kt2 = -0.05325
+ wku0we = 2e-11
+ wkvth0we = 2e-12
+ llc = 0
+ ku0we = -0.0007
+ lln = 1
+ lu0 = -4e-12
+ mjd = 0.26
+ mjs = 0.26
+ beta0 = 13
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ leta0 = -1.6000000000000003e-9
+ njs = 1.02
+ pa0 = 0
+ mobmod = 0
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 1.44e-11
+ pbs = 0.52
+ lint = 6.5375218e-9
+ trnqsmod = 0
+ pu0 = -1.2e-18
+ prt = 0
+ pud = 0
+ lkt1 = -2.4e-10
+ lmax = 2.001e-5
+ lmin = 8.9991e-6
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 1.2299687e-9
+ ub1 = -7.2455506e-19
+ uc1 = 3.028e-11
+ dlcig = 2.5e-9
+ tpb = 0.0014
+ lpe0 = 9.2e-8
+ njtsswg = 9
+ bgidl = 2320000000.0
+ lpeb = 2.5e-7
+ wa0 = 0
+ ute = -1.007
+ wat = 0
+ web = 6843.8
+ wec = -25529.0
+ wlc = 0
+ wln = 1
+ wu0 = 3.6000000000000005e-11
+ xgl = -1.09e-8
+ xgw = 0
+ wud = 0
+ wwc = 0
+ minv = -0.3
+ wwl = 0
+ wwn = 1
+ xtsswgd = 0.18
+ wvfbsdoff = 0
+ xtsswgs = 0.18
+ lvfbsdoff = 0
+ lub1 = 2.4000000000000004e-27
+ ndep = 1e+18
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.018555248
+ lwlc = 0
+ rgatemod = 0
+ dmcgt = 0
+ pdiblcb = -0.3
+ moin = 5.1
+ tcjsw = 0.000357
+ tnjtsswg = 1
+ nigc = 3.083
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ bigsd = 0.00125
+ bigbacc = 0.002588
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ wvoff = -3.2000000000000003e-10
+ ntox = 1.0
+ pcit = 1.2000000000000001e-17
+ kvth0we = 0.00018
+ pclm = 1.4
+ wvsat = 0
+ wvth0 = 2.4e-9
+ lintnoi = -1.5e-8
+ bigbinv = 0.004953
+ phin = 0.15
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ pkt1 = -1.76e-16
+ a0 = 3.25
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 72000
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.026201254
+ k3 = -1.8419
+ em = 1000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.01599
+ w0 = 0
+ ua = -1.8237726e-9
+ ub = 2.103696e-18
+ xpart = 1
+ uc = 7.33e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 3.4e-9
+ toxref = 3e-9
+ rbdb = 50
+ prwb = 0
+ prwg = 0
+ pub1 = 1.6e-34
+ egidl = 0.29734
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ rdsw = 100
+ ijthsfwd = 0.01
+ ltvoff = 0
+ nfactor = 1
+ rshg = 15.6
+ ijthsrev = 0.01
+ pvoff = -4e-17
+ lku0we = 2.5e-11
+ cdscb = 0
+ cdscd = 0
+ epsrox = 3.9
+ pvsat = 1.44e-11
+ wk2we = 5e-12
+ pvth0 = 1.2e-16
+ drout = 0.56
+ nigbacc = 10
+ rdsmod = 0
+ igbmod = 1
+ voffl = 0
+ tnom = 25
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ weta0 = 0
+ pbswgd = 0.95
+ pbswgs = 0.95
+ nigbinv = 10
+ igcmod = 1
+ cgidl = 0.22
+ wags = 8e-9
+ wcit = -4.0000000000000004e-11
+ voff = -0.1128204
+ fnoimod = 1
+ pbswd = 0.8
+ pbsws = 0.8
+ acde = 0.4
+ pkvth0we = -1.3e-19
+ eigbinv = 1.1
+ vsat = 102860
+ wint = 0
+ vth0 = 0.37631089
+ wkt1 = 2.5600000000000003e-9
+ pvfbsdoff = 0
+ wmax = 0.00090001
+ aigc = 0.011769394
+ wmin = 9.0026e-6
+ pdits = 0
+ vfbsdoff = 0.02
+ permod = 1
+ cigsd = 0.069865
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ bigc = 0.001442
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ paramchk = 1
+ wwlc = 0
+ cigbacc = 0.32875
+ voffcv = -0.16942
+ wpemod = 1
+ cdsc = 0
+ tnoia = 0
+ tnoimod = 0
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ peta0 = 0.0
+ cigbinv = 0.006
+ tpbsw = 0.0019
+ ijthdfwd = 0.01
+ cjswd = 8.6592e-11
+ cjsws = 8.6592e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ version = 4.5
+ tempmod = 0
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ tpbswg = 0.0009
+ ijthdrev = 0.01
+ aigbacc = 0.02
+ k2we = 5e-5
+ dsub = 0.75
+ dtox = 2.7e-10
+ scref = 1e-6
+ ptvoff = 0
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ pigcd = 2.621
+ aigsd = 0.01077322
+ lvoff = 1.6e-11
+ eta0 = 0.3
+ aigbinv = 0.0163
+ diomod = 1
+ etab = -0.25
+ wtvfbsdoff = 0
+ lvsat = 0.00016
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 2.9779200000000003e-10
+ pku0we = -1.5e-18
+ lvth0 = 4.0000000000000007e-10
+ cjswgs = 2.9779200000000003e-10
+ lkvth0we = -2e-12
+ delta = 0.007595625
+ ltvfbsdoff = 0
+ rnoia = 0
+ rnoib = 0
+ mjswgd = 0.85
+ mjswgs = 0.85
+ acnqsmod = 0
+ ngate = 8e+20
+ tcjswg = 0.001
+ ngcon = 1
+ poxedge = 1
+ rbodymod = 0
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ binunit = 2
+ ptvfbsdoff = 0
+ )

.model nch_sf_2 nmos (
+ level = 54
+ wtvoff = 0
+ cgidl = 0.22
+ ijthdfwd = 0.01
+ capmod = 2
+ pbswd = 0.8
+ pbsws = 0.8
+ wku0we = 2e-11
+ rshg = 15.6
+ cigbacc = 0.32875
+ mobmod = 0
+ pvfbsdoff = 0
+ ijthdrev = 0.01
+ tnoimod = 0
+ pdits = 0
+ lpdiblc2 = -5.8501673e-10
+ cigsd = 0.069865
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ cigbinv = 0.006
+ tnom = 25
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ version = 4.5
+ tnoia = 0
+ tempmod = 0
+ lkvth0we = -2e-12
+ peta0 = 0.0
+ tpbsw = 0.0019
+ aigbacc = 0.02
+ wags = 8e-9
+ cjswd = 8.6592e-11
+ cjsws = 8.6592e-11
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ wcit = -4.0000000000000004e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ acnqsmod = 0
+ voff = -0.11120139
+ acde = 0.4
+ vsat = 102860
+ wint = 0
+ rbodymod = 0
+ aigbinv = 0.0163
+ vth0 = 0.37056703
+ wkt1 = 2.5600000000000003e-9
+ wmax = 0.00090001
+ aigc = 0.01178613
+ wmin = 9.0026e-6
+ scref = 1e-6
+ pigcd = 2.621
+ toxref = 3e-9
+ aigsd = 0.01077322
+ bigc = 0.001442
+ wwlc = 0
+ lvoff = -1.4538874e-8
+ poxedge = 1
+ cdsc = 0
+ lvsat = 0.00016
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ lvth0 = 5.2037332e-8
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ delta = 0.007595625
+ binunit = 2
+ laigc = -1.5044982e-10
+ rnoia = 0
+ rnoib = 0
+ ltvoff = -1.4627394e-10
+ a0 = 3.4752469
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ ngate = 8e+20
+ at = 61592.494
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.027688843
+ k3 = -1.8419
+ em = 1000000.0
+ ngcon = 1
+ ll = 0
+ lw = 0
+ u0 = 0.016211951000000002
+ w0 = 0
+ ua = -1.7995884e-9
+ ub = 2.1046515e-18
+ uc = 7.3387901e-11
+ ud = 0
+ wkvth0we = 2e-12
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 3.4e-9
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ lku0we = 2.5e-11
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ trnqsmod = 0
+ epsrox = 3.9
+ k2we = 5e-5
+ rdsmod = 0
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ dsub = 0.75
+ dtox = 2.7e-10
+ igbmod = 1
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ ags = 0.95104901
+ pbswgd = 0.95
+ pbswgs = 0.95
+ eta0 = 0.3
+ cjd = 0.001432992
+ rgatemod = 0
+ etab = -0.25
+ cit = -2.3830864e-5
+ cjs = 0.001432992
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 9.8024918e-9
+ tnjtsswg = 1
+ k3b = 1.9326
+ igcmod = 1
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ tvoff = 0.0019272336
+ la0 = -2.0249698e-6
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = 0.093643481
+ kt1 = -0.19577666
+ lk2 = -1.337342e-8
+ kt2 = -0.051823539
+ xjbvd = 1
+ llc = 0
+ xjbvs = 1
+ lln = 1
+ tvfbsdoff = 0.022
+ lk2we = -1.5e-12
+ lu0 = -1.9993361e-9
+ mjd = 0.26
+ lua = -2.1741579e-16
+ mjs = 0.26
+ lub = -8.5898229e-27
+ luc = -7.902321e-19
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njtsswg = 9
+ njd = 1.02
+ njs = 1.02
+ pa0 = 0
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 1.44e-11
+ pbs = 0.52
+ pu0 = -1.2e-18
+ xtsswgd = 0.18
+ prt = 0
+ pud = 0
+ xtsswgs = 0.18
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 1.2713861e-9
+ ub1 = -7.4616446e-19
+ ku0we = -0.0007
+ uc1 = 2.5703642e-11
+ ckappad = 0.6
+ ckappas = 0.6
+ beta0 = 13
+ tpb = 0.0014
+ wa0 = 0
+ leta0 = -1.6000000000000003e-9
+ pdiblc1 = 0
+ pdiblc2 = 0.018620322
+ pdiblcb = -0.3
+ ute = -1.0077691
+ wat = 0
+ web = 6843.8
+ wec = -25529.0
+ wlc = 0
+ wln = 1
+ wu0 = 3.6000000000000005e-11
+ xgl = -1.09e-8
+ xgw = 0
+ permod = 1
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ bigbacc = 0.002588
+ voffcv = -0.16942
+ wpemod = 1
+ dmcgt = 0
+ tcjsw = 0.000357
+ kvth0we = 0.00018
+ lintnoi = -1.5e-8
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ keta = -0.059896633
+ ijthsfwd = 0.01
+ bigsd = 0.00125
+ lags = -3.1905621e-8
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 1.1212395e-9
+ wvoff = -3.2000000000000003e-10
+ kt1l = 0
+ tpbswg = 0.0009
+ wvsat = 0
+ wvth0 = 2.4e-9
+ ijthsrev = 0.01
+ lint = 6.5375218e-9
+ lkt1 = -4.0239573e-8
+ lkt2 = -1.2823887e-8
+ wtvfbsdoff = 0
+ lmax = 8.9991e-6
+ lmin = 8.9908e-7
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ ptvoff = 0
+ lketa = -9.2926692e-10
+ xpart = 1
+ ltvfbsdoff = 0
+ minv = -0.3
+ lua1 = -3.7234224e-16
+ lub1 = 1.9666850999999998e-25
+ luc1 = 4.1141459e-17
+ nfactor = 1
+ diomod = 1
+ ndep = 1e+18
+ lute = 6.9145309e-9
+ egidl = 0.29734
+ lwlc = 0
+ moin = 5.1
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 2.9779200000000003e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.9779200000000003e-10
+ nigc = 3.083
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ mjswgd = 0.85
+ mjswgs = 0.85
+ nigbacc = 10
+ ptvfbsdoff = 0
+ tcjswg = 0.001
+ ntox = 1.0
+ pkvth0we = -1.3e-19
+ pcit = 1.2000000000000001e-17
+ pclm = 1.4
+ pvoff = -4e-17
+ nigbinv = 10
+ phin = 0.15
+ cdscb = 0
+ cdscd = 0
+ vfbsdoff = 0.02
+ pvsat = 1.44e-11
+ wk2we = 5e-12
+ pkt1 = -1.76e-16
+ pvth0 = 1.2e-16
+ drout = 0.56
+ voffl = 0
+ fprout = 300
+ paramchk = 1
+ rbdb = 50
+ prwb = 0
+ prwg = 0
+ pub1 = 1.6e-34
+ xrcrg1 = 12
+ xrcrg2 = 1
+ fnoimod = 1
+ weta0 = 0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ eigbinv = 1.1
+ rdsw = 100
+ )

.model nch_sf_3 nmos (
+ level = 54
+ ku0we = -0.0007
+ beta0 = 13
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ leta0 = -1.6000000000000003e-9
+ ijthsrev = 0.01
+ kvth0we = 0.00018
+ lintnoi = -1.5e-8
+ k2we = 5e-5
+ bigbinv = 0.004953
+ dlcig = 2.5e-9
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ bgidl = 2320000000.0
+ dsub = 0.75
+ wvfbsdoff = 0
+ dtox = 2.7e-10
+ lvfbsdoff = 0
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ eta0 = 0.3
+ dmcgt = 0
+ etab = -0.25
+ tcjsw = 0.000357
+ bigsd = 0.00125
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ wvoff = -3.2000000000000003e-10
+ pkvth0we = -1.3e-19
+ nfactor = 1
+ wvsat = 0
+ wvth0 = 2.4e-9
+ vfbsdoff = 0.02
+ lketa = -2.6515603e-8
+ toxref = 3e-9
+ xpart = 1
+ nigbacc = 10
+ paramchk = 1
+ egidl = 0.29734
+ nigbinv = 10
+ keta = -0.031147941
+ ltvoff = -6.4393769e-10
+ ijthdfwd = 0.01
+ lags = 4.0889306e-7
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = -1.0251822e-10
+ kt1l = 0
+ lku0we = 2.5e-11
+ fnoimod = 1
+ ijthdrev = 0.01
+ epsrox = 3.9
+ eigbinv = 1.1
+ pvoff = -4e-17
+ lint = 6.5375218e-9
+ cdscb = 0
+ cdscd = 0
+ lkt1 = -1.8004368000000002e-8
+ lkt2 = -1.1493547e-8
+ lmax = 8.9908e-7
+ lpdiblc2 = 3.0380287e-9
+ pvsat = 1.44e-11
+ lmin = 4.4908e-7
+ rdsmod = 0
+ wk2we = 5e-12
+ pvth0 = 1.2e-16
+ drout = 0.56
+ igbmod = 1
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ minv = -0.3
+ voffl = 0
+ lua1 = -1.0281867e-16
+ lub1 = 2.0952992e-26
+ luc1 = 3.7680622e-18
+ pbswgd = 0.95
+ pbswgs = 0.95
+ ndep = 1e+18
+ weta0 = 0
+ lwlc = 0
+ igcmod = 1
+ moin = 5.1
+ a0 = 1.288
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ cigbacc = 0.32875
+ at = 219598.22
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.026610322000000002
+ k3 = -1.8419
+ em = 1000000.0
+ ll = 0
+ nigc = 3.083
+ lw = 0
+ u0 = 0.015710444
+ w0 = 0
+ ua = -1.9429424e-9
+ ub = 2.1566e-18
+ uc = 9.3717778e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 3.4e-9
+ lkvth0we = -2e-12
+ cgidl = 0.22
+ tnoimod = 0
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ cigbinv = 0.006
+ acnqsmod = 0
+ pbswd = 0.8
+ pbsws = 0.8
+ ntox = 1.0
+ pcit = 1.2000000000000001e-17
+ pclm = 1.4
+ pvfbsdoff = 0
+ rbodymod = 0
+ version = 4.5
+ permod = 1
+ phin = 0.15
+ tempmod = 0
+ pdits = 0
+ cigsd = 0.069865
+ pkt1 = -1.76e-16
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ aigbacc = 0.02
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ voffcv = -0.16942
+ wpemod = 1
+ rbdb = 50
+ prwb = 0
+ pub1 = 1.6e-34
+ prwg = 0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ tnoia = 0
+ rdsw = 100
+ aigbinv = 0.0163
+ peta0 = 0.0
+ tpbsw = 0.0019
+ wtvfbsdoff = 0
+ cjswd = 8.6592e-11
+ cjsws = 8.6592e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ tpbswg = 0.0009
+ rshg = 15.6
+ ltvfbsdoff = 0
+ wkvth0we = 2e-12
+ poxedge = 1
+ trnqsmod = 0
+ ptvoff = 0
+ binunit = 2
+ scref = 1e-6
+ pigcd = 2.621
+ aigsd = 0.01077322
+ tnom = 25
+ diomod = 1
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ ptvfbsdoff = 0
+ lvoff = -1.3752912000000001e-8
+ pditsd = 0
+ rgatemod = 0
+ pditsl = 0
+ cjswgd = 2.9779200000000003e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.9779200000000003e-10
+ tnjtsswg = 1
+ lvsat = 0.00016
+ lvth0 = 7.8115504e-9
+ delta = 0.007595625
+ laigc = -5.5724245e-11
+ rnoia = 0
+ rnoib = 0
+ mjswgd = 0.85
+ mjswgs = 0.85
+ wags = 8e-9
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ wcit = -4.0000000000000004e-11
+ tcjswg = 0.001
+ ngate = 8e+20
+ voff = -0.1120845
+ acde = 0.4
+ ngcon = 1
+ vsat = 102860
+ wint = 0
+ vth0 = 0.42025892
+ gbmin = 1e-12
+ wkt1 = 2.5600000000000003e-9
+ jswgd = 1.28e-13
+ wmax = 0.00090001
+ jswgs = 1.28e-13
+ aigc = 0.011679696
+ wmin = 9.0026e-6
+ ags = 0.4557696
+ cjd = 0.001432992
+ cit = 0.0013511778
+ cjs = 0.001432992
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 9.8024918e-9
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ fprout = 300
+ dwg = 0
+ dwj = 0
+ njtsswg = 9
+ bigc = 0.001442
+ xrcrg1 = 12
+ xrcrg2 = 1
+ wwlc = 0
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ la0 = -7.832e-8
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.046981618
+ kt1 = -0.22076004
+ kt2 = -0.053318302
+ lk2 = -1.2413537e-8
+ llc = 0
+ cdsc = 0
+ lln = 1
+ lu0 = -1.5529956e-9
+ ckappad = 0.6
+ ckappas = 0.6
+ mjd = 0.26
+ mjs = 0.26
+ lua = -8.9830708e-17
+ lub = -5.4824e-26
+ luc = -1.8883822e-17
+ lud = 0
+ lwc = 0
+ cgbo = 0
+ wtvoff = 0
+ lwl = 0
+ lwn = 1
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ pdiblc1 = 0
+ pdiblc2 = 0.014549485
+ njd = 1.02
+ xtis = 3
+ njs = 1.02
+ pa0 = 0
+ pdiblcb = -0.3
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 1.44e-11
+ pbs = 0.52
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ pu0 = -1.2e-18
+ tvoff = 0.0024864064
+ prt = 0
+ pud = 0
+ tvfbsdoff = 0.022
+ rsh = 17.5
+ tcj = 0.00076
+ ijthsfwd = 0.01
+ xjbvd = 1
+ ua1 = 9.685506e-10
+ ub1 = -5.4873129e-19
+ xjbvs = 1
+ uc1 = 6.7696222e-11
+ lk2we = -1.5e-12
+ tpb = 0.0014
+ capmod = 2
+ wa0 = 0
+ ute = -1
+ wat = 0
+ web = 6843.8
+ wec = -25529.0
+ wlc = 0
+ wln = 1
+ wku0we = 2e-11
+ wu0 = 3.6000000000000005e-11
+ xgl = -1.09e-8
+ xgw = 0
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ bigbacc = 0.002588
+ mobmod = 0
+ )

.model nch_sf_4 nmos (
+ level = 54
+ minv = -0.3
+ lua1 = -3.0475764e-17
+ pk2we = -1e-19
+ lub1 = -2.7571927e-26
+ luc1 = -4.3987511e-18
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ ndep = 1e+18
+ rgatemod = 0
+ lwlc = 0
+ moin = 5.1
+ tnjtsswg = 1
+ tnoia = 0
+ nigc = 3.083
+ peta0 = 0.0
+ poxedge = 1
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ tpbsw = 0.0019
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ binunit = 2
+ cjswd = 8.6592e-11
+ cjsws = 8.6592e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ ntox = 1.0
+ pcit = 1.2000000000000001e-17
+ pclm = 1.5439223
+ phin = 0.15
+ pkt1 = -1.76e-16
+ toxref = 3e-9
+ scref = 1e-6
+ jtsswgd = 2.3e-7
+ pigcd = 2.621
+ jtsswgs = 2.3e-7
+ aigsd = 0.01077322
+ rbdb = 50
+ prwb = 0
+ pub1 = 1.6e-34
+ prwg = 0
+ lvoff = -6.3056134e-9
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ rdsw = 100
+ lvsat = 0.00016
+ lvth0 = -4.290877999999999e-9
+ delta = 0.007595625
+ ltvoff = -1.206053e-10
+ laigc = -1.9935708e-11
+ rnoia = 0
+ rnoib = 0
+ ijthsfwd = 0.01
+ ngate = 8e+20
+ njtsswg = 9
+ ngcon = 1
+ rshg = 15.6
+ lku0we = 2.5e-11
+ ags = 0.134315598
+ epsrox = 3.9
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ cjd = 0.001432992
+ cit = 0.00073144105
+ ijthsrev = 0.01
+ cjs = 0.001432992
+ clc = 1e-7
+ cle = 0.6
+ gbmin = 1e-12
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 1.30529375e-8
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ k3b = 1.9326
+ ckappad = 0.6
+ ckappas = 0.6
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ rdsmod = 0
+ pdiblc1 = 0
+ pdiblc2 = 0.027331777
+ pdiblcb = -0.3
+ igbmod = 1
+ la0 = -2.4730306e-7
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.016785258
+ kt1 = -0.23920434
+ kt2 = -0.070668297
+ lk2 = -9.6174482e-9
+ llc = -1.18e-13
+ lln = 0.7
+ lu0 = -6.2833887e-10
+ mjd = 0.26
+ mjs = 0.26
+ lua = -1.0757894e-17
+ lub = -4.7838952e-26
+ luc = -6.6488035e-18
+ lud = 0
+ pbswgd = 0.95
+ pbswgs = 0.95
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ tnom = 25
+ njd = 1.02
+ njs = 1.02
+ pa0 = 0
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 1.44e-11
+ pbs = 0.52
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ pu0 = -1.2e-18
+ igcmod = 1
+ prt = 0
+ pud = 0
+ bigbacc = 0.002588
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 8.041349e-10
+ ub1 = -4.3844738e-19
+ uc1 = 8.6257162e-11
+ tpb = 0.0014
+ wa0 = 0
+ ute = -1
+ wat = 0
+ web = 6843.8
+ wec = -25529.0
+ kvth0we = 0.00018
+ wlc = 0
+ wln = 1
+ wu0 = 3.6000000000000005e-11
+ xgl = -1.09e-8
+ xgw = 0
+ tvoff = 0.0012970146
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ tvfbsdoff = 0.022
+ lintnoi = -1.5e-8
+ xjbvd = 1
+ xjbvs = 1
+ wags = 8e-9
+ lk2we = -1.5e-12
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ wcit = -4.0000000000000004e-11
+ voff = -0.12901018
+ acde = 0.4
+ pkvth0we = -1.3e-19
+ ku0we = -0.0007
+ beta0 = 13
+ vsat = 102860
+ wint = 0
+ permod = 1
+ leta0 = -1.6000000000000003e-9
+ vth0 = 0.44776443
+ wkt1 = 2.5600000000000003e-9
+ wmax = 0.00090001
+ aigc = 0.011598359
+ wmin = 9.0026e-6
+ vfbsdoff = 0.02
+ a0 = 1.6720524
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 150970.13
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.020255575
+ k3 = -1.8419
+ em = 1000000.0
+ dlcig = 2.5e-9
+ ll = -1.18e-13
+ wvfbsdoff = 0
+ lw = 0
+ u0 = 0.013608952
+ bgidl = 2320000000.0
+ w0 = 0
+ lvfbsdoff = 0
+ ua = -2.1226533e-9
+ ub = 2.1407249e-18
+ uc = 6.5910917e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 3.4e-9
+ voffcv = -0.16942
+ wpemod = 1
+ bigc = 0.001442
+ paramchk = 1
+ wwlc = 0
+ wtvfbsdoff = 0
+ dmcgt = 0
+ tcjsw = 0.000357
+ nfactor = 1
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ ltvfbsdoff = 0
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ ijthdfwd = 0.01
+ bigsd = 0.00125
+ tpbswg = 0.0009
+ wvoff = -3.2000000000000003e-10
+ nigbacc = 10
+ wvsat = 0
+ wvth0 = 2.4e-9
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ ijthdrev = 0.01
+ ptvfbsdoff = 0
+ lpdiblc2 = -2.58618e-9
+ ptvoff = 0
+ nigbinv = 10
+ k2we = 5e-5
+ dsub = 0.75
+ lketa = -2.2644187e-8
+ dtox = 2.7e-10
+ xpart = 1
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ diomod = 1
+ pditsd = 0
+ pditsl = 0
+ egidl = 0.29734
+ cjswgd = 2.9779200000000003e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.9779200000000003e-10
+ eta0 = 0.3
+ etab = -0.25
+ fnoimod = 1
+ eigbinv = 1.1
+ lkvth0we = -2e-12
+ mjswgd = 0.85
+ mjswgs = 0.85
+ tcjswg = 0.001
+ acnqsmod = 0
+ rbodymod = 0
+ pvoff = -4e-17
+ cigbacc = 0.32875
+ cdscb = 0
+ cdscd = 0
+ pvsat = 1.44e-11
+ wk2we = 5e-12
+ pvth0 = 1.2e-16
+ drout = 0.56
+ tnoimod = 0
+ fprout = 300
+ voffl = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ cigbinv = 0.006
+ weta0 = 0
+ lpclm = -6.3325799e-8
+ wtvoff = 0
+ version = 4.5
+ cgidl = 0.22
+ tempmod = 0
+ keta = -0.039946614
+ capmod = 2
+ lags = 5.5033282e-7
+ wku0we = 2e-11
+ aigbacc = 0.02
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 1.7016594e-10
+ pbswd = 0.8
+ mobmod = 0
+ pbsws = 0.8
+ kt1l = 0
+ wkvth0we = 2e-12
+ pvfbsdoff = 0
+ lint = 9.7879675e-9
+ trnqsmod = 0
+ pdits = 0
+ lkt1 = -9.8888734e-9
+ lkt2 = -3.8595493e-9
+ aigbinv = 0.0163
+ lmax = 4.4908e-7
+ cigsd = 0.069865
+ lmin = 2.1577e-7
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ laigsd = -8.1082969e-17
+ )

.model nch_sf_5 nmos (
+ level = 54
+ nigbinv = 10
+ bigsd = 0.00125
+ wags = 8e-9
+ wcit = -4.0000000000000004e-11
+ acnqsmod = 0
+ wvoff = -3.2000000000000003e-10
+ voff = -0.15746310460000001
+ acde = 0.4
+ wvsat = 0
+ vsat = 102521.2852
+ wvth0 = 2.4e-9
+ rbodymod = 0
+ wint = 0
+ vth0 = 0.4637613742
+ wkt1 = 2.5600000000000003e-9
+ wmax = 0.00090001
+ aigc = 0.011526753
+ wmin = 9.0026e-6
+ fnoimod = 1
+ eigbinv = 1.1
+ toxref = 3e-9
+ lketa = -1.1430034e-8
+ xpart = 1
+ bigc = 0.001442
+ wwlc = 0
+ egidl = 0.29734
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ ltvoff = 1.4850105e-11
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ cigbacc = 0.32875
+ tnoimod = 0
+ lku0we = 2.5e-11
+ cigbinv = 0.006
+ epsrox = 3.9
+ wkvth0we = 2e-12
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ pvoff = -4e-17
+ rdsmod = 0
+ trnqsmod = 0
+ cdscb = 0
+ cdscd = 0
+ igbmod = 1
+ pvsat = 1.44e-11
+ version = 4.5
+ wk2we = 5e-12
+ pvth0 = 1.2e-16
+ k2we = 5e-5
+ drout = 0.56
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ tempmod = 0
+ dsub = 0.75
+ dtox = 2.7e-10
+ pbswgd = 0.95
+ pbswgs = 0.95
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ voffl = 0
+ igcmod = 1
+ aigbacc = 0.02
+ weta0 = 0
+ eta0 = 0.3
+ rgatemod = 0
+ etab = -0.25
+ lpclm = -2.4377173e-8
+ tnjtsswg = 1
+ cgidl = 0.22
+ aigbinv = 0.0163
+ pbswd = 0.8
+ pbsws = 0.8
+ pvfbsdoff = 0
+ permod = 1
+ wtvfbsdoff = 0
+ pdits = 0
+ cigsd = 0.069865
+ dvt0w = 0
+ dvt1w = 0
+ poxedge = 1
+ dvt2w = 0
+ ltvfbsdoff = 0
+ voffcv = -0.16942
+ wpemod = 1
+ binunit = 2
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ tnoia = 0
+ peta0 = 0.0
+ wketa = 0
+ keta = -0.093093889
+ ptvfbsdoff = 0
+ tpbsw = 0.0019
+ ijthsfwd = 0.01
+ cjswd = 8.6592e-11
+ cjsws = 8.6592e-11
+ a0 = 0.66068814
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ mjswd = 0.11
+ lags = 3.3904274e-13
+ mjsws = 0.11
+ agidl = 9.41e-8
+ tpbswg = 0.0009
+ at = 79499.116
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = -0.014512077999999998
+ k3 = -1.8419
+ em = 1000000.0
+ jswd = 1.28e-13
+ ll = -1.18e-13
+ jsws = 1.28e-13
+ lw = 0
+ u0 = 0.011606872
+ w0 = 0
+ lcit = 9.2591162e-11
+ ua = -2.2893587e-9
+ ub = 2.089788886e-18
+ uc = 4.5969231e-11
+ ud = 0
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 3.4e-9
+ kt1l = 0
+ ijthsrev = 0.01
+ lint = 9.7879675e-9
+ ptvoff = 0
+ lkt1 = -3.5475226e-9
+ lkt2 = -6.0180086e-10
+ lmax = 2.1577e-7
+ lmin = 9e-8
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ scref = 1e-6
+ diomod = 1
+ pigcd = 2.621
+ minv = -0.3
+ aigsd = 0.01077322
+ lua1 = 7.6861327e-18
+ lub1 = -4.9942255999999997e-26
+ luc1 = -4.2210821e-18
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 2.9779200000000003e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.9779200000000003e-10
+ ndep = 1e+18
+ lvoff = -3.020626000000001e-10
+ njtsswg = 9
+ lwlc = 0
+ moin = 5.1
+ lvsat = 0.0002314843
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ lvth0 = -7.6662159e-9
+ nigc = 3.083
+ delta = 0.007595625
+ mjswgd = 0.85
+ mjswgs = 0.85
+ laigc = -4.8268328e-12
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.02163037
+ pdiblcb = -0.3
+ tcjswg = 0.001
+ rnoia = 0
+ rnoib = 0
+ ags = 2.7425264
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ cjd = 0.001432992
+ cit = 0.001099094
+ cjs = 0.001432992
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 1.30529375e-8
+ pketa = 0
+ ngate = 8e+20
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ ngcon = 1
+ pkvth0we = -1.3e-19
+ ntox = 1.0
+ pcit = 1.2000000000000001e-17
+ pclm = 1.3593316
+ bigbacc = 0.002588
+ la0 = -3.3904685e-8
+ gbmin = 1e-12
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.0017048735
+ kt1 = -0.26925814
+ kt2 = -0.086107863
+ lk2 = -2.2814734e-9
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ llc = -1.18e-13
+ lln = 0.7
+ phin = 0.15
+ lu0 = -2.0589995000000002e-10
+ mjd = 0.26
+ mjs = 0.26
+ lua = 2.4416942e-17
+ lub = -3.7091512499999996e-26
+ luc = -2.4411077e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ vfbsdoff = 0.02
+ njd = 1.02
+ njs = 1.02
+ pa0 = 0
+ nsd = 1e+20
+ kvth0we = 0.00018
+ pbd = 0.52
+ pat = 1.44e-11
+ pbs = 0.52
+ pkt1 = -1.76e-16
+ pu0 = -1.2e-18
+ prt = 0
+ fprout = 300
+ pub = 0
+ pud = 0
+ lintnoi = -1.5e-8
+ rsh = 17.5
+ xrcrg1 = 12
+ xrcrg2 = 1
+ tcj = 0.00076
+ ua1 = 6.2327283e-10
+ ub1 = -3.3242687e-19
+ uc1 = 8.5415128e-11
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ tpb = 0.0014
+ wa0 = 0
+ ute = -1
+ paramchk = 1
+ wat = 0
+ web = 6843.8
+ wec = -25529.0
+ wlc = 0
+ wln = 1
+ wu0 = 3.6000000000000005e-11
+ rbdb = 50
+ xgl = -1.09e-8
+ prwb = 0
+ pub1 = 1.6e-34
+ prwg = 0
+ xgw = 0
+ wub = 0
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ rbpb = 50
+ rbpd = 50
+ wtvoff = 0
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ rdsw = 100
+ tvfbsdoff = 0.022
+ tvoff = 0.00065504585
+ capmod = 2
+ ijthdfwd = 0.01
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ wku0we = 2e-11
+ mobmod = 0
+ rshg = 15.6
+ ku0we = -0.0007
+ beta0 = 13
+ leta0 = -1.6000000000000003e-9
+ ijthdrev = 0.01
+ nfactor = 1
+ lpdiblc2 = -1.3831831e-9
+ wvfbsdoff = 0
+ dlcig = 2.5e-9
+ lvfbsdoff = 0
+ bgidl = 2320000000.0
+ laigsd = 3.3904273e-17
+ tnom = 25
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ nigbacc = 10
+ dmcgt = 0
+ tcjsw = 0.000357
+ lkvth0we = -2e-12
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ )

.model nch_sf_6 nmos (
+ level = 54
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ vfbsdoff = 0.02
+ toxref = 3e-9
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.0069155858
+ scref = 1e-6
+ pdiblcb = -0.3
+ pigcd = 2.621
+ aigsd = 0.01077322
+ paramchk = 1
+ lvoff = -2.04841089e-9
+ ags = 2.74253
+ lvsat = 0.0017264268699999999
+ ltvoff = 1.0839662e-10
+ lvth0 = 2.64929317e-9
+ bigbacc = 0.002588
+ cjd = 0.001432992
+ cit = 0.00031861111
+ cjs = 0.001432992
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ delta = 0.007595625
+ dlc = 3.26497e-9
+ k3b = 1.9326
+ laigc = -2.2427226e-11
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ keta = -0.52835722
+ rnoia = 0
+ rnoib = 0
+ ijthdfwd = 0.01
+ kvth0we = 0.00018
+ la0 = 3.0288889e-8
+ jsd = 6.11e-7
+ lintnoi = -1.5e-8
+ jss = 6.11e-7
+ lat = -0.00030029214
+ kt1 = -0.40872879
+ kt2 = -0.10088778
+ lk2 = -4.8654938e-10
+ lku0we = 2.5e-11
+ pketa = 0
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ ngate = 8e+20
+ bigbinv = 0.004953
+ llc = 0
+ lln = 1
+ lu0 = 9.883078000000001e-11
+ lcit = 1.6595656e-10
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ mjd = 0.26
+ mjs = 0.26
+ lua = 3.5218789e-17
+ lub = -1.9869262700000004e-26
+ luc = 2.2716666e-18
+ lud = 0
+ epsrox = 3.9
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ ngcon = 1
+ njd = 1.02
+ njs = 1.02
+ kt1l = 0
+ pa0 = 0
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 1.44e-11
+ pbs = 0.52
+ pu0 = -1.2e-18
+ prt = 0
+ pub = 0
+ puc = 0
+ pud = 0
+ rdsmod = 0
+ ijthdrev = 0.01
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ rsh = 17.5
+ jswgs = 1.28e-13
+ lint = 0
+ tcj = 0.00076
+ igbmod = 1
+ ua1 = 8.897383e-10
+ ub1 = -8.0235504e-19
+ uc1 = -6.3390556e-11
+ tpb = 0.0014
+ lkt1 = 9.5627184e-9
+ lkt2 = 7.8751111e-10
+ wa0 = 0
+ lpdiblc2 = 6.6256944e-15
+ lmax = 9e-8
+ ute = -1
+ wat = 0
+ web = 6843.8
+ pscbe1 = 1000000000.0
+ wec = -25529.0
+ pscbe2 = 1e-20
+ lmin = 5.4e-8
+ wlc = 0
+ wln = 1
+ wu0 = 3.6000000000000005e-11
+ xgl = -1.09e-8
+ xgw = 0
+ wub = 0
+ wuc = 0
+ wud = 0
+ lpe0 = 9.2e-8
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ pbswgd = 0.95
+ lpeb = 2.5e-7
+ pbswgs = 0.95
+ minv = -0.3
+ igcmod = 1
+ lua1 = -1.7361621e-17
+ lub1 = -5.7690078e-27
+ luc1 = 9.7666522e-18
+ ndep = 1e+18
+ lwlc = 0
+ moin = 5.1
+ nigc = 3.083
+ tvfbsdoff = 0.022
+ nfactor = 1
+ lkvth0we = -2e-12
+ tvoff = -0.00034012981
+ wtvfbsdoff = 0
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ acnqsmod = 0
+ ltvfbsdoff = 0
+ permod = 1
+ ntox = 1.0
+ pcit = 1.2000000000000001e-17
+ ku0we = -0.0007
+ pclm = 1.2209944
+ beta0 = 13
+ rbodymod = 0
+ leta0 = 1.4288888999999997e-9
+ nigbacc = 10
+ letab = -2.2684433e-8
+ phin = 0.15
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ pkt1 = -1.76e-16
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ voffcv = -0.16942
+ wpemod = 1
+ nigbinv = 10
+ ptvfbsdoff = 0
+ rbdb = 50
+ prwb = 0
+ pub1 = 1.6e-34
+ prwg = 0
+ dmcgt = 0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ tcjsw = 0.000357
+ rdsw = 100
+ fnoimod = 1
+ eigbinv = 1.1
+ bigsd = 0.00125
+ tpbswg = 0.0009
+ wvoff = -3.2000000000000003e-10
+ rshg = 15.6
+ wkvth0we = 2e-12
+ wvsat = 0.0
+ wvth0 = 2.4e-9
+ ptvoff = 0
+ trnqsmod = 0
+ cigbacc = 0.32875
+ diomod = 1
+ lketa = 2.9484719e-8
+ xpart = 1
+ pditsd = 0
+ pditsl = 0
+ tnoimod = 0
+ cjswgd = 2.9779200000000003e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.9779200000000003e-10
+ tnom = 25
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ egidl = 0.29734
+ a0 = -0.02222221999999996
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ rgatemod = 0
+ at = 64556.761
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = -0.033607015000000004
+ k3 = -1.8419
+ em = 1000000.0
+ cigbinv = 0.006
+ ll = 0
+ lw = 0
+ u0 = 0.0083650556
+ tnjtsswg = 1
+ w0 = 0
+ ua = -2.404272e-9
+ ub = 1.906573466e-18
+ uc = -4.166667e-12
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 3.4e-9
+ mjswgd = 0.85
+ mjswgs = 0.85
+ tcjswg = 0.001
+ version = 4.5
+ wags = 8e-9
+ tempmod = 0
+ wcit = -4.0000000000000004e-11
+ voff = -0.138884931
+ acde = 0.4
+ aigbacc = 0.02
+ vsat = 86617.64
+ wint = 0
+ vth0 = 0.354021916
+ pvoff = -4e-17
+ wkt1 = 2.5600000000000003e-9
+ wmax = 0.00090001
+ aigc = 0.011713991
+ wmin = 9.0026e-6
+ cdscb = 0
+ cdscd = 0
+ pvsat = 1.44e-11
+ wk2we = 5e-12
+ pvth0 = 1.2e-16
+ fprout = 300
+ drout = 0.56
+ xrcrg1 = 12
+ xrcrg2 = 1
+ aigbinv = 0.0163
+ voffl = 0
+ bigc = 0.001442
+ wwlc = 0
+ wtvoff = 0
+ weta0 = 0
+ lpclm = -1.1373478e-8
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ cgidl = 0.22
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ capmod = 2
+ wku0we = 2e-11
+ ijthsfwd = 0.01
+ poxedge = 1
+ mobmod = 0
+ pbswd = 0.8
+ pvfbsdoff = 0
+ pbsws = 0.8
+ binunit = 2
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ ijthsrev = 0.01
+ pdits = 0
+ cigsd = 0.069865
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ k2we = 5e-5
+ dsub = 0.75
+ dtox = 2.7e-10
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ eta0 = 0.26777778
+ etab = -0.0086762422
+ tnoia = 0
+ peta0 = 0.0
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ wketa = 0
+ tpbsw = 0.0019
+ cjswd = 8.6592e-11
+ cjsws = 8.6592e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ pkvth0we = -1.3e-19
+ njtsswg = 9
+ )

.model nch_sf_7 nmos (
+ level = 54
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ ltvoff = -2.4740506e-10
+ aigbacc = 0.02
+ rdsw = 100
+ ijthsfwd = 0.01
+ lku0we = 2.5e-11
+ aigbinv = 0.0163
+ epsrox = 3.9
+ rshg = 15.6
+ rdsmod = 0
+ igbmod = 1
+ ijthsrev = 0.01
+ pvoff = -4e-17
+ cdscb = 0
+ cdscd = 0
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ pvsat = 1.44e-11
+ wk2we = 5e-12
+ pvth0 = 1.2e-16
+ drout = 0.56
+ pbswgd = 0.95
+ pbswgs = 0.95
+ igcmod = 1
+ poxedge = 1
+ wtvfbsdoff = 0
+ voffl = 0
+ tnom = 25
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ weta0 = 0
+ binunit = 2
+ lpclm = -7.2871722e-8
+ ltvfbsdoff = 0
+ cgidl = 0.22
+ wags = 8e-9
+ wcit = -4.0000000000000004e-11
+ pvfbsdoff = 0
+ permod = 1
+ pbswd = 0.8
+ pbsws = 0.8
+ voff = -0.112415764
+ pkvth0we = -1.3e-19
+ acde = 0.4
+ ptvfbsdoff = 0
+ vsat = 86759.482
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ wint = 0
+ vth0 = 0.351917597
+ wkt1 = 2.5600000000000003e-9
+ wmax = 0.00090001
+ aigc = 0.011692671
+ pdits = 0
+ wmin = 9.0026e-6
+ vfbsdoff = 0.02
+ cigsd = 0.069865
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ voffcv = -0.16942
+ wpemod = 1
+ wub1 = 0.0
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ bigc = 0.001442
+ paramchk = 1
+ wwlc = 0
+ tnoia = 0
+ cdsc = 0
+ cgbo = 0
+ njtsswg = 9
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ peta0 = 0.0
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ tpbsw = 0.0019
+ ijthdfwd = 0.01
+ tpbswg = 0.0009
+ ckappad = 0.6
+ cjswd = 8.6592e-11
+ ckappas = 0.6
+ cjsws = 8.6592e-11
+ mjswd = 0.11
+ pdiblc1 = 0
+ pdiblc2 = 0.0069157
+ mjsws = 0.11
+ agidl = 9.41e-8
+ pdiblcb = -0.3
+ ptvoff = 0
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ ijthdrev = 0.01
+ bigbacc = 0.002588
+ diomod = 1
+ k2we = 5e-5
+ dsub = 0.75
+ scref = 1e-6
+ dtox = 2.7e-10
+ pditsd = 0
+ pditsl = 0
+ kvth0we = 0.00018
+ cjswgd = 2.9779200000000003e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.9779200000000003e-10
+ ags = 2.74253
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ pigcd = 2.621
+ aigsd = 0.01077322
+ cjd = 0.001432992
+ cit = -0.0027423847
+ cjs = 0.001432992
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ lintnoi = -1.5e-8
+ dlc = 3.26497e-9
+ bigbinv = 0.004953
+ k3b = 1.9326
+ lvoff = -3.5836221999999995e-9
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ eta0 = 0.35179556
+ etab = -1.0973583
+ lvsat = 0.0017182000999999996
+ mjswgd = 0.85
+ mjswgs = 0.85
+ lvth0 = 2.7713433000000007e-9
+ la0 = -3.1577778e-7
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = 0.0076586667
+ lkvth0we = -2e-12
+ kt1 = 0.010917511
+ kt2 = -0.10990444
+ lk2 = -1.5787889e-9
+ delta = 0.007595625
+ tcjswg = 0.001
+ llc = 0
+ laigc = -2.1190647e-11
+ lln = 1
+ lu0 = 5.429271100000001e-10
+ mjd = 0.26
+ mjs = 0.26
+ lua = 7.8730998e-17
+ lub = -4.3148946000000005e-26
+ luc = 1.578889e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 0
+ rnoia = 0
+ rnoib = 0
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 1.44e-11
+ pbs = 0.52
+ pu0 = -1.2e-18
+ prt = 0
+ pub = 0
+ puc = 0
+ pud = 0
+ acnqsmod = 0
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 3.744227e-10
+ ngate = 8e+20
+ ub1 = -1.4506222e-18
+ uc1 = -1.6722222e-10
+ tpb = 0.0014
+ ngcon = 1
+ wa0 = 0
+ ute = -1
+ wat = 0.0
+ web = 6843.8
+ wec = -25529.0
+ wlc = 0
+ wln = 1
+ wu0 = 3.6000000000000005e-11
+ xgl = -1.09e-8
+ xgw = 0
+ wub = 0
+ wuc = 0
+ wud = 0
+ rbodymod = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ a0 = 5.9444444
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = -72666.667
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = -0.014775298999999999
+ k3 = -1.8419
+ em = 1000000.0
+ fprout = 300
+ ll = 0
+ lw = 0
+ u0 = 0.0007082222200000001
+ nfactor = 1
+ w0 = 0
+ ua = -3.1544825e-9
+ ub = 2.30794738e-18
+ uc = 7.77778e-12
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 3.4e-9
+ xrcrg1 = 12
+ xrcrg2 = 1
+ wtvoff = 0
+ tvfbsdoff = 0.022
+ nigbacc = 10
+ capmod = 2
+ tvoff = 0.0057943818
+ wku0we = 2e-11
+ keta = 0.088888889
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ mobmod = 0
+ nigbinv = 10
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 3.4349431000000004e-10
+ kt1l = 0
+ ku0we = -0.0007
+ wkvth0we = 2e-12
+ beta0 = 13
+ leta0 = -3.4441422000000003e-9
+ letab = 4.0459126e-8
+ lint = 0
+ trnqsmod = 0
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ lkt1 = -1.4776766999999999e-8
+ lkt2 = 1.3104778e-9
+ lmax = 5.4e-8
+ lmin = 4.5e-8
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ lpe0 = 9.2e-8
+ fnoimod = 1
+ lpeb = 2.5e-7
+ eigbinv = 1.1
+ minv = -0.3
+ lua1 = 1.2526683e-17
+ lub1 = 3.1830488999999997e-26
+ luc1 = 1.5788889e-17
+ ndep = 1e+18
+ dmcgt = 0
+ rgatemod = 0
+ lwlc = 0
+ tcjsw = 0.000357
+ moin = 5.1
+ tnjtsswg = 1
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ nigc = 3.083
+ bigsd = 0.00125
+ noff = 2.7195
+ cigbacc = 0.32875
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ wvoff = -3.2000000000000003e-10
+ tnoimod = 0
+ ntox = 1.0
+ pcit = 1.2000000000000001e-17
+ pclm = 2.281309
+ wvsat = 0.0
+ wvth0 = 2.4e-9
+ cigbinv = 0.006
+ phin = 0.15
+ toxref = 3e-9
+ pkt1 = -1.76e-16
+ lketa = -6.3155556e-9
+ version = 4.5
+ xpart = 1
+ tempmod = 0
+ egidl = 0.29734
+ rbdb = 50
+ prwb = 0
+ pub1 = 1.6e-34
+ prwg = 0
+ )

.model nch_sf_8 nmos (
+ level = 54
+ ngate = 8e+20
+ ngcon = 1
+ wpclm = 0
+ rdsmod = 0
+ wkvth0we = 2e-12
+ wtvfbsdoff = 0
+ igbmod = 1
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ trnqsmod = 0
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ nigbacc = 10
+ ltvfbsdoff = 0
+ pbswgd = 0.95
+ pbswgs = 0.95
+ k2we = 5e-5
+ igcmod = 1
+ dsub = 0.75
+ dtox = 2.7e-10
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ nigbinv = 10
+ rgatemod = 0
+ eta0 = -0.001232
+ etab = -0.88502038
+ tnjtsswg = 1
+ tvfbsdoff = 0.022
+ ptvfbsdoff = 0
+ tvoff = 0.0030235155
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ fnoimod = 1
+ permod = 1
+ eigbinv = 1.1
+ ku0we = -0.0007
+ beta0 = 13
+ leta0 = 1.3854208e-8
+ letab = 3.0054568e-8
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ ppclm = 0
+ voffcv = -0.16942
+ wpemod = 1
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ cigbacc = 0.32875
+ dmcgt = 0
+ tnoimod = 0
+ tcjsw = 0.000357
+ cigbinv = 0.006
+ tpbswg = 0.0009
+ keta = 0.44888889
+ ijthsfwd = 0.01
+ bigsd = 0.00125
+ version = 4.5
+ wvoff = -3.2000000000000003e-10
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 3.7725569000000003e-10
+ tempmod = 0
+ kt1l = 0
+ ptvoff = 0
+ wvsat = 0.0
+ wvth0 = 2.4e-9
+ ijthsrev = 0.01
+ lint = 0
+ aigbacc = 0.02
+ lkt1 = -4.1488498e-9
+ lkt2 = 1.6072e-9
+ diomod = 1
+ lmax = 4.5e-8
+ lmin = 3.6e-8
+ lpe0 = 9.2e-8
+ pditsd = 0
+ pditsl = 0
+ lketa = -2.3955556e-8
+ lpeb = 2.5e-7
+ cjswgd = 2.9779200000000003e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.9779200000000003e-10
+ xpart = 1
+ minv = -0.3
+ aigbinv = 0.0163
+ lua1 = 7.1708778e-18
+ lub1 = -2.1542999e-26
+ luc1 = -1.63268e-17
+ egidl = 0.29734
+ ndep = 1e+18
+ lwlc = 0
+ mjswgd = 0.85
+ mjswgs = 0.85
+ moin = 5.1
+ nigc = 3.083
+ tcjswg = 0.001
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ poxedge = 1
+ pkvth0we = -1.3e-19
+ ntox = 1.0
+ pcit = 1.2000000000000001e-17
+ pclm = 2.10165423
+ binunit = 2
+ pvoff = -4e-17
+ fprout = 300
+ phin = 0.15
+ cdscb = 0
+ cdscd = 0
+ vfbsdoff = 0.02
+ pvsat = 1.44e-11
+ xrcrg1 = 12
+ xrcrg2 = 1
+ wk2we = 5e-12
+ pvth0 = 1.2e-16
+ drout = 0.56
+ pkt1 = -1.76e-16
+ voffl = 0
+ wtvoff = 0
+ paramchk = 1
+ weta0 = 0
+ rbdb = 50
+ prwb = 0
+ pub1 = 1.6e-34
+ prwg = 0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ lpclm = -6.406864000000001e-8
+ rdsw = 100
+ capmod = 2
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ cgidl = 0.22
+ wku0we = 2e-11
+ mobmod = 0
+ ijthdfwd = 0.01
+ a0 = 3.6555556
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 123237.73
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.025756861000000002
+ k3 = -1.8419
+ em = 1000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.005247777299999999
+ pvfbsdoff = 0
+ w0 = 0
+ ua = -2.2580401200000003e-9
+ ub = 1.5627388499999998e-18
+ uc = 2.4e-10
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 3.4e-9
+ pbswd = 0.8
+ pbsws = 0.8
+ rshg = 15.6
+ ijthdrev = 0.01
+ pdits = 0
+ njtsswg = 9
+ cigsd = 0.069865
+ laigsd = -2.1777778e-17
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ ckappad = 0.6
+ ckappas = 0.6
+ pk2we = -1e-19
+ tnom = 25
+ pdiblc1 = 0
+ pdiblc2 = 0.0069157
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ pdiblcb = -0.3
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ tnoia = 0
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ peta0 = 0.0
+ lkvth0we = -2e-12
+ bigbacc = 0.002588
+ tpbsw = 0.0019
+ wags = 8e-9
+ cjswd = 8.6592e-11
+ cjsws = 8.6592e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ wcit = -4.0000000000000004e-11
+ kvth0we = 0.00018
+ acnqsmod = 0
+ voff = -0.039834349000000005
+ acde = 0.4
+ lintnoi = -1.5e-8
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ vsat = 76593.03200000002
+ rbodymod = 0
+ vtsswgs = 4.2
+ wint = 0
+ vth0 = 0.355739103
+ toxref = 3e-9
+ wkt1 = 2.5600000000000003e-9
+ ags = 2.74253
+ wmax = 0.00090001
+ aigc = 0.011387162
+ wmin = 9.0026e-6
+ cjd = 0.001432992
+ cit = -0.0034313898000000002
+ cjs = 0.001432992
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 3.26497e-9
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ scref = 1e-6
+ wub1 = 0.0
+ pigcd = 2.621
+ aigsd = 0.010773221
+ la0 = -2.0362223e-7
+ bigc = 0.001442
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.0019406488000000002
+ kt1 = -0.20597876
+ kt2 = -0.11596
+ lk2 = -3.5648647e-9
+ wwlc = 0
+ llc = 0
+ lvoff = -7.140111900000001e-9
+ lln = 1
+ lu0 = 3.2048887e-10
+ mjd = 0.26
+ mjs = 0.26
+ lua = 3.4805321000000004e-17
+ lub = -6.633731000000002e-27
+ luc = -9.7999999e-18
+ lud = 0
+ ltvoff = -1.1163261e-10
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 0
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 1.44e-11
+ pbs = 0.52
+ pk2 = 0
+ lvsat = 0.0022163563900000002
+ cdsc = 0
+ pu0 = -1.2e-18
+ lvth0 = 2.5840918800000004e-9
+ prt = 0
+ cgbo = 0
+ pua = 0
+ pub = 0
+ puc = 0
+ pud = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ delta = 0.007595625
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 4.8372486e-10
+ ub1 = -3.6136738e-19
+ cigc = 0.000625
+ laigc = -6.2207351e-12
+ uc1 = 4.882e-10
+ tpb = 0.0014
+ wa0 = 0
+ rnoia = 0
+ rnoib = 0
+ nfactor = 1
+ ute = -1
+ wat = 0.0
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 0
+ wlc = 0
+ lku0we = 2.5e-11
+ wln = 1
+ wu0 = 3.6000000000000005e-11
+ xgl = -1.09e-8
+ xgw = 0
+ wua = 0
+ wub = 0
+ wuc = 0
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ epsrox = 3.9
+ )

.model nch_sf_9 nmos (
+ level = 54
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ ptvfbsdoff = 0
+ voffl = 0
+ minv = -0.3
+ lub1 = 2.4000000000000004e-27
+ weta0 = 0
+ ndep = 1e+18
+ wetab = -1.0073378e-8
+ lwlc = 0
+ moin = 5.1
+ nigc = 3.083
+ cgidl = 0.22
+ lkvth0we = -2e-12
+ njtsswg = 9
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ pvfbsdoff = 0
+ noic = 45200000.0
+ permod = 1
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ acnqsmod = 0
+ pbswd = 0.8
+ pbsws = 0.8
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.018557155
+ pdiblcb = -0.3
+ ntox = 1.0
+ pcit = 1.2000000000000001e-17
+ pclm = 1.4152454
+ rbodymod = 0
+ phin = 0.15
+ voffcv = -0.16942
+ wpemod = 1
+ pdits = 0
+ cigsd = 0.069865
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ pkt1 = -1.76e-16
+ bigbacc = 0.002588
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ kvth0we = 0.00018
+ rbdb = 50
+ prwb = 0
+ pub1 = 1.6e-34
+ prwg = 0
+ wpdiblc2 = -1.7177628e-11
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ lintnoi = -1.5e-8
+ tnoia = 0
+ bigbinv = 0.004953
+ rdsw = 100
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ peta0 = 0.0
+ tpbswg = 0.0009
+ wketa = 3.3422159e-8
+ tpbsw = 0.0019
+ cjswd = 8.6592e-11
+ cjsws = 8.6592e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ ags = 0.9568331400000001
+ ptvoff = 0
+ cjd = 0.001432992
+ cit = 4.8708935e-5
+ cjs = 0.001432992
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ wkvth0we = 2e-12
+ bvs = 8.7
+ rshg = 15.6
+ waigsd = 3.0716751e-12
+ dlc = 9.8024918e-9
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ trnqsmod = 0
+ diomod = 1
+ la0 = 0
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = 8e-5
+ kt1 = -0.19515831
+ kt2 = -0.052853133
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 2.9779200000000003e-10
+ llc = 0
+ pku0we = -1.5e-18
+ lln = 1
+ cjswgs = 2.9779200000000003e-10
+ lu0 = -4e-12
+ mjd = 0.26
+ mjs = 0.26
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ scref = 1e-6
+ njd = 1.02
+ njs = 1.02
+ pa0 = 0
+ nfactor = 1
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 1.44e-11
+ pbs = 0.52
+ pigcd = 2.621
+ aigsd = 0.010772879
+ pu0 = -1.2e-18
+ prt = 0
+ pud = 0
+ tnom = 25
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 1.311952e-9
+ toxe = 2.43e-9
+ ub1 = -8.0649865e-19
+ toxm = 2.43e-9
+ lvoff = 1.6e-11
+ uc1 = 3.0375074e-11
+ mjswgd = 0.85
+ mjswgs = 0.85
+ tpb = 0.0014
+ rgatemod = 0
+ wa0 = -2.5183444e-7
+ ute = -0.96248296
+ wat = 0
+ tnjtsswg = 1
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -3.7920026e-9
+ lvsat = 0.00016
+ wlc = 0
+ tcjswg = 0.001
+ wln = 1
+ wu0 = -2.2590781999999998e-10
+ xgl = -1.09e-8
+ xgw = 0
+ lvth0 = 4.0000000000000007e-10
+ wua = -4.0765791e-17
+ wub = 4.0599742e-26
+ wuc = -7.8572347e-18
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ delta = 0.007595625
+ nigbacc = 10
+ rnoia = 0
+ rnoib = 0
+ wags = -7.6054279e-8
+ wcit = 4.2192733e-10
+ ngate = 8e+20
+ voff = -0.11308442
+ ngcon = 1
+ wpclm = -1.3730014e-7
+ acde = 0.4
+ nigbinv = 10
+ vsat = 103058.98
+ wint = 0
+ gbmin = 1e-12
+ vth0 = 0.37754845
+ fprout = 300
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ wkt1 = -4.3079654e-8
+ wkt2 = -3.5741805e-9
+ wmax = 9.0026e-6
+ xrcrg1 = 12
+ xrcrg2 = 1
+ aigc = 0.011766468
+ wmin = 9.025999999999999e-7
+ wtvoff = -8.3463378e-10
+ wua1 = -7.3834184e-16
+ wub1 = 7.3798399e-25
+ wuc1 = -8.5623711e-19
+ fnoimod = 1
+ bigc = 0.001442
+ wute = -4.0092044e-7
+ eigbinv = 1.1
+ wwlc = 0
+ tvfbsdoff = 0.022
+ capmod = 2
+ cdsc = 0
+ cgbo = 0
+ wku0we = 2e-11
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ tvoff = 0.0020036382
+ cigc = 0.000625
+ mobmod = 0
+ xjbvd = 1
+ ijthsfwd = 0.01
+ xjbvs = 1
+ lk2we = -1.5e-12
+ cigbacc = 0.32875
+ ku0we = -0.0007
+ beta0 = 13
+ leta0 = -1.6000000000000003e-9
+ tnoimod = 0
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ ijthsrev = 0.01
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ cigbinv = 0.006
+ dlcig = 2.5e-9
+ k2we = 5e-5
+ bgidl = 2320000000.0
+ dsub = 0.75
+ dtox = 2.7e-10
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ a0 = 3.277963
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ version = 4.5
+ at = 72000
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.026622307
+ k3 = -1.8419
+ em = 1000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.016019082
+ dmcgt = 0
+ w0 = 0
+ tempmod = 0
+ ua = -1.8192461e-9
+ ub = 2.0991879e-18
+ uc = 7.4172444e-11
+ ud = 0
+ eta0 = 0.3
+ tcjsw = 0.000357
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ alpha0 = 2e-10
+ ww = 0
+ alpha1 = 3.6
+ xw = 3.4e-9
+ etab = -0.24888148
+ aigbacc = 0.02
+ bigsd = 0.00125
+ wvoff = 2.0577201e-9
+ pkvth0we = -1.3e-19
+ aigbinv = 0.0163
+ wvsat = -0.0017920539
+ wvth0 = -8.745485e-9
+ toxref = 3e-9
+ waigc = 2.6350949e-11
+ vfbsdoff = 0.02
+ xpart = 1
+ paramchk = 1
+ ltvoff = 0
+ egidl = 0.29734
+ poxedge = 1
+ binunit = 2
+ wtvfbsdoff = 0
+ keta = -0.063711099
+ lku0we = 2.5e-11
+ ijthdfwd = 0.01
+ epsrox = 3.9
+ ltvfbsdoff = 0
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 8e-12
+ rdsmod = 0
+ kt1l = 0
+ igbmod = 1
+ ijthdrev = 0.01
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ pvoff = -4e-17
+ lint = 6.5375218e-9
+ pbswgd = 0.95
+ cdscb = 0
+ cdscd = 0
+ pbswgs = 0.95
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ lkt1 = -2.4e-10
+ pvsat = 1.44e-11
+ lmax = 2.001e-5
+ wk2we = 5e-12
+ pvth0 = 1.2e-16
+ lmin = 8.9991e-6
+ drout = 0.56
+ igcmod = 1
+ )

.model nch_sf_10 nmos (
+ level = 54
+ xrcrg1 = 12
+ xrcrg2 = 1
+ cgidl = 0.22
+ vfbsdoff = 0.02
+ wtvoff = -8.9580408e-10
+ nfactor = 1
+ pbswd = 0.8
+ pbsws = 0.8
+ paramchk = 1
+ capmod = 2
+ wku0we = 2e-11
+ mobmod = 0
+ pdits = 0
+ cigsd = 0.069865
+ nigbacc = 10
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ ijthdfwd = 0.01
+ keta = -0.064075044
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ nigbinv = 10
+ lags = -6.3328546e-8
+ wtvfbsdoff = 0
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 1.1417416e-9
+ tnoia = 0
+ laigsd = 1.1048614e-17
+ ijthdrev = 0.01
+ kt1l = 0
+ peta0 = 0.0
+ ltvfbsdoff = 0
+ lpdiblc2 = -6.1589259e-10
+ wketa = 3.7630763e-8
+ lint = 6.5375218e-9
+ tpbsw = 0.0019
+ lkt1 = -4.5777316e-8
+ lkt2 = -1.2972142e-8
+ cjswd = 8.6592e-11
+ lmax = 8.9991e-6
+ cjsws = 8.6592e-11
+ lmin = 8.9908e-7
+ fnoimod = 1
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ lpe0 = 9.2e-8
+ eigbinv = 1.1
+ lpeb = 2.5e-7
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ minv = -0.3
+ lua1 = -4.3996966e-16
+ lub1 = 2.6300002e-25
+ luc1 = 3.9191378e-17
+ ndep = 1e+18
+ lute = -3.7058959e-8
+ lwlc = 0
+ ptvfbsdoff = 0
+ moin = 5.1
+ lkvth0we = -2e-12
+ nigc = 3.083
+ scref = 1e-6
+ pigcd = 2.621
+ aigsd = 0.010772879
+ cigbacc = 0.32875
+ acnqsmod = 0
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ lvoff = -1.4226682e-8
+ toxref = 3e-9
+ tnoimod = 0
+ pags = 2.8299487e-13
+ rbodymod = 0
+ lvsat = 0.00016
+ lvth0 = 5.1655324e-8
+ ntox = 1.0
+ pcit = -1.726418e-16
+ pclm = 1.4152454
+ cigbinv = 0.006
+ delta = 0.007595625
+ laigc = -1.4938914e-10
+ tvfbsdoff = 0.022
+ rnoia = 0
+ rnoib = 0
+ phin = 0.15
+ pkt1 = 4.9696912e-14
+ pkt2 = 1.3351872e-15
+ pketa = -3.7835355e-14
+ version = 4.5
+ ngate = 8e+20
+ ltvoff = -2.0733557e-10
+ ngcon = 1
+ tempmod = 0
+ wpclm = -1.3730014e-7
+ wpdiblc2 = -4.8108443e-11
+ gbmin = 1e-12
+ rbdb = 50
+ pua1 = 6.0905252e-22
+ prwb = 0
+ prwg = 0
+ pub1 = -5.972215799999999e-31
+ jswgd = 1.28e-13
+ puc1 = 1.7562426e-23
+ jswgs = 1.28e-13
+ rbpb = 50
+ rbpd = 50
+ aigbacc = 0.02
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ pute = 3.9602525e-13
+ lku0we = 2.5e-11
+ rdsw = 100
+ wvfbsdoff = 0
+ epsrox = 3.9
+ lvfbsdoff = 0
+ rdsmod = 0
+ aigbinv = 0.0163
+ igbmod = 1
+ wkvth0we = 2e-12
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ pbswgd = 0.95
+ pbswgs = 0.95
+ rshg = 15.6
+ trnqsmod = 0
+ tvoff = 0.0020267011
+ igcmod = 1
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ poxedge = 1
+ ku0we = -0.0007
+ beta0 = 13
+ tnom = 25
+ rgatemod = 0
+ leta0 = -1.6000000000000003e-9
+ binunit = 2
+ tnjtsswg = 1
+ toxe = 2.43e-9
+ paigsd = -9.9503825e-23
+ toxm = 2.43e-9
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ permod = 1
+ wags = -1.0753313e-7
+ wcit = 4.4246590999999995e-10
+ dmcgt = 0
+ tcjsw = 0.000357
+ voff = -0.11150014
+ acde = 0.4
+ voffcv = -0.16942
+ wpemod = 1
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ vsat = 103058.98
+ wint = 0
+ vth0 = 0.37184708
+ wkt1 = -4.8627253e-8
+ wkt2 = -3.7226997e-9
+ wmax = 9.0026e-6
+ aigc = 0.011783086
+ bigsd = 0.00125
+ wmin = 9.025999999999999e-7
+ wvoff = 2.3704676e-9
+ wua1 = -8.0608962e-16
+ wub1 = 8.0443355e-25
+ wuc1 = -2.8097884e-18
+ wvsat = -0.0017920539
+ wvth0 = -9.128173e-9
+ bigc = 0.001442
+ wute = -4.4497219e-7
+ wwlc = 0
+ waigc = 2.7413515e-11
+ tpbswg = 0.0009
+ njtsswg = 9
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ lketa = 3.2718606e-9
+ xtsswgd = 0.18
+ cgsl = 3.31989e-12
+ ijthsfwd = 0.01
+ cgso = 4.90562e-11
+ xtsswgs = 0.18
+ cigc = 0.000625
+ xpart = 1
+ ckappad = 0.6
+ ckappas = 0.6
+ ptvoff = 5.4992103e-16
+ pdiblc1 = 0
+ pdiblc2 = 0.018625664
+ pdiblcb = -0.3
+ waigsd = 3.0716862e-12
+ egidl = 0.29734
+ diomod = 1
+ ijthsrev = 0.01
+ pditsd = 0
+ pditsl = 0
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ cjswgd = 2.9779200000000003e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.9779200000000003e-10
+ ags = 0.9638774700000001
+ bigbacc = 0.002588
+ cjd = 0.001432992
+ cit = -7.7402473e-5
+ cjs = 0.001432992
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 9.8024918e-9
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ k2we = 5e-5
+ kvth0we = 0.00018
+ dsub = 0.75
+ dtox = 2.7e-10
+ mjswgd = 0.85
+ mjswgs = 0.85
+ pvfbsdoff = 0
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ la0 = -2.0592205e-6
+ lintnoi = -1.5e-8
+ ppdiblc2 = 2.7806803e-16
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = 0.094562725
+ tcjswg = 0.001
+ kt1 = -0.19009298
+ lk2 = -1.3154073e-8
+ kt2 = -0.051410181
+ bigbinv = 0.004953
+ llc = 0
+ vtsswgd = 4.2
+ lln = 1
+ vtsswgs = 4.2
+ lu0 = -2.0004409e-9
+ mjd = 0.26
+ lua = -2.2049077e-16
+ mjs = 0.26
+ lub = -1.5408759e-27
+ luc = 1.1211784e-18
+ lud = 0
+ pvoff = -2.8516001e-15
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 3.0846188e-13
+ eta0 = 0.3
+ nsd = 1e+20
+ pbd = 0.52
+ pat = -8.264318700000001e-9
+ pbs = 0.52
+ pk2 = -1.9754424e-15
+ cdscb = 0
+ cdscd = 0
+ etab = -0.24888148
+ pu0 = 8.7503831e-18
+ pvsat = 1.44e-11
+ prt = 0
+ pua = 2.7693259e-23
+ pub = -6.3482817e-32
+ puc = -1.7214163e-23
+ pud = 0
+ wk2we = 5e-12
+ pvth0 = 3.5603639e-15
+ drout = 0.56
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 1.3608919e-9
+ ub1 = -8.3548641e-19
+ uc1 = 2.6015633e-11
+ paigc = -9.5524673e-18
+ tpb = 0.0014
+ wa0 = -2.8614611e-7
+ ute = -0.95836072
+ wat = 0.00092088084
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -3.5722648e-9
+ voffl = 0
+ wlc = 0
+ wln = 1
+ wu0 = -2.2701464999999998e-10
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -4.3846243e-17
+ wub = 4.7661234e-26
+ wuc = -5.9424224e-18
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ a0 = 3.5070197
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ weta0 = 0
+ pkvth0we = -1.3e-19
+ at = 61490.242
+ cf = 8.15e-11
+ wetab = -1.0073378e-8
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.028085497
+ k3 = -1.8419
+ em = 1000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.016241155
+ fprout = 300
+ w0 = 0
+ ua = -1.7947198e-9
+ ub = 2.0993593e-18
+ uc = 7.4047731e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 3.4e-9
+ )

.model nch_sf_11 nmos (
+ level = 54
+ ku0we = -0.0007
+ beta0 = 13
+ wku0we = 2e-11
+ leta0 = -1.6000000000000003e-9
+ rbdb = 50
+ mobmod = 0
+ pua1 = 9.7840116e-23
+ prwb = 0
+ prwg = 0
+ pub1 = -1.2224721e-31
+ puc1 = -3.5940917e-24
+ a0 = 1.2386098
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ wtvfbsdoff = 0
+ at = 220073.87
+ cf = 8.15e-11
+ rbpb = 50
+ rbpd = 50
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.027332723
+ k3 = -1.8419
+ rbps = 50
+ em = 1000000.0
+ rbsb = 50
+ pvag = 1.2
+ ll = 0
+ lw = 0
+ u0 = 0.015741688
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ w0 = 0
+ ua = -1.9419497e-9
+ ub = 2.1613601e-18
+ uc = 9.7509556e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 3.4e-9
+ rdsw = 100
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ ijthsfwd = 0.01
+ ltvfbsdoff = 0
+ dmcgt = 0
+ tcjsw = 0.000357
+ laigsd = -9.7335958e-18
+ ijthsrev = 0.01
+ rshg = 15.6
+ njtsswg = 9
+ bigsd = 0.00125
+ ptvfbsdoff = 0
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ wvoff = -8.1064574e-9
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.014827337
+ pdiblcb = -0.3
+ wvsat = -0.0017920539
+ ppdiblc2 = 2.4623293e-15
+ tnom = 25
+ wvth0 = 1.1738105999999999e-9
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ waigc = -9.5733062e-12
+ lketa = -3.0044615e-8
+ bigbacc = 0.002588
+ xpart = 1
+ wags = 1.2540313e-6
+ kvth0we = 0.00018
+ toxref = 3e-9
+ egidl = 0.29734
+ pkvth0we = -1.3e-19
+ wcit = 1.1976377e-10
+ ags = 0.31741392
+ cjd = 0.001432992
+ cit = 0.0013334381
+ voff = -0.11121991
+ lintnoi = -1.5e-8
+ cjs = 0.001432992
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ acde = 0.4
+ dlc = 9.8024918e-9
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ k3b = 1.9326
+ vtsswgs = 4.2
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ vsat = 103058.98
+ wint = 0
+ vfbsdoff = 0.02
+ vth0 = 0.42039507
+ wkt1 = 2.0388643e-8
+ wkt2 = -3.7425887e-9
+ wmax = 9.0026e-6
+ la0 = -4.0335612e-8
+ aigc = 0.011680759
+ wmin = 9.025999999999999e-7
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.046576700000000006
+ kt1 = -0.22273968
+ lk2 = -1.2484105e-8
+ kt2 = -0.052902736
+ llc = 0
+ lln = 1
+ lu0 = -1.5559156e-9
+ mjd = 0.26
+ ltvoff = -6.7137092e-10
+ lua = -8.9456155e-17
+ mjs = 0.26
+ lub = -5.6721601e-26
+ luc = -1.9759846e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = -3.420874e-13
+ nsd = 1e+20
+ pbd = 0.52
+ pat = -3.6322881000000003e-9
+ pbs = 0.52
+ pk2 = 6.3553328e-16
+ pvfbsdoff = 0
+ paramchk = 1
+ pu0 = 2.5098232e-17
+ wua1 = -2.3169366e-16
+ wub1 = 2.7075449e-25
+ prt = 0
+ wuc1 = 2.096158e-17
+ pua = -3.3732216e-24
+ pub = 1.7089792e-32
+ puc = 7.8894695e-24
+ pud = 0
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 9.9427719e-10
+ bigc = 0.001442
+ ub1 = -5.7879508e-19
+ uc1 = 6.536871e-11
+ pvoff = 6.4728631e-15
+ tpb = 0.0014
+ wwlc = 0
+ wa0 = 4.4480813e-7
+ ute = -1
+ wat = -0.0042836479
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -6.5059453e-9
+ cdscb = 0
+ cdscd = 0
+ lku0we = 2.5e-11
+ wlc = 0
+ wln = 1
+ wu0 = -2.4538301999999994e-10
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -8.9400845e-18
+ wub = -4.2869787e-26
+ pvsat = 1.44e-11
+ wuc = -3.4148751e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ epsrox = 3.9
+ cdsc = 0
+ wk2we = 5e-12
+ pvth0 = -5.6084018e-15
+ drout = 0.56
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ ijthdfwd = 0.01
+ cgsl = 3.31989e-12
+ paigc = 2.3365803e-17
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ rdsmod = 0
+ nfactor = 1
+ voffl = 0
+ igbmod = 1
+ weta0 = 0
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ wetab = -1.0073378e-8
+ pbswgd = 0.95
+ pbswgs = 0.95
+ ijthdrev = 0.01
+ igcmod = 1
+ cgidl = 0.22
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ lpdiblc2 = 2.7646188e-9
+ nigbacc = 10
+ k2we = 5e-5
+ pbswd = 0.8
+ pbsws = 0.8
+ dsub = 0.75
+ dtox = 2.7e-10
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ nigbinv = 10
+ paigsd = 8.7660773e-23
+ eta0 = 0.3
+ pdits = 0
+ etab = -0.24888148
+ cigsd = 0.069865
+ lkvth0we = -2e-12
+ permod = 1
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ pk2we = -1e-19
+ fnoimod = 1
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ acnqsmod = 0
+ eigbinv = 1.1
+ voffcv = -0.16942
+ wpemod = 1
+ tnoia = 0
+ rbodymod = 0
+ peta0 = 0.0
+ wketa = -4.0591301e-8
+ tpbsw = 0.0019
+ cjswd = 8.6592e-11
+ cjsws = 8.6592e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ cigbacc = 0.32875
+ wpdiblc2 = -2.5023346e-9
+ tnoimod = 0
+ tpbswg = 0.0009
+ cigbinv = 0.006
+ scref = 1e-6
+ ptvoff = 2.4706364e-16
+ pigcd = 2.621
+ keta = -0.026640801
+ aigsd = 0.010772879
+ waigsd = 3.0714759e-12
+ version = 4.5
+ lvoff = -1.4476081e-8
+ lags = 5.1202402e-7
+ wkvth0we = 2e-12
+ tempmod = 0
+ jswd = 1.28e-13
+ diomod = 1
+ jsws = 1.28e-13
+ lcit = -1.1390653e-10
+ lvsat = 0.00016
+ kt1l = 0
+ lvth0 = 8.4476154e-9
+ pditsd = 0
+ pditsl = 0
+ trnqsmod = 0
+ cjswgd = 2.9779200000000003e-10
+ tvfbsdoff = 0.022
+ pku0we = -1.5e-18
+ cjswgs = 2.9779200000000003e-10
+ delta = 0.007595625
+ laigc = -5.8318716e-11
+ aigbacc = 0.02
+ lint = 6.5375218e-9
+ rnoia = 0
+ rnoib = 0
+ lkt1 = -1.6721753e-8
+ lkt2 = -1.1643768e-8
+ lmax = 8.9908e-7
+ lmin = 4.4908e-7
+ pketa = 3.1782283e-14
+ mjswgd = 0.85
+ lpe0 = 9.2e-8
+ ngate = 8e+20
+ mjswgs = 0.85
+ lpeb = 2.5e-7
+ ngcon = 1
+ wpclm = -1.3730014e-7
+ aigbinv = 0.0163
+ tcjswg = 0.001
+ minv = -0.3
+ rgatemod = 0
+ lua1 = -1.1368255e-16
+ lub1 = 3.4544732e-26
+ luc1 = 4.1671397e-18
+ gbmin = 1e-12
+ tnjtsswg = 1
+ ndep = 1e+18
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ lwlc = 0
+ moin = 5.1
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ nigc = 3.083
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ poxedge = 1
+ fprout = 300
+ xrcrg1 = 12
+ xrcrg2 = 1
+ pags = -9.2879744e-13
+ ntox = 1.0
+ pcit = 1.1456310000000002e-16
+ binunit = 2
+ pclm = 1.4152454
+ tvoff = 0.0025480892
+ wtvoff = -5.5551488e-10
+ xjbvd = 1
+ phin = 0.15
+ xjbvs = 1
+ lk2we = -1.5e-12
+ pkt1 = -1.1727235e-14
+ pkt2 = 1.3528884e-15
+ capmod = 2
+ )

.model nch_sf_12 nmos (
+ level = 54
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ ptvfbsdoff = 0
+ cigbacc = 0.32875
+ laigsd = -9.015225e-17
+ wkvth0we = 2e-12
+ tnoia = 0
+ tnoimod = 0
+ trnqsmod = 0
+ peta0 = 0.0
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ wketa = 1.7936379e-8
+ tpbsw = 0.0019
+ a0 = 1.7327189
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ cigbinv = 0.006
+ at = 153009.14
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.020841707
+ k3 = -1.8419
+ em = 1000000.0
+ cjswd = 8.6592e-11
+ ll = -1.18e-13
+ cjsws = 8.6592e-11
+ lw = 0
+ u0 = 0.013635621
+ w0 = 0
+ mjswd = 0.11
+ ua = -2.1226101e-9
+ ub = 2.1428106e-18
+ uc = 6.8443458e-11
+ ud = 0
+ mjsws = 0.11
+ agidl = 9.41e-8
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 3.4e-9
+ k2we = 5e-5
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ dsub = 0.75
+ dtox = 2.7e-10
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ version = 4.5
+ rgatemod = 0
+ tnjtsswg = 1
+ tempmod = 0
+ eta0 = 0.3
+ etab = -0.24888148
+ aigbacc = 0.02
+ scref = 1e-6
+ pigcd = 2.621
+ aigsd = 0.010772879
+ toxref = 3e-9
+ lvoff = -6.0751145e-9
+ aigbinv = 0.0163
+ lvsat = 0.00016
+ lvth0 = -4.541492e-9
+ tvfbsdoff = 0.022
+ delta = 0.007595625
+ laigc = -1.9233809e-11
+ rnoia = 0
+ rnoib = 0
+ ltvoff = -1.0250882e-10
+ pketa = 6.0301037e-15
+ ngate = 8e+20
+ ngcon = 1
+ wpclm = -2.8227848e-7
+ poxedge = 1
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ lku0we = 2.5e-11
+ wvfbsdoff = 0
+ epsrox = 3.9
+ lvfbsdoff = 0
+ binunit = 2
+ rdsmod = 0
+ ijthsfwd = 0.01
+ igbmod = 1
+ keta = -0.041938217
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ lags = 4.5664516e-7
+ pbswgd = 0.95
+ pbswgs = 0.95
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 1.7714929e-10
+ ijthsrev = 0.01
+ igcmod = 1
+ kt1l = 0
+ tvoff = 0.0012552207
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ lint = 9.7879675e-9
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ lkt1 = -9.8358544e-9
+ lkt2 = -3.7159363e-9
+ lmax = 4.4908e-7
+ lmin = 2.1577e-7
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ ku0we = -0.0007
+ paigsd = 8.167794e-23
+ ppdiblc2 = -2.773275e-15
+ beta0 = 13
+ minv = -0.3
+ lua1 = -3.2594611e-17
+ lub1 = -2.5000430000000002e-26
+ leta0 = -1.6000000000000003e-9
+ luc1 = -3.5163101e-18
+ ndep = 1e+18
+ ppclm = 6.379047e-14
+ lwlc = 0
+ permod = 1
+ moin = 5.1
+ dlcig = 2.5e-9
+ nigc = 3.083
+ bgidl = 2320000000.0
+ njtsswg = 9
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ pkvth0we = -1.3e-19
+ dmcgt = 0
+ voffcv = -0.16942
+ ckappad = 0.6
+ wpemod = 1
+ ckappas = 0.6
+ tcjsw = 0.000357
+ pdiblc1 = 0
+ pdiblc2 = 0.026288388
+ pags = 8.4375107e-13
+ pdiblcb = -0.3
+ ntox = 1.0
+ pcit = -5.0892012e-17
+ pclm = 1.5752657
+ vfbsdoff = 0.02
+ phin = 0.15
+ bigsd = 0.00125
+ pkt1 = -6.5348923e-16
+ pkt2 = -1.2933793e-15
+ bigbacc = 0.002588
+ wvoff = 1.1413397999999999e-8
+ paramchk = 1
+ wvsat = -0.0017920539
+ kvth0we = 0.00018
+ wvth0 = -1.6974895999999998e-8
+ tpbswg = 0.0009
+ rbdb = 50
+ pua1 = 1.9082335e-23
+ prwb = 0
+ prwg = 0
+ pub1 = -2.2998905000000002e-32
+ puc1 = -7.9472634e-24
+ waigc = 5.7897385e-11
+ lintnoi = -1.5e-8
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ rdsw = 100
+ ags = 0.44327497
+ lketa = -2.3313752e-8
+ ijthdfwd = 0.01
+ ptvoff = -1.6297696e-16
+ xpart = 1
+ cjd = 0.001432992
+ cit = 0.00067194759
+ cjs = 0.001432992
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ waigsd = 3.0714895e-12
+ dlc = 1.30529375e-8
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ egidl = 0.29734
+ diomod = 1
+ la0 = -2.5774361e-7
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.017068219
+ pditsd = 0
+ pditsl = 0
+ kt1 = -0.23838945
+ ijthdrev = 0.01
+ lk2 = -9.6280577e-9
+ kt2 = -0.070920535
+ cjswgd = 2.9779200000000003e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.9779200000000003e-10
+ llc = -1.18e-13
+ lln = 0.7
+ rshg = 15.6
+ lu0 = -6.2924579e-10
+ mjd = 0.26
+ lua = -9.9655811e-18
+ mjs = 0.26
+ lub = -4.8559819e-26
+ luc = -6.9707629e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 9.4027643e-14
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 2.5627516999999998e-9
+ lpdiblc2 = -2.2782436e-9
+ pbs = 0.52
+ pk2 = 9.5548939e-17
+ pu0 = 6.9677938e-18
+ prt = 0
+ pua = -7.1355685e-24
+ pub = 6.4921301e-33
+ puc = 2.8995668e-24
+ pud = 0
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 8.0998641e-10
+ ub1 = -4.4346517e-19
+ uc1 = 8.2831095e-11
+ mjswgd = 0.85
+ mjswgs = 0.85
+ tpb = 0.0014
+ wa0 = -5.4636242e-7
+ nfactor = 1
+ pvfbsdoff = 0
+ ute = -1
+ wat = -0.018363284
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -5.2787082e-9
+ tcjswg = 0.001
+ wlc = 0
+ wln = 1
+ wu0 = -2.0417747999999998e-10
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -3.8929611e-19
+ wub = -1.8784192e-26
+ wuc = -2.2808063e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ tnom = 25
+ pvoff = -2.1158734e-15
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ cdscb = 0
+ cdscd = 0
+ lkvth0we = -2e-12
+ pvsat = 1.44e-11
+ wk2we = 5e-12
+ pvth0 = 2.3770293e-15
+ drout = 0.56
+ paigc = -6.3213007e-18
+ nigbacc = 10
+ voffl = 0
+ acnqsmod = 0
+ wags = -2.7744881e-6
+ fprout = 300
+ weta0 = 0
+ wetab = -1.0073378e-8
+ wcit = 4.9579813e-10
+ xrcrg1 = 12
+ xrcrg2 = 1
+ lpclm = -7.0408907e-8
+ voff = -0.13031302
+ rbodymod = 0
+ nigbinv = 10
+ acde = 0.4
+ cgidl = 0.22
+ vsat = 103058.98
+ wtvoff = 3.7639557e-10
+ wint = 0
+ vth0 = 0.44991577
+ wkt1 = -4.7789615999999995e-9
+ wkt2 = 2.2716562e-9
+ wmax = 9.0026e-6
+ wtvfbsdoff = 0
+ aigc = 0.01159193
+ wmin = 9.025999999999999e-7
+ capmod = 2
+ pbswd = 0.8
+ pbsws = 0.8
+ ltvfbsdoff = 0
+ fnoimod = 1
+ wua1 = -5.2698704e-17
+ wub1 = 4.5190152e-26
+ wku0we = 2e-11
+ wuc1 = 3.0855152e-17
+ eigbinv = 1.1
+ wpdiblc2 = 9.3967661e-9
+ bigc = 0.001442
+ mobmod = 0
+ wwlc = 0
+ pdits = 0
+ cigsd = 0.069865
+ cdsc = 0
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ )

.model nch_sf_13 nmos (
+ level = 54
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ lint = 9.7879675e-9
+ bigsd = 0.00125
+ lkt1 = -3.8611259999999994e-9
+ lkt2 = -5.6046527e-10
+ lmax = 2.1577e-7
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ lmin = 9e-8
+ wvoff = -2.553608e-9
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ wvsat = -0.00035982647999999954
+ minv = -0.3
+ wvth0 = -3.4626170000000013e-9
+ lua1 = 8.0644671e-18
+ lub1 = -5.0360301e-26
+ luc1 = -4.6427809e-18
+ ags = 2.6074682
+ ndep = 1e+18
+ waigc = 3.6164887e-11
+ cjd = 0.001432992
+ cit = 0.0010410649
+ cjs = 0.001432992
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ lwlc = 0
+ dlc = 1.30529375e-8
+ k3b = 1.9326
+ moin = 5.1
+ lkvth0we = -2e-12
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ nigc = 3.083
+ lketa = -1.0074554e-8
+ xpart = 1
+ la0 = -3.95931149e-8
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.0017960989
+ toxref = 3e-9
+ kt1 = -0.26670569
+ lk2 = -2.2996724e-9
+ kt2 = -0.085875374
+ llc = -1.18e-13
+ lln = 0.7
+ a0 = 0.69883298
+ a1 = 0
+ a2 = 1
+ lu0 = -2.0339706e-10
+ b0 = 0
+ b1 = 0
+ acnqsmod = 0
+ mjd = 0.26
+ lua = 2.3685126e-17
+ mjs = 0.26
+ lub = -3.581049857e-26
+ luc = -1.971816e-18
+ lud = 0
+ at = 80629.42
+ cf = 8.15e-11
+ lwc = 0
+ noff = 2.7195
+ lwl = 0
+ lwn = 1
+ ef = 1.0
+ k1 = 0.274
+ k2 = -0.013889977
+ k3 = -1.8419
+ em = 1000000.0
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ njd = 1.02
+ njs = 1.02
+ nfactor = 1
+ pa0 = 5.1229998e-14
+ egidl = 0.29734
+ ll = -1.18e-13
+ lw = 0
+ u0 = 0.01161738
+ w0 = 0
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 8.359756599999999e-10
+ pbs = 0.52
+ ua = -2.2820921e-9
+ ub = 2.0823870489000003e-18
+ uc = 4.4751766e-11
+ ud = 0
+ pk2 = 1.6389978e-16
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 3.4e-9
+ pu0 = -2.3741017e-17
+ prt = 0
+ pua = 6.5907354e-24
+ pub = -1.1536808500000001e-32
+ puc = -4.2264406e-24
+ pud = 0
+ pags = -3.4153056e-19
+ rbodymod = 0
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 6.1728936e-10
+ ub1 = -3.2327621e-19
+ uc1 = 8.8169819e-11
+ ntox = 1.0
+ pcit = -4.8109378000000005e-17
+ pclm = 1.3619854
+ tpb = 0.0014
+ wa0 = -3.4353242e-7
+ ute = -1
+ wat = -0.010179511
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -5.6026458e-9
+ wlc = 0
+ wln = 1
+ wu0 = -5.8638093e-11
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -6.5442869e-17
+ wub = 6.6660889e-26
+ wuc = 1.0964484e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ ltvoff = 4.8985213e-12
+ phin = 0.15
+ pvfbsdoff = 0
+ nigbacc = 10
+ pkt1 = 2.6483122e-15
+ pkt2 = -3.7226831e-16
+ wpdiblc2 = -7.3538749e-9
+ lku0we = 2.5e-11
+ pvoff = 8.3114947e-16
+ rbdb = 50
+ pua1 = -3.4072796e-24
+ prwb = 0
+ prwg = 0
+ pub1 = 3.9249133e-33
+ epsrox = 3.9
+ puc1 = 3.7978198e-24
+ cdscb = 0
+ cdscd = 0
+ rbpb = 50
+ rbpd = 50
+ nigbinv = 10
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ pvsat = -2.8779949e-10
+ wk2we = 5e-12
+ pvth0 = -4.740435999999999e-16
+ rdsw = 100
+ drout = 0.56
+ rdsmod = 0
+ igbmod = 1
+ paigc = -1.7357437e-18
+ voffl = 0
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ pbswgd = 0.95
+ pbswgs = 0.95
+ weta0 = 0
+ wetab = -1.0073378e-8
+ wkvth0we = 2e-12
+ fnoimod = 1
+ lpclm = -2.540677e-8
+ igcmod = 1
+ eigbinv = 1.1
+ rshg = 15.6
+ trnqsmod = 0
+ cgidl = 0.22
+ pbswd = 0.8
+ pbsws = 0.8
+ paigsd = -5.1229584e-23
+ rgatemod = 0
+ tnom = 25
+ cigbacc = 0.32875
+ tnjtsswg = 1
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ permod = 1
+ pdits = 0
+ cigsd = 0.069865
+ tnoimod = 0
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ cigbinv = 0.006
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ wags = 1.2243337999999999e-6
+ voffcv = -0.16942
+ wpemod = 1
+ wcit = 4.826102800000001e-10
+ tnoia = 0
+ voff = -0.1572150866
+ version = 4.5
+ acde = 0.4
+ tempmod = 0
+ peta0 = 0.0
+ vsat = 102561.23895
+ wint = 0
+ vth0 = 0.4644123399
+ wketa = 1.0437078e-7
+ wkt1 = -2.0427309999999998e-8
+ wkt2 = -2.0937989e-9
+ tpbsw = 0.0019
+ wmax = 9.0026e-6
+ aigc = 0.011522737
+ wmin = 9.025999999999999e-7
+ cjswd = 8.6592e-11
+ aigbacc = 0.02
+ cjsws = 8.6592e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ wua1 = 5.3887147e-17
+ wub1 = -8.2410881e-26
+ wuc1 = -2.4808749e-17
+ tpbswg = 0.0009
+ bigc = 0.001442
+ wwlc = 0
+ aigbinv = 0.0163
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ ptvoff = 8.9623963e-17
+ ijthsfwd = 0.01
+ scref = 1e-6
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ waigsd = 3.0721194e-12
+ pigcd = 2.621
+ aigsd = 0.010772879
+ diomod = 1
+ lvoff = -3.987924600000001e-10
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 2.9779200000000003e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.9779200000000003e-10
+ lvsat = 0.00026503966000000003
+ tvfbsdoff = 0.022
+ ijthsrev = 0.01
+ lvth0 = -7.60025498e-9
+ poxedge = 1
+ delta = 0.007595625
+ laigc = -4.6341008e-12
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ binunit = 2
+ rnoia = 0
+ rnoib = 0
+ mjswgd = 0.85
+ mjswgs = 0.85
+ k2we = 5e-5
+ pketa = -1.2207451e-14
+ tcjswg = 0.001
+ ngate = 8e+20
+ dsub = 0.75
+ ngcon = 1
+ dtox = 2.7e-10
+ wpclm = -2.3899735e-8
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ ppdiblc2 = 7.6111026e-16
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ eta0 = 0.3
+ etab = -0.24888148
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ fprout = 300
+ wtvfbsdoff = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ pkvth0we = -1.3e-19
+ ltvfbsdoff = 0
+ wtvoff = -8.2076521e-10
+ tvoff = 0.00074618122
+ vfbsdoff = 0.02
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ capmod = 2
+ njtsswg = 9
+ wku0we = 2e-11
+ paramchk = 1
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ ku0we = -0.0007
+ mobmod = 0
+ beta0 = 13
+ leta0 = -1.6000000000000003e-9
+ ckappad = 0.6
+ ptvfbsdoff = 0
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.022446923
+ pdiblcb = -0.3
+ ppclm = 9.2725546e-15
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ ijthdfwd = 0.01
+ keta = -0.10468292
+ bigbacc = 0.002588
+ laigsd = 3.9592657e-17
+ lags = 3.7696529e-13
+ dmcgt = 0
+ tcjsw = 0.000357
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 9.9265533e-11
+ kvth0we = 0.00018
+ ijthdrev = 0.01
+ kt1l = 0
+ lintnoi = -1.5e-8
+ lpdiblc2 = -1.4676946e-9
+ bigbinv = 0.004953
+ )

.model nch_sf_14 nmos (
+ level = 54
+ poxedge = 1
+ binunit = 2
+ scref = 1e-6
+ toxref = 3e-9
+ pigcd = 2.621
+ aigsd = 0.010772879
+ wags = 1.2243302e-6
+ lvoff = -2.035806880000001e-9
+ pkvth0we = -1.3e-19
+ wcit = 1.1125736e-10
+ tvfbsdoff = 0.022
+ voff = -0.13980004150000003
+ lvsat = 0.0016675818900000004
+ lvth0 = 2.63756691e-9
+ acde = 0.4
+ delta = 0.007595625
+ vsat = 87640.57610000002
+ laigc = -2.2637509e-11
+ wint = 0
+ vfbsdoff = 0.02
+ vth0 = 0.3554993353
+ ltvoff = 1.2509019e-10
+ wkt1 = 8.639080600000001e-8
+ wkt2 = 1.6147625e-8
+ rnoia = 0
+ rnoib = 0
+ wmax = 9.0026e-6
+ aigc = 0.011714263
+ wmin = 9.025999999999999e-7
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ pketa = 8.4378567e-15
+ ngate = 8e+20
+ paramchk = 1
+ ngcon = 1
+ wpclm = 3.4675908e-7
+ wua1 = -1.154179e-16
+ wub1 = 3.1505286e-27
+ wuc1 = 9.7519251e-17
+ lku0we = 2.5e-11
+ a0 = -0.035582299999999956
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ bigc = 0.001442
+ gbmin = 1e-12
+ epsrox = 3.9
+ at = 65883.509
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = -0.032987969000000006
+ k3 = -1.8419
+ wvfbsdoff = 0
+ em = 1000000.0
+ wwlc = 0
+ jswgd = 1.28e-13
+ lvfbsdoff = 0
+ jswgs = 1.28e-13
+ ll = 0
+ lw = 0
+ u0 = 0.0081965756
+ w0 = 0
+ ua = -2.421907e-9
+ ub = 1.9130826320999997e-18
+ uc = 4.338735e-12
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 3.4e-9
+ rdsmod = 0
+ cdsc = 0
+ igbmod = 1
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ ijthdfwd = 0.01
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ pbswgd = 0.95
+ pbswgs = 0.95
+ njtsswg = 9
+ igcmod = 1
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ ijthdrev = 0.01
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.006833075
+ pdiblcb = -0.3
+ tvoff = -0.00053245355
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ lpdiblc2 = 7.1362462e-15
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ k2we = 5e-5
+ paigsd = 1.5255572e-23
+ dsub = 0.75
+ dtox = 2.7e-10
+ ku0we = -0.0007
+ bigbacc = 0.002588
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ beta0 = 13
+ leta0 = 1.0128653999999998e-9
+ letab = -2.2297043e-8
+ permod = 1
+ kvth0we = 0.00018
+ ppclm = -2.5569374e-14
+ eta0 = 0.27220356
+ etab = -0.011678893
+ lkvth0we = -2e-12
+ dlcig = 2.5e-9
+ lintnoi = -1.5e-8
+ bgidl = 2320000000.0
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ acnqsmod = 0
+ voffcv = -0.16942
+ wpemod = 1
+ dmcgt = 0
+ tcjsw = 0.000357
+ rbodymod = 0
+ bigsd = 0.00125
+ ags = 2.6074722
+ wvoff = 7.921506600000001e-9
+ cjd = 0.001432992
+ cit = 0.00030181593
+ cjs = 0.001432992
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 3.26497e-9
+ tpbswg = 0.0009
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ wvsat = -0.0092125549
+ nfactor = 1
+ wvth0 = -1.0905709099999997e-8
+ wpdiblc2 = 7.4309162e-10
+ waigc = -2.4473999e-12
+ la0 = 2.94419216e-8
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.00040998333000000003
+ kt1 = -0.41803712
+ lk2 = -5.0446112e-10
+ kt2 = -0.10268076
+ llc = 0
+ lln = 1
+ lu0 = 1.1815857e-10
+ mjd = 0.26
+ lua = 3.6827721e-17
+ mjs = 0.26
+ lub = -1.9895881809999996e-26
+ luc = 1.827009e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ ptvoff = -1.5034232e-16
+ njd = 1.02
+ njs = 1.02
+ pa0 = 7.627786000000002e-15
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 1.00227885e-9
+ pbs = 0.52
+ pk2 = 1.6131306e-16
+ waigsd = 3.0714121e-12
+ lketa = 2.8547804e-8
+ pu0 = -1.7526607e-16
+ prt = 0
+ pua = -1.4490045e-23
+ xpart = 1
+ pub = 2.3973370000000036e-34
+ puc = 4.0045874e-24
+ pud = 0
+ rsh = 17.5
+ keta = -0.51555907
+ tcj = 0.00076
+ ua1 = 9.0255397e-10
+ ub1 = -8.0270486e-19
+ uc1 = -7.4218809e-11
+ diomod = 1
+ tpb = 0.0014
+ nigbacc = 10
+ wa0 = 1.203209e-7
+ egidl = 0.29734
+ ute = -1
+ wat = -0.011948694
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -5.5751276e-9
+ pditsd = 0
+ pditsl = 0
+ wlc = 0
+ wln = 1
+ wkvth0we = 2e-12
+ wu0 = 1.5533305e-9
+ cjswgd = 2.9779200000000003e-10
+ pku0we = -1.5e-18
+ xgl = -1.09e-8
+ cjswgs = 2.9779200000000003e-10
+ xgw = 0
+ wua = 1.5882075e-16
+ wub = -5.862147e-26
+ wuc = -7.6599643e-17
+ wud = 0
+ wwc = 0
+ jswd = 1.28e-13
+ wwl = 0
+ wwn = 1
+ jsws = 1.28e-13
+ lcit = 1.6875494e-10
+ kt1l = 0
+ trnqsmod = 0
+ nigbinv = 10
+ lint = 0
+ mjswgd = 0.85
+ mjswgs = 0.85
+ lkt1 = 1.0364027999999998e-8
+ lkt2 = 1.0192413e-9
+ pvfbsdoff = 0
+ lmax = 9e-8
+ tcjswg = 0.001
+ lmin = 5.4e-8
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ minv = -0.3
+ rgatemod = 0
+ lua1 = -1.8750406e-17
+ wtvfbsdoff = 0
+ lub1 = -5.294006799999999e-27
+ luc1 = 1.062175e-17
+ pvoff = -1.5351133999999976e-16
+ tnjtsswg = 1
+ fnoimod = 1
+ ndep = 1e+18
+ eigbinv = 1.1
+ cdscb = 0
+ cdscd = 0
+ lwlc = 0
+ moin = 5.1
+ pvsat = 5.443570199999999e-10
+ wk2we = 5e-12
+ pvth0 = 2.2560707800000002e-16
+ ltvfbsdoff = 0
+ drout = 0.56
+ nigc = 3.083
+ paigc = 1.8938113e-18
+ fprout = 300
+ voffl = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ weta0 = -3.9858587e-8
+ wetab = 2.7041872e-8
+ lpclm = -8.5343289e-9
+ wtvoff = 1.7320676e-9
+ cigbacc = 0.32875
+ ntox = 1.0
+ pcit = -1.3202202999999999e-17
+ pclm = 1.1824913
+ cgidl = 0.22
+ ptvfbsdoff = 0
+ tnoimod = 0
+ phin = 0.15
+ capmod = 2
+ pkt1 = -7.3925907e-15
+ pkt2 = -2.0869621e-15
+ wku0we = 2e-11
+ cigbinv = 0.006
+ pbswd = 0.8
+ pbsws = 0.8
+ mobmod = 0
+ rbdb = 50
+ pua1 = 1.2507395e-23
+ prwb = 0
+ prwg = 0
+ pub1 = -4.1178592e-33
+ puc1 = -7.7010123e-24
+ version = 4.5
+ pdits = 0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ cigsd = 0.069865
+ tempmod = 0
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ rdsw = 100
+ ijthsfwd = 0.01
+ aigbacc = 0.02
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ laigsd = -1.6939346e-18
+ tnoia = 0
+ ijthsrev = 0.01
+ rshg = 15.6
+ peta0 = 3.7467072e-15
+ aigbinv = 0.0163
+ petab = -3.4888335e-15
+ wketa = -1.1526014e-7
+ tpbsw = 0.0019
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ cjswd = 8.6592e-11
+ cjsws = 8.6592e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ ppdiblc2 = -4.5980291e-21
+ tnom = 25
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ )

.model nch_sf_15 nmos (
+ level = 54
+ fnoimod = 1
+ ltvoff = -2.8596488e-10
+ eigbinv = 1.1
+ pvfbsdoff = 0
+ lku0we = 2.5e-11
+ epsrox = 3.9
+ pvoff = 8.455401999999991e-16
+ cdscb = 0
+ cdscd = 0
+ rdsmod = 0
+ cigbacc = 0.32875
+ pvsat = -2.7975772999999997e-9
+ igbmod = 1
+ wk2we = 5e-12
+ pvth0 = -6.148169999999998e-16
+ drout = 0.56
+ ijthsfwd = 0.01
+ paigc = 1.0773556e-18
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ tnoimod = 0
+ voffl = 0
+ pbswgd = 0.95
+ pbswgs = 0.95
+ keta = 0.067264197
+ cigbinv = 0.006
+ weta0 = 3.2678994e-7
+ igcmod = 1
+ wetab = -1.4667966e-7
+ lpclm = -8.0899178e-8
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 3.3511574e-10
+ ijthsrev = 0.01
+ kt1l = 0
+ cgidl = 0.22
+ version = 4.5
+ a0 = 5.6809619
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = -88751.793
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = -0.013351152
+ k3 = -1.8419
+ em = 1000000.0
+ ll = 0
+ tempmod = 0
+ lw = 0
+ lint = 0
+ u0 = 0.00071525646
+ w0 = 0
+ ua = -3.0786989e-9
+ ub = 2.197681248e-18
+ uc = -5.08518e-12
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 3.4e-9
+ lkt1 = -1.6213163e-8
+ lkt2 = 1.223943e-9
+ lmax = 5.4e-8
+ lmin = 4.5e-8
+ paigsd = -3.180948e-23
+ pbswd = 0.8
+ lpe0 = 9.2e-8
+ pbsws = 0.8
+ lpeb = 2.5e-7
+ aigbacc = 0.02
+ minv = -0.3
+ permod = 1
+ lua1 = 1.293984e-17
+ lub1 = 3.95094339e-26
+ luc1 = 1.790810823e-17
+ ndep = 1e+18
+ pdits = 0
+ lwlc = 0
+ cigsd = 0.069865
+ moin = 5.1
+ aigbinv = 0.0163
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ nigc = 3.083
+ voffcv = -0.16942
+ wpemod = 1
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ pkvth0we = -1.3e-19
+ tnoia = 0
+ ntox = 1.0
+ pcit = 8.745740299999999e-17
+ pclm = 2.4301611
+ peta0 = -1.7518907e-14
+ petab = 6.5870154e-15
+ vfbsdoff = 0.02
+ wketa = 1.9475197e-7
+ poxedge = 1
+ tpbsw = 0.0019
+ phin = 0.15
+ cjswd = 8.6592e-11
+ cjsws = 8.6592e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ binunit = 2
+ pkt1 = 1.276018e-14
+ pkt2 = 7.7933247e-16
+ tpbswg = 0.0009
+ paramchk = 1
+ rbdb = 50
+ pua1 = -3.7208869e-24
+ prwb = 0
+ prwg = 0
+ pub1 = -6.899657900000001e-32
+ puc1 = -1.9085691e-23
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ ptvoff = 3.472697e-16
+ waigsd = 3.0722235e-12
+ rdsw = 100
+ ijthdfwd = 0.01
+ scref = 1e-6
+ diomod = 1
+ pigcd = 2.621
+ aigsd = 0.010772879
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ pditsd = 0
+ pditsl = 0
+ lvoff = -3.6819500800000004e-9
+ cjswgd = 2.9779200000000003e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.9779200000000003e-10
+ tvfbsdoff = 0.022
+ lvsat = 0.00203043379
+ ijthdrev = 0.01
+ lvth0 = 2.8529352400000006e-9
+ rshg = 15.6
+ delta = 0.007595625
+ laigc = -2.1310273e-11
+ wtvfbsdoff = 0
+ mjswgd = 0.85
+ mjswgs = 0.85
+ rnoia = 0
+ rnoib = 0
+ tcjswg = 0.001
+ ltvfbsdoff = 0
+ pketa = -9.5428465e-15
+ ngate = 8e+20
+ ngcon = 1
+ wpclm = -1.3405624e-6
+ njtsswg = 9
+ tnom = 25
+ wvfbsdoff = 0
+ gbmin = 1e-12
+ lvfbsdoff = 0
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ jswgd = 1.28e-13
+ toxe = 2.43e-9
+ jswgs = 1.28e-13
+ toxm = 2.43e-9
+ ckappad = 0.6
+ lkvth0we = -2e-12
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.0068331981
+ pdiblcb = -0.3
+ fprout = 300
+ ptvfbsdoff = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ acnqsmod = 0
+ wags = 1.2243302e-6
+ wcit = -1.6242531e-9
+ wtvoff = -6.84745e-9
+ bigbacc = 0.002588
+ rbodymod = 0
+ voff = -0.111418263
+ acde = 0.4
+ vsat = 81384.50940000001
+ tvoff = 0.0065547027
+ kvth0we = 0.00018
+ wint = 0
+ vth0 = 0.351786088
+ wkt1 = -2.6107076e-7
+ wkt2 = -3.3271248e-8
+ xjbvd = 1
+ xjbvs = 1
+ wmax = 9.0026e-6
+ lk2we = -1.5e-12
+ capmod = 2
+ aigc = 0.011691379
+ wmin = 9.025999999999999e-7
+ lintnoi = -1.5e-8
+ bigbinv = 0.004953
+ wku0we = 2e-11
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ mobmod = 0
+ ku0we = -0.0007
+ wua1 = 1.6438006e-16
+ wub1 = 1.12174916e-24
+ wuc1 = 2.9380698399999997e-16
+ beta0 = 13
+ wpdiblc2 = 7.4301235e-10
+ leta0 = -1.4988938100000002e-9
+ letab = 3.9727723e-8
+ bigc = 0.001442
+ wwlc = 0
+ ppclm = 7.229527e-14
+ cdsc = 0
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ laigsd = 3.532034e-18
+ dmcgt = 0
+ wkvth0we = 2e-12
+ tcjsw = 0.000357
+ nfactor = 1
+ ags = 2.6074722
+ trnqsmod = 0
+ cjd = 0.001432992
+ cit = -0.0025664738
+ cjs = 0.001432992
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ dlc = 3.26497e-9
+ k3b = 1.9326
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ bigsd = 0.00125
+ k2we = 5e-5
+ wvoff = -9.303523999999996e-9
+ la0 = -3.0211764e-7
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = 0.0085588642
+ dsub = 0.75
+ kt1 = 0.040190302
+ lk2 = -1.6433965e-9
+ kt2 = -0.1062101
+ dtox = 2.7e-10
+ llc = 0
+ lln = 1
+ lu0 = 5.5207508e-10
+ mjd = 0.26
+ nigbacc = 10
+ lua = 7.492165e-17
+ mjs = 0.26
+ lub = -3.6402602300000003e-26
+ luc = 2.373596e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ wvsat = 0.048407002000000005
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ njd = 1.02
+ njs = 1.02
+ pa0 = -1.230232e-13
+ rgatemod = 0
+ wvth0 = 3.584367999999999e-9
+ nsd = 1e+20
+ pbd = 0.52
+ pat = -8.0927789e-9
+ pbs = 0.52
+ pk2 = 5.8185614e-16
+ tnjtsswg = 1
+ pu0 = -8.3586575e-17
+ prt = 0
+ pua = 3.4306982e-23
+ pub = -6.0757564e-32
+ puc = -7.1571349e-24
+ pud = 0
+ waigc = 1.1629424e-11
+ eta0 = 0.31550975
+ rsh = 17.5
+ etab = -1.0810714
+ tcj = 0.00076
+ ua1 = 3.5617042e-10
+ ub1 = -1.575178019e-18
+ uc1 = -1.9984569999999999e-10
+ tpb = 0.0014
+ wa0 = 2.372924e-6
+ ute = -1
+ wat = 0.14486265
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -1.282587e-8
+ nigbinv = 10
+ lketa = -5.2559457e-9
+ toxref = 3e-9
+ wlc = 0
+ wln = 1
+ wu0 = -2.7350354e-11
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -6.825073e-16
+ wub = 9.9305604e-25
+ wuc = 1.1584384e-16
+ wud = 0
+ wwc = 0
+ xpart = 1
+ wwl = 0
+ wwn = 1
+ egidl = 0.29734
+ )

.model nch_sf_16 nmos (
+ level = 54
+ pketa = 8.7750313e-15
+ pkt1 = -1.1108479599999999e-15
+ pkt2 = 1.5926682e-15
+ ngate = 8e+20
+ lku0we = 2.5e-11
+ ngcon = 1
+ wpclm = -1.03603352e-6
+ epsrox = 3.9
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ wpdiblc2 = 7.4301235e-10
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ rdsmod = 0
+ bigbacc = 0.002588
+ rbdb = 50
+ pua1 = -1.9060214e-23
+ prwb = 0
+ prwg = 0
+ pub1 = 4.8648331000000004e-32
+ puc1 = 2.02154738e-23
+ igbmod = 1
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ rdsw = 100
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ kvth0we = 0.00018
+ pbswgd = 0.95
+ pbswgs = 0.95
+ lintnoi = -1.5e-8
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ igcmod = 1
+ wkvth0we = 2e-12
+ rshg = 15.6
+ trnqsmod = 0
+ tvoff = 0.002919136
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ paigsd = 4.3875156e-23
+ ku0we = -0.0007
+ permod = 1
+ beta0 = 13
+ rgatemod = 0
+ leta0 = 1.4143207e-8
+ tnom = 25
+ letab = 3.0329695e-8
+ tnjtsswg = 1
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ nfactor = 1
+ ppclm = 5.7373356e-14
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ voffcv = -0.16942
+ wpemod = 1
+ a0 = 3.2177147
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 125884.31
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.026615951000000002
+ k3 = -1.8419
+ em = 1000000.0
+ ll = 0
+ lw = 0
+ ags = 2.6074722
+ u0 = 0.0051989103
+ w0 = 0
+ ua = -2.19661343e-9
+ ub = 1.4860819409999996e-18
+ uc = 2.2595638e-10
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ wags = 1.2243302e-6
+ xl = 4e-9
+ ww = 0
+ xw = 3.4e-9
+ cjd = 0.001432992
+ cit = -0.0038023049
+ cjs = 0.001432992
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dmcgt = 0
+ dlc = 3.26497e-9
+ wcit = 3.3004264e-9
+ tcjsw = 0.000357
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ nigbacc = 10
+ voff = -0.04075972859999999
+ acde = 0.4
+ la0 = -1.8141853e-7
+ vsat = 70170.28169999999
+ wint = 0
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.0019583049
+ vth0 = 0.35751746059999995
+ kt1 = -0.20813859
+ lk2 = -3.6017846e-9
+ kt2 = -0.11042259
+ llc = 0
+ lln = 1
+ lu0 = 3.3237593e-10
+ wkt1 = 2.2011446e-8
+ wkt2 = -4.9869936e-8
+ mjd = 0.26
+ bigsd = 0.00125
+ lua = 3.1699464000000005e-17
+ mjs = 0.26
+ lub = -1.5342368999999952e-27
+ luc = -8.94744e-18
+ lud = 0
+ wmax = 9.0026e-6
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ aigc = 0.011397597
+ wmin = 9.025999999999999e-7
+ njs = 1.02
+ pa0 = -1.9996651e-13
+ nsd = 1e+20
+ nigbinv = 10
+ pbd = 0.52
+ pat = 1.734101e-10
+ pbs = 0.52
+ pk2 = 3.3250012e-16
+ tpbswg = 0.0009
+ pu0 = -1.08255347e-16
+ prt = 0
+ pua = 2.7971342e-23
+ pub = -4.5926045000000006e-32
+ puc = -7.6781524e-24
+ pud = 0
+ wvoff = 8.01398399999999e-9
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 4.3071269e-10
+ ub1 = -2.19332361e-19
+ uc1 = 5.446354900000001e-10
+ wua1 = 4.7742754e-16
+ tpb = 0.0014
+ wub1 = -1.27916739e-24
+ wuc1 = -5.08258e-16
+ wvsat = 0.057843828
+ wa0 = 3.9431957e-6
+ wvth0 = -1.3615896999999985e-8
+ ute = -1
+ wat = -0.023835087
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -7.7369724e-9
+ bigc = 0.001442
+ wlc = 0
+ wln = 1
+ wu0 = 4.7609764e-10
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -5.5320853e-16
+ wub = 6.903720200000001e-25
+ wuc = 1.2647685e-16
+ wud = 0
+ wwlc = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ waigc = -9.3979847e-11
+ ptvoff = -3.4317401e-17
+ waigsd = 3.0706789e-12
+ fnoimod = 1
+ cdsc = 0
+ eigbinv = 1.1
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ lketa = -2.4929909e-8
+ xtis = 3
+ ijthsfwd = 0.01
+ diomod = 1
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ xpart = 1
+ wtvfbsdoff = 0
+ cigc = 0.000625
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 2.9779200000000003e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.9779200000000003e-10
+ egidl = 0.29734
+ ltvfbsdoff = 0
+ ijthsrev = 0.01
+ mjswgd = 0.85
+ mjswgs = 0.85
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ cigbacc = 0.32875
+ pvfbsdoff = 0
+ tcjswg = 0.001
+ tnoimod = 0
+ k2we = 5e-5
+ dsub = 0.75
+ dtox = 2.7e-10
+ ptvfbsdoff = 0
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ cigbinv = 0.006
+ pvoff = -3.0173800000002723e-18
+ cdscb = 0
+ cdscd = 0
+ eta0 = -0.003716791
+ etab = -0.88927493
+ pvsat = -3.2599810500000005e-9
+ wk2we = 5e-12
+ pvth0 = 2.2799515999999984e-16
+ drout = 0.56
+ version = 4.5
+ fprout = 300
+ paigc = 6.2522098e-18
+ tempmod = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ voffl = 0
+ weta0 = 2.2378028e-8
+ pkvth0we = -1.3e-19
+ wetab = 3.831648e-8
+ aigbacc = 0.02
+ wtvoff = 9.4004181e-10
+ lpclm = -7.043921000000001e-8
+ cgidl = 0.22
+ vfbsdoff = 0.02
+ capmod = 2
+ aigbinv = 0.0163
+ wku0we = 2e-11
+ mobmod = 0
+ pbswd = 0.8
+ pbsws = 0.8
+ paramchk = 1
+ pdits = 0
+ cigsd = 0.069865
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ poxedge = 1
+ ijthdfwd = 0.01
+ laigsd = -2.6649547e-17
+ pk2we = -1e-19
+ keta = 0.46877367
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ binunit = 2
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ tnoia = 0
+ lcit = 3.9567143e-10
+ ijthdrev = 0.01
+ kt1l = 0
+ peta0 = -2.6027237e-15
+ petab = -2.4777955e-15
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ wketa = -1.7908228e-7
+ tpbsw = 0.0019
+ lint = 0
+ cjswd = 8.6592e-11
+ cjsws = 8.6592e-11
+ lkt1 = -4.045047e-9
+ lkt2 = 1.4303548e-9
+ mjswd = 0.11
+ lmax = 4.5e-8
+ mjsws = 0.11
+ agidl = 9.41e-8
+ lmin = 3.6e-8
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ minv = -0.3
+ lua1 = 9.2872684e-18
+ lub1 = -2.69270018e-26
+ luc1 = -1.8571467190000002e-17
+ ndep = 1e+18
+ lwlc = 0
+ lkvth0we = -2e-12
+ moin = 5.1
+ toxref = 3e-9
+ nigc = 3.083
+ scref = 1e-6
+ pigcd = 2.621
+ aigsd = 0.01077288
+ acnqsmod = 0
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ lvoff = -7.14421828e-9
+ tvfbsdoff = 0.022
+ njtsswg = 9
+ rbodymod = 0
+ lvsat = 0.002579933613
+ lvth0 = 2.5720960299999997e-9
+ ntox = 1.0
+ ltvoff = -1.0782211e-10
+ pcit = -1.5385171000000001e-16
+ pclm = 2.21669238
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ delta = 0.007595625
+ laigc = -6.9149623e-12
+ ckappad = 0.6
+ ckappas = 0.6
+ rnoia = 0
+ rnoib = 0
+ pdiblc1 = 0
+ pdiblc2 = 0.0068331981
+ phin = 0.15
+ pdiblcb = -0.3
+ )

.model nch_sf_17 nmos (
+ level = 54
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ pbswgd = 0.95
+ xtis = 3
+ pbswgs = 0.95
+ ijthdfwd = 0.01
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ aigbinv = 0.0163
+ cigc = 0.000625
+ voffl = 0
+ igcmod = 1
+ weta0 = -1.09928e-7
+ wetab = 2.7482e-8
+ ijthdrev = 0.01
+ cgidl = 0.22
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ poxedge = 1
+ k2we = 5e-5
+ pbswd = 0.8
+ pbsws = 0.8
+ dsub = 0.75
+ permod = 1
+ dtox = 2.7e-10
+ binunit = 2
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ pdits = 0
+ eta0 = 0.42133333
+ cigsd = 0.069865
+ etab = -0.29033333
+ lkvth0we = -2e-12
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ voffcv = -0.16942
+ wpemod = 1
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ acnqsmod = 0
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ tnoia = 0
+ rbodymod = 0
+ peta0 = 0.0
+ wketa = -3.7974654e-8
+ tpbsw = 0.0019
+ cjswd = 8.6592e-11
+ tpbswg = 0.0009
+ cjsws = 8.6592e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ wtvfbsdoff = 0
+ a0 = 2.2098167
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 72000
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.018286228
+ k3 = -1.8419
+ em = 1000000.0
+ wpdiblc2 = -6.449088e-9
+ ll = 0
+ lw = 0
+ u0 = 0.0158665
+ w0 = 0
+ ua = -1.7855187e-9
+ ub = 2.0636167e-18
+ uc = 7.8391667e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ptvoff = 0
+ ww = 0
+ xw = 3.4e-9
+ njtsswg = 9
+ ltvfbsdoff = 0
+ waigsd = 3.0876027e-12
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ diomod = 1
+ scref = 1e-6
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.025656394
+ pigcd = 2.621
+ pdiblcb = -0.3
+ pditsd = 0
+ pditsl = 0
+ aigsd = 0.010772862
+ cjswgd = 2.9779200000000003e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.9779200000000003e-10
+ keta = 0.015093331
+ tvfbsdoff = 0.022
+ lvoff = 1.6e-11
+ wkvth0we = 2e-12
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lvsat = 0.00016
+ lcit = 8e-12
+ lvth0 = 4.0000000000000007e-10
+ ptvfbsdoff = 0
+ kt1l = 0
+ mjswgd = 0.85
+ mjswgs = 0.85
+ trnqsmod = 0
+ delta = 0.007595625
+ bigbacc = 0.002588
+ tcjswg = 0.001
+ rnoia = 0
+ rnoib = 0
+ lint = 6.5375218e-9
+ kvth0we = 0.00018
+ lkt1 = -2.4e-10
+ lmax = 2.001e-5
+ lmin = 8.9991e-6
+ ngate = 8e+20
+ lintnoi = -1.5e-8
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ ngcon = 1
+ bigbinv = 0.004953
+ wpclm = 5.7423639e-7
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ rgatemod = 0
+ minv = -0.3
+ lub1 = 2.4000000000000004e-27
+ gbmin = 1e-12
+ tnjtsswg = 1
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ ndep = 1e+18
+ lwlc = 0
+ moin = 5.1
+ fprout = 300
+ nigc = 3.083
+ xrcrg1 = 12
+ xrcrg2 = 1
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ wtvoff = 9.3503662e-10
+ ntox = 1.0
+ pcit = 1.2000000000000001e-17
+ pclm = 0.629885
+ tvoff = 5.0359625e-5
+ capmod = 2
+ nfactor = 1
+ wku0we = 2e-11
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ phin = 0.15
+ mobmod = 0
+ pkt1 = -1.76e-16
+ ku0we = -0.0007
+ beta0 = 13
+ leta0 = -1.6000000000000003e-9
+ nigbacc = 10
+ rbdb = 50
+ prwb = 0
+ prwg = 0
+ pub1 = 1.6e-34
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ ags = 0.73720097
+ dlcig = 2.5e-9
+ rdsw = 100
+ bgidl = 2320000000.0
+ cjd = 0.001432992
+ cit = 6.2896875e-5
+ cjs = 0.001432992
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 9.8024918e-9
+ ijthsfwd = 0.01
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ nigbinv = 10
+ la0 = 0
+ jsd = 6.11e-7
+ dmcgt = 0
+ jss = 6.11e-7
+ lat = 8e-5
+ kt1 = -0.28314411
+ kt2 = -0.074391698
+ tcjsw = 0.000357
+ llc = 0
+ lln = 1
+ lu0 = -4e-12
+ mjd = 0.26
+ mjs = 0.26
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 0
+ ijthsrev = 0.01
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 1.44e-11
+ pbs = 0.52
+ rshg = 15.6
+ pu0 = -1.2e-18
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ prt = 0
+ pud = 0
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = -6.8749055e-10
+ ub1 = 1.0341951e-18
+ uc1 = 4.5339833e-11
+ fnoimod = 1
+ bigsd = 0.00125
+ tpb = 0.0014
+ wa0 = 7.159061e-7
+ eigbinv = 1.1
+ ute = -2.01925
+ wat = 0
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 3.760485e-9
+ wlc = 0
+ wln = 1
+ wu0 = -8.766899999999998e-11
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -7.132277e-17
+ wub = 7.28273e-26
+ wuc = -1.167985e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ wvoff = 6.981215e-10
+ wvsat = -0.0045771271
+ wvth0 = -6.3727395e-9
+ tnom = 25
+ toxe = 2.43e-9
+ waigc = 5.0140497e-11
+ toxm = 2.43e-9
+ toxref = 3e-9
+ cigbacc = 0.32875
+ xpart = 1
+ tnoimod = 0
+ wags = 1.2293247e-7
+ egidl = 0.29734
+ pkvth0we = -1.3e-19
+ wcit = 4.0907306e-10
+ cigbinv = 0.006
+ voff = -0.11158375
+ ltvoff = 0
+ acde = 0.4
+ vsat = 106133.02
+ vfbsdoff = 0.02
+ wint = 0
+ pvfbsdoff = 0
+ vth0 = 0.37492953
+ wkt1 = 3.6635480999999995e-8
+ wkt2 = 1.5939759e-8
+ wmax = 9.025999999999999e-7
+ aigc = 0.011740211
+ wmin = 5.426e-7
+ version = 4.5
+ tempmod = 0
+ lku0we = 2.5e-11
+ epsrox = 3.9
+ paramchk = 1
+ wua1 = 1.0731531e-15
+ wub1 = -9.2968455e-25
+ wuc1 = -1.4414309e-17
+ aigbacc = 0.02
+ rdsmod = 0
+ bigc = 0.001442
+ pvoff = -4e-17
+ wute = 5.565105e-7
+ wwlc = 0
+ igbmod = 1
+ cdscb = 0
+ cdscd = 0
+ pvsat = 1.44e-11
+ wk2we = 5e-12
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ pvth0 = 1.2e-16
+ cdsc = 0
+ drout = 0.56
+ )

.model nch_sf_18 nmos (
+ level = 54
+ kt1l = 0
+ nigbacc = 10
+ tvoff = -0.0002433276
+ paigsd = 1.3573222e-22
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ lint = 6.5375218e-9
+ lkt1 = 8.600640500000001e-8
+ lkt2 = 5.1456509e-9
+ lmax = 8.9991e-6
+ lmin = 8.9908e-7
+ permod = 1
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ nigbinv = 10
+ ags = 0.69161289
+ ku0we = -0.0007
+ ppdiblc2 = 1.9760389e-14
+ beta0 = 13
+ cjd = 0.001432992
+ leta0 = -1.6000000000000003e-9
+ cit = -0.00011782923
+ cjs = 0.001432992
+ minv = -0.3
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ lua1 = 1.38467e-15
+ lub1 = -1.4868591e-24
+ luc1 = 1.0686128e-16
+ dlc = 9.8024918e-9
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ ndep = 1e+18
+ lute = 1.0068051e-6
+ lwlc = 0
+ moin = 5.1
+ dlcig = 2.5e-9
+ voffcv = -0.16942
+ wpemod = 1
+ bgidl = 2320000000.0
+ la0 = -1.1479603e-6
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ nigc = 3.083
+ lat = 0.085425067
+ kt1 = -0.2927377
+ lk2 = -1.3507419e-8
+ kt2 = -0.074964073
+ llc = 0
+ lln = 1
+ lu0 = -2.0044396e-9
+ fnoimod = 1
+ mjd = 0.26
+ lua = -1.5028094e-16
+ mjs = 0.26
+ lub = -1.4426347e-25
+ luc = -5.2935673e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = -5.1713984e-13
+ eigbinv = 1.1
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 1.44e-11
+ pbs = 0.52
+ pk2 = -1.6553107e-15
+ pu0 = 1.2373224e-17
+ prt = 0
+ noff = 2.7195
+ pua = -3.5916841e-23
+ pub = 6.5823852e-32
+ puc = 3.1761344e-23
+ pud = 0
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ pkvth0we = -1.3e-19
+ dmcgt = 0
+ rsh = 17.5
+ tcjsw = 0.000357
+ tcj = 0.00076
+ ua1 = -8.4151391e-10
+ ub1 = 1.1998524e-18
+ uc1 = 3.3453151e-11
+ tpb = 0.0014
+ wa0 = 7.7343e-7
+ pags = -1.4569295e-13
+ ute = -2.1312417
+ wtvfbsdoff = 0
+ wat = 0
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 3.944613e-9
+ wlc = 0
+ wln = 1
+ ntox = 1.0
+ wu0 = -8.917881e-11
+ pcit = -6.1747523e-16
+ xgl = -1.09e-8
+ pclm = 0.629885
+ xgw = 0
+ wua = -6.7327571e-17
+ wub = 6.5505403e-26
+ wuc = -1.5212814e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ vfbsdoff = 0.02
+ tpbswg = 0.0009
+ bigsd = 0.00125
+ ltvfbsdoff = 0
+ phin = 0.15
+ cigbacc = 0.32875
+ wvoff = 5.020811499999999e-10
+ pkt1 = -6.969914000000001e-14
+ pkt2 = -1.5079533e-14
+ paramchk = 1
+ tnoimod = 0
+ wvsat = -0.0045771271
+ wvth0 = -6.6760901e-9
+ ptvoff = -2.0299898e-15
+ waigsd = 3.0875876e-12
+ waigc = 5.030718e-11
+ rbdb = 50
+ pua1 = -1.044071e-21
+ prwb = 0
+ prwg = 0
+ pub1 = 9.881508100000001e-31
+ cigbinv = 0.006
+ puc1 = -4.3746501e-23
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ pute = -5.4971558e-13
+ diomod = 1
+ rdsw = 100
+ ptvfbsdoff = 0
+ lketa = -1.3350472e-7
+ ijthdfwd = 0.01
+ pditsd = 0
+ xpart = 1
+ pditsl = 0
+ cjswgd = 2.9779200000000003e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.9779200000000003e-10
+ version = 4.5
+ tempmod = 0
+ egidl = 0.29734
+ mjswgd = 0.85
+ mjswgs = 0.85
+ ijthdrev = 0.01
+ aigbacc = 0.02
+ a0 = 2.3375097
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ rshg = 15.6
+ at = 62506.667
+ cf = 8.15e-11
+ tcjswg = 0.001
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.019788722
+ k3 = -1.8419
+ em = 1000000.0
+ pvfbsdoff = 0
+ ll = 0
+ lw = 0
+ u0 = 0.016089018
+ lpdiblc2 = -2.2119558e-8
+ w0 = 0
+ ua = -1.7688022e-9
+ ub = 2.0796638e-18
+ uc = 8.4279951e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 3.4e-9
+ aigbinv = 0.0163
+ tnom = 25
+ pvoff = 1.7224031e-15
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ cdscb = 0
+ cdscd = 0
+ fprout = 300
+ pvsat = 1.44e-11
+ lkvth0we = -2e-12
+ wk2we = 5e-12
+ pvth0 = 2.8471227e-15
+ drout = 0.56
+ xrcrg1 = 12
+ xrcrg2 = 1
+ paigc = -1.4984839e-18
+ voffl = 0
+ poxedge = 1
+ acnqsmod = 0
+ wtvoff = 1.1608419e-9
+ wags = 1.3913858999999998e-7
+ weta0 = -1.09928e-7
+ wetab = 2.7482e-8
+ wcit = 4.7909255e-10
+ binunit = 2
+ rbodymod = 0
+ voff = -0.1094379
+ acde = 0.4
+ capmod = 2
+ cgidl = 0.22
+ vsat = 106133.02
+ wint = 0
+ wku0we = 2e-11
+ vth0 = 0.36914059
+ wkt1 = 4.4368867e-8
+ wkt2 = 1.7617127e-8
+ wmax = 9.025999999999999e-7
+ mobmod = 0
+ aigc = 0.011757817
+ wmin = 5.426e-7
+ pbswd = 0.8
+ pbsws = 0.8
+ wua1 = 1.1892901e-15
+ wub1 = -1.0395834e-24
+ wuc1 = -9.5481798e-18
+ wpdiblc2 = -8.647129e-9
+ bigc = 0.001442
+ wute = 6.1765795e-7
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ wwlc = 0
+ pdits = 0
+ cigsd = 0.069865
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ laigsd = -2.4859383e-16
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ wkvth0we = 2e-12
+ tnoia = 0
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ trnqsmod = 0
+ peta0 = 0.0
+ njtsswg = 9
+ wketa = -4.7550208e-8
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ tpbsw = 0.0019
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ cjswd = 8.6592e-11
+ cjsws = 8.6592e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.028116857
+ k2we = 5e-5
+ pdiblcb = -0.3
+ dsub = 0.75
+ dtox = 2.7e-10
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ rgatemod = 0
+ tnjtsswg = 1
+ toxref = 3e-9
+ eta0 = 0.42133333
+ etab = -0.29033333
+ bigbacc = 0.002588
+ scref = 1e-6
+ pigcd = 2.621
+ aigsd = 0.010772862
+ kvth0we = 0.00018
+ tvfbsdoff = 0.022
+ lvoff = -1.9275251e-8
+ lintnoi = -1.5e-8
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ ltvoff = 2.6402481e-9
+ lvsat = 0.00016
+ lvth0 = 5.2442565999999996e-8
+ delta = 0.007595625
+ laigc = -1.5827875e-10
+ rnoia = 0
+ rnoib = 0
+ lku0we = 2.5e-11
+ pketa = 8.6084224e-14
+ epsrox = 3.9
+ ngate = 8e+20
+ ngcon = 1
+ wvfbsdoff = 0
+ wpclm = 5.7423639e-7
+ lvfbsdoff = 0
+ rdsmod = 0
+ gbmin = 1e-12
+ igbmod = 1
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ pbswgd = 0.95
+ pbswgs = 0.95
+ nfactor = 1
+ ijthsfwd = 0.01
+ igcmod = 1
+ keta = 0.029943688
+ lags = 4.0983681e-7
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 1.6327276999999999e-9
+ ijthsrev = 0.01
+ )

.model nch_sf_19 nmos (
+ level = 54
+ rgatemod = 0
+ tnom = 25
+ tnjtsswg = 1
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ pdits = 0
+ cigsd = 0.069865
+ voffcv = -0.16942
+ wpemod = 1
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ njtsswg = 9
+ wtvfbsdoff = 0
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ ltvfbsdoff = 0
+ ckappad = 0.6
+ ckappas = 0.6
+ wags = -7.75542e-7
+ pdiblc1 = 0
+ pdiblc2 = -0.019237439
+ pdiblcb = -0.3
+ wcit = -4.9548514e-10
+ tnoia = 0
+ voff = -0.12566406
+ acde = 0.4
+ peta0 = 0.0
+ vsat = 106133.02
+ wketa = 9.2259042e-8
+ wint = 0
+ tpbswg = 0.0009
+ vth0 = 0.42734179
+ tpbsw = 0.0019
+ wkt1 = -6.739324899999999e-8
+ wkt2 = 3.7202325e-9
+ wmax = 9.025999999999999e-7
+ bigbacc = 0.002588
+ cjswd = 8.6592e-11
+ aigc = 0.01160027
+ cjsws = 8.6592e-11
+ wmin = 5.426e-7
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ ptvfbsdoff = 0
+ kvth0we = 0.00018
+ ptvoff = 9.96032e-16
+ wua1 = 1.1798319e-17
+ wub1 = 1.8760115e-25
+ wuc1 = -8.2926019e-17
+ lintnoi = -1.5e-8
+ waigsd = 3.0878745e-12
+ bigbinv = 0.004953
+ bigc = 0.001442
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ wwlc = 0
+ diomod = 1
+ cdsc = 0
+ cgbo = 0
+ pditsd = 0
+ pditsl = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ cjswgd = 2.9779200000000003e-10
+ ijthsfwd = 0.01
+ scref = 1e-6
+ pku0we = -1.5e-18
+ cjswgs = 2.9779200000000003e-10
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ pigcd = 2.621
+ tvfbsdoff = 0.022
+ aigsd = 0.010772861
+ lvoff = -4.8339703e-9
+ mjswgd = 0.85
+ mjswgs = 0.85
+ lvsat = 0.00016
+ lvth0 = 6.434924000000001e-10
+ ijthsrev = 0.01
+ tcjswg = 0.001
+ delta = 0.007595625
+ laigc = -1.8062176e-11
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ rnoia = 0
+ rnoib = 0
+ nfactor = 1
+ pketa = -3.8346008e-14
+ ngate = 8e+20
+ k2we = 5e-5
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ ngcon = 1
+ dsub = 0.75
+ wpclm = 5.7423639e-7
+ dtox = 2.7e-10
+ ppdiblc2 = -1.3176269e-14
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ fprout = 300
+ eta0 = 0.42133333
+ etab = -0.29033333
+ xrcrg1 = 12
+ xrcrg2 = 1
+ nigbacc = 10
+ a0 = 1.6362276
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 209176.65
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.016538798
+ k3 = -1.8419
+ em = 1000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.015567274
+ w0 = 0
+ ua = -1.7708735e-9
+ ub = 1.8600147e-18
+ uc = 2.580063e-11
+ ud = 0
+ wtvoff = -2.2391826e-9
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 3.4e-9
+ pkvth0we = -1.3e-19
+ nigbinv = 10
+ capmod = 2
+ wku0we = 2e-11
+ tvoff = 0.004406442
+ vfbsdoff = 0.02
+ mobmod = 0
+ ags = 2.557561
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ cjd = 0.001432992
+ cit = 0.0020125208
+ cjs = 0.001432992
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 9.8024918e-9
+ k3b = 1.9326
+ fnoimod = 1
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ eigbinv = 1.1
+ paramchk = 1
+ ku0we = -0.0007
+ beta0 = 13
+ la0 = -5.2381924e-7
+ leta0 = -1.6000000000000003e-9
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.04511122
+ kt1 = -0.12585017
+ lk2 = -1.0614987e-8
+ kt2 = -0.061139846
+ llc = 0
+ lln = 1
+ lu0 = -1.5400873e-9
+ mjd = 0.26
+ lua = -1.4843753e-16
+ mjs = 0.26
+ lub = 5.1224193e-26
+ luc = -8.8907704e-19
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 9.5948774e-14
+ nsd = 1e+20
+ pbd = 0.52
+ pat = -4.9600129999999994e-9
+ pbs = 0.52
+ laigsd = 2.1900591e-16
+ pk2 = -1.0578878e-15
+ pu0 = 1.0757724e-17
+ dlcig = 2.5e-9
+ prt = 0
+ pua = 5.0063903e-23
+ pub = -8.0709098e-32
+ puc = -9.2074471e-24
+ pud = 0
+ bgidl = 2320000000.0
+ ijthdfwd = 0.01
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 7.2552224e-10
+ ub1 = -4.8701436e-19
+ uc1 = 1.8003493e-10
+ tpb = 0.0014
+ wa0 = 8.4566389e-8
+ ute = -1
+ wat = 0.0055892281
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 3.2733514e-9
+ keta = -0.17327473
+ cigbacc = 0.32875
+ wlc = 0
+ wln = 1
+ wu0 = -8.736364e-11
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -1.6393515e-16
+ wub = 2.3014917e-25
+ wuc = 3.0819536e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ dmcgt = 0
+ tcjsw = 0.000357
+ lags = -1.250857e-6
+ tnoimod = 0
+ jswd = 1.28e-13
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ jsws = 1.28e-13
+ lcit = -2.6328379999999997e-10
+ ijthdrev = 0.01
+ kt1l = 0
+ cigbinv = 0.006
+ lpdiblc2 = 2.0025765e-8
+ bigsd = 0.00125
+ lint = 6.5375218e-9
+ lkt1 = -6.2523496e-8
+ lkt2 = -7.1579117e-9
+ lmax = 8.9908e-7
+ lmin = 4.4908e-7
+ wvoff = 4.979937800000001e-9
+ lpe0 = 9.2e-8
+ version = 4.5
+ lpeb = 2.5e-7
+ tempmod = 0
+ wvsat = -0.0045771271
+ wvth0 = -5.119922700000001e-9
+ minv = -0.3
+ lua1 = -9.9922063e-18
+ lub1 = 1.4452288e-26
+ luc1 = -2.3596511e-17
+ toxref = 3e-9
+ waigc = 6.3350032e-11
+ ndep = 1e+18
+ aigbacc = 0.02
+ lwlc = 0
+ lkvth0we = -2e-12
+ moin = 5.1
+ lketa = 4.735968e-8
+ nigc = 3.083
+ xpart = 1
+ acnqsmod = 0
+ aigbinv = 0.0163
+ egidl = 0.29734
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ ltvoff = -1.4980468e-9
+ rbodymod = 0
+ pags = 6.6837277e-13
+ ntox = 1.0
+ pvfbsdoff = 0
+ pcit = 2.4989891e-16
+ pclm = 0.629885
+ phin = 0.15
+ lku0we = 2.5e-11
+ epsrox = 3.9
+ pkt1 = 2.9769144e-14
+ pkt2 = -2.7112972e-15
+ poxedge = 1
+ rdsmod = 0
+ igbmod = 1
+ wpdiblc2 = 2.8360352e-8
+ pvoff = -2.2628893999999997e-15
+ binunit = 2
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ rbdb = 50
+ pua1 = 3.8966634e-24
+ prwb = 0
+ prwg = 0
+ pub1 = -1.0404345999999999e-31
+ cdscb = 0
+ cdscd = 0
+ puc1 = 2.1559776e-23
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ pvsat = 1.44e-11
+ rbsb = 50
+ pvag = 1.2
+ pbswgd = 0.95
+ pbswgs = 0.95
+ wk2we = 5e-12
+ pvth0 = 1.4621336999999999e-15
+ drout = 0.56
+ rdsw = 100
+ igcmod = 1
+ paigc = -1.3106622e-17
+ voffl = 0
+ weta0 = -1.09928e-7
+ wetab = 2.7482e-8
+ wkvth0we = 2e-12
+ trnqsmod = 0
+ cgidl = 0.22
+ rshg = 15.6
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ paigsd = -1.1957726e-22
+ permod = 1
+ pbswd = 0.8
+ pbsws = 0.8
+ )

.model nch_sf_20 nmos (
+ level = 54
+ rgatemod = 0
+ tnom = 25
+ tnjtsswg = 1
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ pdits = 0
+ cigsd = 0.069865
+ voffcv = -0.16942
+ wpemod = 1
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ njtsswg = 9
+ wtvfbsdoff = 0
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ ltvfbsdoff = 0
+ ckappad = 0.6
+ ckappas = 0.6
+ wags = 2.522663e-6
+ pdiblc1 = 0
+ pdiblc2 = 0.041730695
+ pdiblcb = -0.3
+ wcit = 1.1646633e-10
+ tnoia = 0
+ voff = -0.11119538
+ acde = 0.4
+ peta0 = 0.0
+ vsat = 99029.765
+ wketa = 8.4379468e-9
+ wint = 0
+ tpbswg = 0.0009
+ vth0 = 0.43569989
+ tpbsw = 0.0019
+ wkt1 = 1.2876763e-8
+ wkt2 = -6.4493333e-9
+ wmax = 9.025999999999999e-7
+ bigbacc = 0.002588
+ cjswd = 8.6592e-11
+ aigc = 0.011620363
+ cjsws = 8.6592e-11
+ wmin = 5.426e-7
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ ptvfbsdoff = 0
+ kvth0we = 0.00018
+ ptvoff = -1.0913215e-16
+ wua1 = 2.6150731e-17
+ wub1 = -7.4432483e-26
+ wuc1 = -3.5091334e-17
+ lintnoi = -1.5e-8
+ waigsd = 3.0877293e-12
+ bigbinv = 0.004953
+ bigc = 0.001442
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ wwlc = 0
+ diomod = 1
+ cdsc = 0
+ cgbo = 0
+ pditsd = 0
+ pditsl = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ cjswgd = 2.9779200000000003e-10
+ ijthsfwd = 0.01
+ scref = 1e-6
+ pku0we = -1.5e-18
+ cjswgs = 2.9779200000000003e-10
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ pigcd = 2.621
+ tvfbsdoff = 0.022
+ aigsd = 0.010772861
+ lvoff = -1.120019e-8
+ mjswgd = 0.85
+ mjswgs = 0.85
+ lvsat = 0.0032854309
+ lvth0 = -3.0340680000000002e-9
+ ijthsrev = 0.01
+ tcjswg = 0.001
+ delta = 0.007595625
+ laigc = -2.6902885e-11
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ rnoia = 0
+ rnoib = 0
+ nfactor = 1
+ pketa = -1.4647263e-15
+ ngate = 8e+20
+ k2we = 5e-5
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ ngcon = 1
+ dsub = 0.75
+ wpclm = 5.7423639e-7
+ dtox = 2.7e-10
+ ppdiblc2 = 1.3236303e-15
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ fprout = 300
+ eta0 = 0.42133333
+ etab = -0.29033333
+ xrcrg1 = 12
+ xrcrg2 = 1
+ nigbacc = 10
+ a0 = -0.63009793
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 152816.98
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.01550817
+ k3 = -1.8419
+ em = 1000000.0
+ ll = -1.18e-13
+ lw = 0
+ u0 = 0.013490665
+ w0 = 0
+ ua = -2.0345741e-9
+ ub = 2.0265059e-18
+ uc = 2.0750138e-11
+ ud = 0
+ wtvoff = 2.7255415e-10
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 3.4e-9
+ pkvth0we = -1.3e-19
+ nigbinv = 10
+ capmod = 2
+ wku0we = 2e-11
+ tvoff = 0.001369836
+ vfbsdoff = 0.02
+ mobmod = 0
+ ags = -5.4034702
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ cjd = 0.001432992
+ cit = 0.0010906361
+ cjs = 0.001432992
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 1.30529375e-8
+ k3b = 1.9326
+ fnoimod = 1
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ eigbinv = 1.1
+ paramchk = 1
+ ku0we = -0.0007
+ beta0 = 13
+ la0 = 4.73364e-7
+ leta0 = -1.6000000000000003e-9
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.020312964
+ kt1 = -0.257877
+ lk2 = -1.0161511e-8
+ kt2 = -0.061294719
+ llc = -1.18e-13
+ lln = 0.7
+ lu0 = -6.2637936e-10
+ mjd = 0.26
+ lua = -3.2409276e-17
+ mjs = 0.26
+ lub = -2.2031936e-26
+ luc = 1.3331392e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = -5.6835585e-13
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 5.5024901e-9
+ pbs = 0.52
+ laigsd = 6.148791e-17
+ pk2 = 5.7885716e-16
+ pu0 = 4.3708054e-18
+ dlcig = 2.5e-9
+ prt = 0
+ pua = 1.3198419e-23
+ pub = -1.7542132e-32
+ puc = -4.6237685e-24
+ pud = 0
+ bgidl = 2320000000.0
+ ijthdfwd = 0.01
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 7.2295613e-10
+ ub1 = -3.1143135e-19
+ uc1 = 1.5561971e-10
+ tpb = 0.0014
+ wa0 = 1.5943496e-6
+ ute = -1
+ wat = -0.018189188
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -4.4652352e-10
+ keta = -0.031454297
+ cigbacc = 0.32875
+ wlc = 0
+ wln = 1
+ wu0 = -7.284792e-11
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -8.0149958e-17
+ wub = 8.6587882e-26
+ wuc = 2.0402085e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ dmcgt = 0
+ tcjsw = 0.000357
+ lags = 2.2519967e-6
+ tnoimod = 0
+ jswd = 1.28e-13
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ jsws = 1.28e-13
+ lcit = 1.4234545e-10
+ ijthdrev = 0.01
+ kt1l = 0
+ cigbinv = 0.006
+ lpdiblc2 = -6.8002141e-9
+ bigsd = 0.00125
+ lint = 9.7879675e-9
+ lkt1 = -4.4316909e-9
+ lkt2 = -7.0897675e-9
+ lmax = 4.4908e-7
+ lmin = 2.1577e-7
+ wvoff = -5.9071857e-9
+ lpe0 = 9.2e-8
+ version = 4.5
+ lpeb = 2.5e-7
+ tempmod = 0
+ wvsat = 0.0018584193
+ wvth0 = -4.0953081e-9
+ minv = -0.3
+ lua1 = -8.8631172e-18
+ lub1 = -6.280423399999999e-26
+ luc1 = -1.2853813e-17
+ toxref = 3e-9
+ waigc = 3.2137522e-11
+ ndep = 1e+18
+ aigbacc = 0.02
+ lwlc = 0
+ lkvth0we = -2e-12
+ moin = 5.1
+ lketa = -1.5041313e-8
+ nigc = 3.083
+ xpart = 1
+ acnqsmod = 0
+ aigbinv = 0.0163
+ egidl = 0.29734
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ ltvoff = -1.6194017e-10
+ rbodymod = 0
+ pags = -7.8283743e-13
+ ntox = 1.0
+ pvfbsdoff = 0
+ pcit = -1.9359734999999997e-17
+ pclm = 0.629885
+ phin = 0.15
+ lku0we = 2.5e-11
+ epsrox = 3.9
+ pkt1 = -5.5496613e-15
+ pkt2 = 1.7633117e-15
+ poxedge = 1
+ rdsmod = 0
+ igbmod = 1
+ wpdiblc2 = -4.5939646e-9
+ pvoff = 2.527445e-15
+ binunit = 2
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ rbdb = 50
+ pua1 = -2.4183981e-24
+ prwb = 0
+ prwg = 0
+ pub1 = 1.1251342e-32
+ cdscb = 0
+ cdscd = 0
+ puc1 = 5.125141e-25
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ pvsat = -2.8172404000000002e-9
+ rbsb = 50
+ pvag = 1.2
+ pbswgd = 0.95
+ pbswgs = 0.95
+ wk2we = 5e-12
+ pvth0 = 1.0113032399999999e-15
+ drout = 0.56
+ rdsw = 100
+ igcmod = 1
+ paigc = 6.2688273e-19
+ voffl = 0
+ weta0 = -1.09928e-7
+ wetab = 2.7482e-8
+ wkvth0we = 2e-12
+ trnqsmod = 0
+ cgidl = 0.22
+ rshg = 15.6
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ paigsd = -5.5708045e-23
+ permod = 1
+ pbswd = 0.8
+ pbsws = 0.8
+ )

.model nch_sf_21 nmos (
+ level = 54
+ acnqsmod = 0
+ dmcgt = 0
+ version = 4.5
+ tcjsw = 0.000357
+ ptvfbsdoff = 0
+ tempmod = 0
+ rbodymod = 0
+ tpbswg = 0.0009
+ aigbacc = 0.02
+ bigsd = 0.00125
+ wvoff = 1.0089489999999996e-10
+ ptvoff = 6.7086074e-18
+ wvsat = -0.0116031636
+ waigsd = 3.0872445e-12
+ aigbinv = 0.0163
+ wvth0 = 1.0690214590000001e-8
+ wpdiblc2 = 3.4958017e-9
+ waigc = 1.7847398e-12
+ diomod = 1
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 2.9779200000000003e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.9779200000000003e-10
+ lketa = -3.6124213e-8
+ xpart = 1
+ keta = 0.068466797
+ egidl = 0.29734
+ mjswgd = 0.85
+ mjswgs = 0.85
+ wkvth0we = 2e-12
+ poxedge = 1
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ tcjswg = 0.001
+ lcit = 6.9521194e-11
+ pvfbsdoff = 0
+ kt1l = 0
+ trnqsmod = 0
+ binunit = 2
+ lint = 9.7879675e-9
+ lkt1 = 4.7588252e-10
+ lkt2 = 9.4878496e-10
+ lmax = 2.1577e-7
+ lmin = 9e-8
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ rgatemod = 0
+ minv = -0.3
+ lua1 = 1.428412e-17
+ pvoff = 1.2597136100000002e-15
+ lub1 = -6.086010399999999e-26
+ luc1 = -3.3484914000000002e-18
+ tnjtsswg = 1
+ fprout = 300
+ ndep = 1e+18
+ cdscb = 0
+ cdscd = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ pvsat = 2.315286599999985e-11
+ lwlc = 0
+ wk2we = 5e-12
+ pvth0 = -2.10841744e-15
+ moin = 5.1
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ drout = 0.56
+ nigc = 3.083
+ paigc = 7.0313197e-18
+ wtvoff = -2.7645419e-10
+ voffl = 0
+ noff = 2.7195
+ weta0 = -1.09928e-7
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ wetab = 2.7482e-8
+ lpclm = 5.9671804e-8
+ capmod = 2
+ wku0we = 2e-11
+ ntox = 1.0
+ cgidl = 0.22
+ pcit = -2.1161006999999998e-17
+ pclm = 0.34708024
+ mobmod = 0
+ njtsswg = 9
+ phin = 0.15
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ pkt1 = -1.2810175000000001e-15
+ pkt2 = -1.739649e-15
+ pbswd = 0.8
+ pbsws = 0.8
+ a0 = 1.2892878
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 51380.779
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = -0.031682087000000005
+ k3 = -1.8419
+ em = 1000000.0
+ ckappad = 0.6
+ ckappas = 0.6
+ ll = -1.18e-13
+ lw = 0
+ u0 = 0.011619764000000001
+ w0 = 0
+ ua = -2.2703742e-9
+ ub = 2.053795462e-18
+ uc = 5.2246809e-11
+ ud = 0
+ pdiblc1 = 0
+ pdiblc2 = 0.010471563
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 3.4e-9
+ pdiblcb = -0.3
+ rbdb = 50
+ pua1 = -9.0422848e-24
+ prwb = 0
+ pdits = 0
+ laigsd = -6.8373623e-17
+ prwg = 0
+ pub1 = 1.3437735999999999e-32
+ puc1 = 2.6251991999999997e-24
+ cigsd = 0.069865
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ rdsw = 100
+ ijthsfwd = 0.01
+ bigbacc = 0.002588
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ kvth0we = 0.00018
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ tnoia = 0
+ ijthsrev = 0.01
+ lintnoi = -1.5e-8
+ bigbinv = 0.004953
+ peta0 = 0.0
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ rshg = 15.6
+ wketa = -5.2502872e-8
+ tpbsw = 0.0019
+ cjswd = 8.6592e-11
+ cjsws = 8.6592e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ ppdiblc2 = -3.8331042e-16
+ toxref = 3e-9
+ tnom = 25
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ scref = 1e-6
+ tvfbsdoff = 0.022
+ pigcd = 2.621
+ aigsd = 0.010772862
+ nfactor = 1
+ ltvoff = 9.6416574e-11
+ wags = -1.187467e-6
+ lvoff = -8.718213999999996e-10
+ pkvth0we = -1.3e-19
+ wcit = 1.2500316e-10
+ lvsat = -7.817471000000006e-5
+ lvth0 = -5.796310299999999e-9
+ voff = -0.16014500000000004
+ acde = 0.4
+ delta = 0.007595625
+ laigc = -1.4310771e-11
+ vfbsdoff = 0.02
+ vsat = 114971.1026
+ wint = 0
+ vth0 = 0.44879110699999997
+ rnoia = 0
+ rnoib = 0
+ lku0we = 2.5e-11
+ wkt1 = -7.3537768e-9
+ wkt2 = 1.0152376e-8
+ nigbacc = 10
+ wmax = 9.025999999999999e-7
+ epsrox = 3.9
+ aigc = 0.011560684
+ wmin = 5.426e-7
+ wvfbsdoff = 0
+ pketa = 1.139354e-14
+ lvfbsdoff = 0
+ ngate = 8e+20
+ rdsmod = 0
+ ngcon = 1
+ paramchk = 1
+ wpclm = 8.9560432e-7
+ igbmod = 1
+ wua1 = 5.7543559e-17
+ wub1 = -8.4794537e-26
+ wuc1 = -4.510386400000001e-17
+ gbmin = 1e-12
+ nigbinv = 10
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ bigc = 0.001442
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ wwlc = 0
+ pbswgd = 0.95
+ pbswgs = 0.95
+ cdsc = 0
+ igcmod = 1
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ ijthdfwd = 0.01
+ xtis = 3
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ fnoimod = 1
+ eigbinv = 1.1
+ ags = 5.2695
+ ijthdrev = 0.01
+ cjd = 0.001432992
+ cit = 0.0014357747
+ cjs = 0.001432992
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 1.30529375e-8
+ paigsd = 4.6587859e-23
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ tvoff = 0.00014539643
+ lpdiblc2 = -2.045371e-10
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ permod = 1
+ la0 = 6.8373618e-8
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = 0.0010900743
+ kt1 = -0.28113564
+ lk2 = -2.0436616e-10
+ kt2 = -0.099392124
+ llc = -1.18e-13
+ lln = 0.7
+ wtvfbsdoff = 0
+ lu0 = -2.3161917000000002e-10
+ mjd = 0.26
+ lua = 1.7344554e-17
+ mjs = 0.26
+ lub = -2.7790142600000004e-26
+ luc = -5.3126584e-18
+ lud = 0
+ k2we = 5e-5
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = -4.6587862e-14
+ nsd = 1e+20
+ dsub = 0.75
+ pbd = 0.52
+ pat = -1.7788972999999999e-9
+ pbs = 0.52
+ pk2 = -1.7344476e-15
+ cigbacc = 0.32875
+ dtox = 2.7e-10
+ ku0we = -0.0007
+ pu0 = 1.828211e-18
+ beta0 = 13
+ prt = 0
+ pua = 1.2335294e-23
+ pub = -1.88032504e-32
+ puc = -1.1996375e-24
+ pud = 0
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ leta0 = -1.6000000000000003e-9
+ ltvfbsdoff = 0
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 6.1325358e-10
+ ub1 = -3.2064524e-19
+ uc1 = 1.1057065000000001e-10
+ tnoimod = 0
+ tpb = 0.0014
+ ppclm = -6.7808634e-14
+ wa0 = -8.7848444e-7
+ voffcv = -0.16942
+ wpemod = 1
+ ute = -1
+ wat = 0.016319757
+ eta0 = 0.42133333
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 1.0517006e-8
+ lkvth0we = -2e-12
+ etab = -0.29033333
+ wlc = 0
+ wln = 1
+ wu0 = -6.079771099999999e-11
+ xgl = -1.09e-8
+ xgw = 0
+ dlcig = 2.5e-9
+ wua = -7.6059319e-17
+ wub = 9.256491399999999e-26
+ wuc = 4.1739756e-18
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ bgidl = 2320000000.0
+ cigbinv = 0.006
+ )

.model nch_sf_22 nmos (
+ level = 54
+ phin = 0.15
+ cjswd = 8.6592e-11
+ cjsws = 8.6592e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ pkt1 = -2.623551e-15
+ pkt2 = 8.0276583e-16
+ ptvoff = -9.1490879e-17
+ nfactor = 1
+ paramchk = 1
+ waigsd = 3.0879615e-12
+ diomod = 1
+ rbdb = 50
+ pua1 = -1.6477593e-25
+ prwb = 0
+ prwg = 0
+ pub1 = 1.4693022e-32
+ puc1 = 5.722749999999999e-24
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ pditsd = 0
+ pditsl = 0
+ rbsb = 50
+ pvag = 1.2
+ cjswgd = 2.9779200000000003e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.9779200000000003e-10
+ rdsw = 100
+ ijthdfwd = 0.01
+ scref = 1e-6
+ tvfbsdoff = 0.022
+ nigbacc = 10
+ pigcd = 2.621
+ aigsd = 0.010772861
+ mjswgd = 0.85
+ mjswgs = 0.85
+ lvoff = -4.808304999999992e-10
+ tcjswg = 0.001
+ lvsat = 0.0014054919840000002
+ ijthdrev = 0.01
+ lvth0 = 6.877404000000001e-10
+ nigbinv = 10
+ delta = 0.007595625
+ rshg = 15.6
+ laigc = -8.7106488e-12
+ lpdiblc2 = -4.1841324e-15
+ rnoia = 0
+ rnoib = 0
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ pketa = -2.7052976e-14
+ ngate = 8e+20
+ ngcon = 1
+ wpclm = 4.0103412e-7
+ fnoimod = 1
+ fprout = 300
+ eigbinv = 1.1
+ gbmin = 1e-12
+ tnom = 25
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ xrcrg1 = 12
+ xrcrg2 = 1
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ lkvth0we = -2e-12
+ wtvoff = 7.682212e-10
+ ags = 5.2695
+ cjd = 0.001432992
+ cit = 0.00076911293
+ cjs = 0.001432992
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ acnqsmod = 0
+ dlc = 3.26497e-9
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ wags = -1.187467e-6
+ capmod = 2
+ wcit = -3.1211371e-10
+ cigbacc = 0.32875
+ rbodymod = 0
+ wku0we = 2e-11
+ la0 = -1.9182963e-7
+ voff = -0.164304478
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.00161425008
+ acde = 0.4
+ kt1 = -0.33033037
+ lk2 = -1.3785596e-9
+ kt2 = -0.066210327
+ mobmod = 0
+ llc = 0
+ lln = 1
+ lu0 = -7.115591899999999e-11
+ tnoimod = 0
+ mjd = 0.26
+ tvoff = 0.00053139469
+ lua = 2.7860169e-17
+ mjs = 0.26
+ lub = -2.7395085e-26
+ luc = 1.41139916e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ vsat = 99187.40900000001
+ njs = 1.02
+ pa0 = 2.0809981e-13
+ wint = 0
+ vth0 = 0.379811848
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 2.0933444199999996e-9
+ pbs = 0.52
+ pk2 = 9.5324632e-16
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ wkt1 = 6.9284939e-9
+ wkt2 = -1.689459e-8
+ pu0 = -3.7471417e-18
+ wmax = 9.025999999999999e-7
+ prt = 0
+ pua = -6.3654423e-24
+ pub = 7.034010899999999e-33
+ puc = -7.127418999999999e-24
+ pud = 0
+ cigbinv = 0.006
+ aigc = 0.011501109
+ wmin = 5.426e-7
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 8.1588744e-10
+ ub1 = -6.9089562e-19
+ uc1 = 1.1957352299999998e-10
+ tpb = 0.0014
+ wa0 = -3.5879278e-6
+ ute = -1
+ wat = -0.024874303599999998
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -1.8075483e-8
+ ku0we = -0.0007
+ wlc = 0
+ wln = 1
+ wu0 = -1.4854479999999955e-12
+ xgl = -1.09e-8
+ xgw = 0
+ beta0 = 13
+ wua = 1.2288469e-16
+ wub = -1.8229956900000002e-25
+ wua1 = -3.6898024e-17
+ wuc = 6.7235478e-17
+ wud = 0
+ wub1 = -9.8148649e-26
+ wuc1 = -7.8056508e-17
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ leta0 = -1.2426782e-8
+ wpdiblc2 = -5.8202891e-10
+ letab = -2.2164189e-8
+ version = 4.5
+ bigc = 0.001442
+ laigsd = 3.8113519e-17
+ tempmod = 0
+ wwlc = 0
+ ppclm = -2.1319035e-14
+ dlcig = 2.5e-9
+ cdsc = 0
+ bgidl = 2320000000.0
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ aigbacc = 0.02
+ xtis = 3
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ dmcgt = 0
+ tcjsw = 0.000357
+ wkvth0we = 2e-12
+ aigbinv = 0.0163
+ a0 = 4.0574074
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 80150.18699999999
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = -0.019190666999999998
+ k3 = -1.8419
+ em = 1000000.0
+ ll = 0
+ lw = 0
+ trnqsmod = 0
+ u0 = 0.009912708000000001
+ w0 = 0
+ ua = -2.3822425e-9
+ ub = 2.049592666e-18
+ uc = -1.5441968e-10
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 3.4e-9
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ bigsd = 0.00125
+ wvoff = 3.0122529e-8
+ k2we = 5e-5
+ dsub = 0.75
+ dtox = 2.7e-10
+ wvsat = -0.019673989999999995
+ toxref = 3e-9
+ wvth0 = -3.2932843000000014e-8
+ rgatemod = 0
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ tnjtsswg = 1
+ poxedge = 1
+ waigc = 1.9067031e-10
+ eta0 = 0.53651186
+ etab = -0.054544089
+ binunit = 2
+ lketa = 6.7720908e-8
+ xpart = 1
+ ltvoff = 6.0132739e-11
+ egidl = 0.29734
+ pvfbsdoff = 0
+ lku0we = 2.5e-11
+ epsrox = 3.9
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ rdsmod = 0
+ igbmod = 1
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ pvoff = -1.5623199999999997e-15
+ pbswgd = 0.95
+ pbswgs = 0.95
+ cdscb = 0
+ cdscd = 0
+ pvsat = 7.818105999999996e-10
+ wk2we = 5e-12
+ igcmod = 1
+ pvth0 = 1.99215e-15
+ drout = 0.56
+ paigc = -1.0723924e-17
+ ijthsfwd = 0.01
+ njtsswg = 9
+ voffl = 0
+ keta = -1.0362685
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ weta0 = -2.7932191e-7
+ wetab = 6.5877739e-8
+ wtvfbsdoff = 0
+ lpclm = -1.3225653e-8
+ ckappad = 0.6
+ ckappas = 0.6
+ jswd = 1.28e-13
+ pdiblc1 = 0
+ jsws = 1.28e-13
+ pdiblc2 = 0.0082956805
+ lcit = 1.3218741e-10
+ paigsd = -2.0809977e-23
+ pdiblcb = -0.3
+ ijthsrev = 0.01
+ kt1l = 0
+ cgidl = 0.22
+ ltvfbsdoff = 0
+ permod = 1
+ lint = 0
+ lkt1 = 5.1001869e-9
+ lkt2 = -2.1703039e-9
+ lmax = 9e-8
+ lmin = 5.4e-8
+ pbswd = 0.8
+ pbsws = 0.8
+ bigbacc = 0.002588
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ ppdiblc2 = 5.6582339e-21
+ minv = -0.3
+ kvth0we = 0.00018
+ lua1 = -4.7634626e-18
+ lub1 = -2.6056569000000004e-26
+ luc1 = -4.194757189999999e-18
+ voffcv = -0.16942
+ wpemod = 1
+ pdits = 0
+ ndep = 1e+18
+ lintnoi = -1.5e-8
+ cigsd = 0.069865
+ ptvfbsdoff = 0
+ lwlc = 0
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ moin = 5.1
+ vtsswgs = 4.2
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ nigc = 3.083
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ pkvth0we = -1.3e-19
+ tnoia = 0
+ tpbswg = 0.0009
+ peta0 = 1.5923028e-14
+ ntox = 1.0
+ pcit = 1.99279785e-17
+ petab = -3.6091995e-15
+ pclm = 1.1225851
+ vfbsdoff = 0.02
+ wketa = 3.5650261e-7
+ tpbsw = 0.0019
+ )

.model nch_sf_23 nmos (
+ level = 54
+ pditsl = 0
+ cjswgd = 2.9779200000000003e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.9779200000000003e-10
+ cdsc = 0
+ lketa = -2.0578185e-8
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ ijthsfwd = 0.01
+ xtid = 3
+ xtis = 3
+ xpart = 1
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ mjswgd = 0.85
+ mjswgs = 0.85
+ egidl = 0.29734
+ tcjswg = 0.001
+ pvfbsdoff = 0
+ ijthsrev = 0.01
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ njtsswg = 9
+ k2we = 5e-5
+ dsub = 0.75
+ dtox = 2.7e-10
+ fprout = 300
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ xrcrg1 = 12
+ xrcrg2 = 1
+ pvoff = -3.96509854e-15
+ ckappad = 0.6
+ ckappas = 0.6
+ cdscb = 0
+ pdiblc1 = 0
+ pdiblc2 = 0.0082956083
+ cdscd = 0
+ pdiblcb = -0.3
+ pvsat = 3.6118091109999995e-9
+ eta0 = 0.49180426
+ etab = -1.1686036
+ wk2we = 5e-12
+ pvth0 = 4.8634049e-15
+ drout = 0.56
+ wtvoff = -4.625476e-9
+ paigc = -1.7630641e-18
+ voffl = 0
+ weta0 = 1.6706711e-7
+ capmod = 2
+ bigbacc = 0.002588
+ wetab = -6.7375536e-8
+ pkvth0we = -1.3e-19
+ lpclm = -4.9784452e-8
+ wku0we = 2e-11
+ mobmod = 0
+ kvth0we = 0.00018
+ cgidl = 0.22
+ vfbsdoff = 0.02
+ lintnoi = -1.5e-8
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ pbswd = 0.8
+ pbsws = 0.8
+ paramchk = 1
+ laigsd = -3.1577826e-17
+ pdits = 0
+ cigsd = 0.069865
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ ijthdfwd = 0.01
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ keta = 0.48612964
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ nfactor = 1
+ tnoia = 0
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ ijthdrev = 0.01
+ lcit = 3.9401345000000003e-10
+ peta0 = -9.9675358e-15
+ kt1l = 0
+ petab = 4.1194905e-15
+ wketa = -1.8474011e-7
+ tpbsw = 0.0019
+ lint = 0
+ cjswd = 8.6592e-11
+ cjsws = 8.6592e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ lkt1 = -1.5114128e-8
+ lkt2 = -1.4213753e-9
+ lmax = 5.4e-8
+ lmin = 4.5e-8
+ nigbacc = 10
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ toxref = 3e-9
+ minv = -0.3
+ lua1 = 7.7308837e-17
+ lub1 = -1.5651426199999998e-25
+ luc1 = -7.947051999999997e-18
+ ndep = 1e+18
+ lkvth0we = -2e-12
+ nigbinv = 10
+ lwlc = 0
+ moin = 5.1
+ a0 = 11.080765
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 31524.241299999994
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ tvfbsdoff = 0.022
+ k2 = 0.014747898
+ k3 = -1.8419
+ em = 1000000.0
+ ll = 0
+ lw = 0
+ u0 = -0.00036107273999999996
+ scref = 1e-6
+ nigc = 3.083
+ w0 = 0
+ ua = -5.2066121e-9
+ ub = 5.20056154e-18
+ uc = 2.7090556e-10
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 3.4e-9
+ pigcd = 2.621
+ aigsd = 0.010772862
+ ltvoff = -1.4697355e-10
+ acnqsmod = 0
+ lvoff = 1.6278058999999974e-9
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ fnoimod = 1
+ lvsat = -0.00504394337
+ rbodymod = 0
+ lvth0 = -3.1936672999999985e-9
+ eigbinv = 1.1
+ ntox = 1.0
+ delta = 0.007595625
+ pcit = 3.4096077e-17
+ lku0we = 2.5e-11
+ pclm = 1.7529092
+ laigc = -1.8175152e-11
+ epsrox = 3.9
+ rnoia = 0
+ rnoib = 0
+ wvfbsdoff = 0
+ phin = 0.15
+ lvfbsdoff = 0
+ rdsmod = 0
+ pketa = 4.339103e-15
+ igbmod = 1
+ ngate = 8e+20
+ pkt1 = 1.1764455e-14
+ pkt2 = 3.1759909e-15
+ ngcon = 1
+ wpclm = -7.2697212e-7
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ wpdiblc2 = -5.8193135e-10
+ pbswgd = 0.95
+ gbmin = 1e-12
+ pbswgs = 0.95
+ cigbacc = 0.32875
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ ags = 5.2695
+ rbdb = 50
+ pua1 = -6.2039198e-23
+ prwb = 0
+ prwg = 0
+ pub1 = 1.08600889e-31
+ puc1 = 4.339185599999997e-24
+ igcmod = 1
+ wtvfbsdoff = 0
+ cjd = 0.001432992
+ cit = -0.0037451293
+ cjs = 0.001432992
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ dlc = 3.26497e-9
+ k3b = 1.9326
+ tnoimod = 0
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ rdsw = 100
+ ltvfbsdoff = 0
+ cigbinv = 0.006
+ la0 = -5.9918439e-7
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = 0.0012060548200000004
+ kt1 = 0.018192305
+ lk2 = -3.3469964e-9
+ kt2 = -0.079122889
+ llc = 0
+ lln = 1
+ lu0 = 5.2472336e-10
+ mjd = 0.26
+ lua = 1.9167361e-16
+ mjs = 0.26
+ lub = -2.101512744e-25
+ luc = -1.0554871600000002e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 1.4611928e-13
+ wkvth0we = 2e-12
+ nsd = 1e+20
+ pbd = 0.52
+ pat = -1.4311335800000002e-9
+ pbs = 0.52
+ pk2 = 2.1253177e-15
+ paigsd = 1.0451534e-29
+ pu0 = -5.8805924e-17
+ prt = 0
+ pua = -7.1470289e-23
+ pub = 9.665873609999999e-32
+ puc = 4.556057900000002e-24
+ pud = 0
+ version = 4.5
+ rsh = 17.5
+ trnqsmod = 0
+ tcj = 0.00076
+ ua1 = -5.9915221e-10
+ ub1 = 1.5583749700000001e-18
+ uc1 = 1.8426858999999987e-10
+ rshg = 15.6
+ tempmod = 0
+ tvoff = 0.0041021928
+ tpb = 0.0014
+ wa0 = -2.5192978e-6
+ permod = 1
+ ute = -1
+ wat = 0.035892558
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -3.8283609e-8
+ xjbvd = 1
+ xjbvs = 1
+ wlc = 0
+ wln = 1
+ lk2we = -1.5e-12
+ wu0 = 9.478039e-10
+ xgl = -1.09e-8
+ xgw = 0
+ wua = 1.2453821e-15
+ wub = -1.72755342e-24
+ wuc = -1.3420376999999993e-16
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ ptvfbsdoff = 0
+ aigbacc = 0.02
+ ku0we = -0.0007
+ beta0 = 13
+ rgatemod = 0
+ leta0 = -9.833740899999999e-9
+ letab = 4.245126e-8
+ voffcv = -0.16942
+ wpemod = 1
+ tnom = 25
+ tnjtsswg = 1
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ aigbinv = 0.0163
+ ppclm = 4.4105328e-14
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ wags = -1.187467e-6
+ dmcgt = 0
+ tcjsw = 0.000357
+ wcit = -5.5639126e-10
+ tpbswg = 0.0009
+ voff = -0.20066027000000003
+ acde = 0.4
+ poxedge = 1
+ vsat = 210384.59399999995
+ wint = 0
+ vth0 = 0.44673267
+ bigsd = 0.00125
+ binunit = 2
+ wkt1 = -2.4114058e-7
+ wkt2 = -5.7812263e-8
+ wmax = 9.025999999999999e-7
+ aigc = 0.01166429
+ wmin = 5.426e-7
+ ptvoff = 2.2134356e-16
+ wvoff = 7.154973409999999e-8
+ waigsd = 3.0876027e-12
+ wvsat = -0.06846706247
+ wua1 = 1.0299024e-15
+ wub1 = -1.71724981e-24
+ wuc1 = -5.4200488999999977e-17
+ wvth0 = -8.243723199999998e-8
+ diomod = 1
+ bigc = 0.001442
+ waigc = 3.6172725e-11
+ wwlc = 0
+ pditsd = 0
+ )

.model nch_sf_24 nmos (
+ level = 54
+ lvsat = -0.0034499051999999993
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lvth0 = 2.938582699999999e-9
+ lcit = 2.9117288e-10
+ trnqsmod = 0
+ kt1l = 0
+ cigbacc = 0.32875
+ delta = 0.007595625
+ laigc = -7.4258513e-12
+ rnoia = 0
+ rnoib = 0
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ tnoimod = 0
+ lint = 0
+ lkt1 = 7.714149e-10
+ lkt2 = 6.4873536e-9
+ lmax = 4.5e-8
+ pketa = 3.05233408e-14
+ ags = 5.2695
+ ngate = 8e+20
+ lmin = 3.6e-8
+ cigbinv = 0.006
+ ngcon = 1
+ lpe0 = 9.2e-8
+ cjd = 0.001432992
+ cit = -0.001646336
+ fprout = 300
+ cjs = 0.001432992
+ clc = 1e-7
+ wpclm = 9.524622100000001e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ lpeb = 2.5e-7
+ dlc = 3.26497e-9
+ k3b = 1.9326
+ xrcrg1 = 12
+ xrcrg2 = 1
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ rgatemod = 0
+ gbmin = 1e-12
+ minv = -0.3
+ tnjtsswg = 1
+ lua1 = -6.7547343e-17
+ lub1 = 1.3220925399999999e-25
+ luc1 = 3.2044560000000004e-17
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ ndep = 1e+18
+ la0 = -5.581062559999999e-7
+ version = 4.5
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.00159504779
+ wtvoff = -5.6534448e-10
+ lwlc = 0
+ kt1 = -0.30600245
+ lk2 = -3.4047834e-9
+ kt2 = -0.24052552
+ llc = 0
+ moin = 5.1
+ lln = 1
+ lu0 = 6.9334295e-10
+ tempmod = 0
+ mjd = 0.26
+ lua = 1.9963428e-16
+ mjs = 0.26
+ lub = -1.86515944e-25
+ luc = -1.3855022100000003e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 1.41312605e-13
+ nigc = 3.083
+ nsd = 1e+20
+ pbd = 0.52
+ pat = -1.5570081000000008e-10
+ pbs = 0.52
+ pk2 = 1.540171e-16
+ pu0 = -4.3529201000000005e-16
+ prt = 0
+ pua = -1.24177601e-22
+ pub = 1.2166737845000001e-31
+ puc = -3.231882900000001e-24
+ pud = 0
+ aigbacc = 0.02
+ capmod = 2
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 2.3570964e-9
+ ub1 = -4.3339417e-18
+ uc1 = -6.318859999999999e-10
+ tpb = 0.0014
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ wku0we = 2e-11
+ wa0 = -2.4212027299999997e-6
+ ute = -1
+ wat = 0.009863318999999999
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 1.947015e-9
+ wlc = 0
+ wln = 1
+ wu0 = 8.6311905e-9
+ xgl = -1.09e-8
+ mobmod = 0
+ xgw = 0
+ wua = 2.32104147e-15
+ wub = -2.2379339299999998e-24
+ wuc = 2.4733810000000014e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ ntox = 1.0
+ pcit = -5.917525700000001e-17
+ pclm = 0.021884800000000038
+ tvoff = 0.0045807103
+ aigbinv = 0.0163
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ phin = 0.15
+ pkt1 = -5.4745624e-15
+ pkt2 = -2.9889728e-15
+ ku0we = -0.0007
+ beta0 = 13
+ laigsd = 2.1777751e-17
+ leta0 = 4.423777099999998e-9
+ letab = 3.2196399e-8
+ ppclm = -3.8186956000000005e-14
+ rbdb = 50
+ pua1 = 5.0551945e-23
+ prwb = 0
+ prwg = 0
+ pub1 = -9.5529116e-32
+ puc1 = -2.5642617899999998e-23
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ poxedge = 1
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ rdsw = 100
+ ijthsfwd = 0.01
+ binunit = 2
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ dmcgt = 0
+ tcjsw = 0.000357
+ ijthsrev = 0.01
+ rshg = 15.6
+ bigsd = 0.00125
+ wvoff = -4.4038220999999975e-8
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ toxref = 3e-9
+ wvsat = -0.03971696100000001
+ wvth0 = 1.8939272999999993e-8
+ tnom = 25
+ waigc = -1.3685053e-10
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ lketa = -4.89346675e-8
+ xpart = 1
+ ltvoff = -1.7042091e-10
+ egidl = 0.29734
+ njtsswg = 9
+ wags = -1.187467e-6
+ pkvth0we = -1.3e-19
+ pvfbsdoff = 0
+ wcit = 1.3471085999999997e-9
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ voff = 0.016693055000000012
+ lku0we = 2.5e-11
+ acde = 0.4
+ ckappad = 0.6
+ epsrox = 3.9
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.0082956083
+ vfbsdoff = 0.02
+ pdiblcb = -0.3
+ vsat = 177853.19600000003
+ wint = 0
+ vth0 = 0.32158466499999994
+ wkt1 = 1.1067611e-7
+ wkt2 = 6.8003321e-8
+ rdsmod = 0
+ wtvfbsdoff = 0
+ wmax = 9.025999999999999e-7
+ aigc = 0.011444916
+ wmin = 5.426e-7
+ igbmod = 1
+ a0 = 10.24243689
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 88689.602
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.015927223
+ k3 = -1.8419
+ em = 1000000.0
+ ll = 0
+ lw = 0
+ u0 = -0.0038022958
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ paramchk = 1
+ w0 = 0
+ ua = -5.369074800000001e-9
+ ub = 4.718207719999999e-18
+ uc = 3.3825556e-10
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 3.4e-9
+ ltvfbsdoff = 0
+ pbswgd = 0.95
+ pbswgs = 0.95
+ wua1 = -1.2678761e-15
+ wub1 = 2.44866871e-24
+ wuc1 = 5.576703800000001e-16
+ bigbacc = 0.002588
+ pvoff = 1.6987133300000001e-15
+ bigc = 0.001442
+ igcmod = 1
+ wwlc = 0
+ cdscb = 0
+ cdscd = 0
+ kvth0we = 0.00018
+ pvsat = 2.20305333e-9
+ wk2we = 5e-12
+ pvth0 = -1.0404569999999977e-16
+ drout = 0.56
+ cdsc = 0
+ lintnoi = -1.5e-8
+ paigc = 6.7150752e-18
+ cgbo = 0
+ ijthdfwd = 0.01
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ voffl = 0
+ cigc = 0.000625
+ ptvfbsdoff = 0
+ weta0 = -1.6294544599999998e-7
+ wetab = 1.0177792e-7
+ paigsd = 4.9710031e-30
+ lpclm = 3.5035747999999996e-8
+ ijthdrev = 0.01
+ cgidl = 0.22
+ permod = 1
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ pbswd = 0.8
+ pbsws = 0.8
+ k2we = 5e-5
+ dsub = 0.75
+ dtox = 2.7e-10
+ voffcv = -0.16942
+ wpemod = 1
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ nfactor = 1
+ pdits = 0
+ cigsd = 0.069865
+ eta0 = 0.20083450200000003
+ lkvth0we = -2e-12
+ etab = -0.95932067
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ acnqsmod = 0
+ nigbacc = 10
+ tpbswg = 0.0009
+ tnoia = 0
+ rbodymod = 0
+ peta0 = 6.20307972e-15
+ petab = -4.1690291e-15
+ wketa = -7.1911233e-7
+ tpbsw = 0.0019
+ nigbinv = 10
+ cjswd = 8.6592e-11
+ cjsws = 8.6592e-11
+ ptvoff = 2.2397114e-17
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ waigsd = 3.0876027e-12
+ diomod = 1
+ wpdiblc2 = -5.8193135e-10
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 2.9779200000000003e-10
+ pku0we = -1.5e-18
+ fnoimod = 1
+ cjswgs = 2.9779200000000003e-10
+ eigbinv = 1.1
+ tvfbsdoff = 0.022
+ scref = 1e-6
+ pigcd = 2.621
+ mjswgd = 0.85
+ aigsd = 0.010772861
+ mjswgs = 0.85
+ keta = 1.06483334
+ tcjswg = 0.001
+ lvoff = -9.022509e-9
+ wkvth0we = 2e-12
+ )

.model nch_sf_25 nmos (
+ level = 54
+ fprout = 300
+ xrcrg1 = 12
+ xrcrg2 = 1
+ pvoff = -4e-17
+ tnom = 25
+ cdscb = 0
+ cdscd = 0
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ wtvoff = 0
+ pvsat = 1.44e-11
+ lkvth0we = -2e-12
+ wk2we = 5e-12
+ pvth0 = 1.2e-16
+ drout = 0.56
+ voffl = 0
+ capmod = 2
+ acnqsmod = 0
+ wku0we = 2e-11
+ weta0 = -1.1162667e-8
+ wags = -5.746904e-8
+ wetab = 2.2325333e-8
+ mobmod = 0
+ wcit = 2.563688e-10
+ rbodymod = 0
+ nfactor = 1
+ voff = -0.13478422
+ acde = 0.4
+ cgidl = 0.22
+ vsat = 102889.02
+ wint = 0
+ vth0 = 0.39140512
+ wkt1 = 2.4629406130000002e-9
+ wkt2 = -5.3296152e-9
+ wmax = 5.426e-7
+ aigc = 0.011779434
+ wmin = 2.726e-7
+ pbswd = 0.8
+ pbsws = 0.8
+ wua1 = -1.874362e-16
+ nigbacc = 10
+ wub1 = 1.1464267e-25
+ wuc1 = -2.7527136e-17
+ wpdiblc2 = 4.9914968e-9
+ bigc = 0.001442
+ pdits = 0
+ wwlc = 0
+ cigsd = 0.069865
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ nigbinv = 10
+ xtis = 3
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ wkvth0we = 2e-12
+ tnoia = 0
+ trnqsmod = 0
+ peta0 = 0.0
+ fnoimod = 1
+ wketa = 1.6322115e-8
+ eigbinv = 1.1
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ tpbsw = 0.0019
+ dmdg = 0
+ cjswd = 8.6592e-11
+ cjsws = 8.6592e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ toxref = 3e-9
+ k2we = 5e-5
+ dsub = 0.75
+ dtox = 2.7e-10
+ rgatemod = 0
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ tnjtsswg = 1
+ tvfbsdoff = 0.022
+ eta0 = 0.24044444
+ etab = -0.28088889
+ cigbacc = 0.32875
+ ltvoff = 0
+ scref = 1e-6
+ pigcd = 2.621
+ tnoimod = 0
+ aigsd = 0.010772818
+ wtvfbsdoff = 0
+ lvoff = 1.6e-11
+ cigbinv = 0.006
+ lvsat = 0.00016
+ lku0we = 2.5e-11
+ lvth0 = 4.0000000000000007e-10
+ ltvfbsdoff = 0
+ epsrox = 3.9
+ delta = 0.007595625
+ ags = 1.06760667
+ wvfbsdoff = 0
+ cjd = 0.001432992
+ cit = 0.000342575
+ version = 4.5
+ cjs = 0.001432992
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ lvfbsdoff = 0
+ rnoia = 0
+ rnoib = 0
+ rdsmod = 0
+ dlc = 9.8024918e-9
+ k3b = 1.9326
+ tempmod = 0
+ igbmod = 1
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ ngate = 8e+20
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ ngcon = 1
+ la0 = 0
+ wpclm = 9.3989653e-8
+ pbswgd = 0.95
+ jsd = 6.11e-7
+ pbswgs = 0.95
+ jss = 6.11e-7
+ lat = 8e-5
+ aigbacc = 0.02
+ kt1 = -0.22055704
+ kt2 = -0.0354368
+ llc = 0
+ lln = 1
+ lu0 = -4e-12
+ mjd = 0.26
+ mjs = 0.26
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ gbmin = 1e-12
+ njs = 1.02
+ pa0 = 0
+ igcmod = 1
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 1.44e-11
+ jswgd = 1.28e-13
+ ptvfbsdoff = 0
+ pbs = 0.52
+ jswgs = 1.28e-13
+ pu0 = -1.2e-18
+ prt = 0
+ pud = 0
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 1.6212811e-9
+ ub1 = -8.7849211e-19
+ uc1 = 6.9356e-11
+ tpb = 0.0014
+ aigbinv = 0.0163
+ wa0 = -1.17208e-8
+ ijthsfwd = 0.01
+ ute = -1
+ wat = 0.071441067
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 1.8596306e-9
+ wlc = 0
+ wln = 1
+ wu0 = -1.2477067e-9
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -1.3097991e-16
+ wub = 9.54408e-26
+ wuc = -2.4557867e-18
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ keta = -0.084351302
+ a0 = 3.5424667
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = -58844.444
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.021767646
+ k3 = -1.8419
+ em = 1000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.017991111
+ jswd = 1.28e-13
+ w0 = 0
+ jsws = 1.28e-13
+ ijthsrev = 0.01
+ ua = -1.6762565e-9
+ ub = 2.0222e-18
+ uc = 6.1497778e-11
+ ud = 0
+ lcit = 8e-12
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 3.4e-9
+ permod = 1
+ kt1l = 0
+ tvoff = 0.0017628809
+ xjbvd = 1
+ xjbvs = 1
+ poxedge = 1
+ lk2we = -1.5e-12
+ lint = 6.5375218e-9
+ lkt1 = -2.4e-10
+ lmax = 2.001e-5
+ binunit = 2
+ lmin = 8.9991e-6
+ lpe0 = 9.2e-8
+ voffcv = -0.16942
+ wpemod = 1
+ lpeb = 2.5e-7
+ ku0we = -0.0007
+ beta0 = 13
+ leta0 = -1.6000000000000003e-9
+ minv = -0.3
+ lub1 = 2.4000000000000004e-27
+ ndep = 1e+18
+ lwlc = 0
+ dlcig = 2.5e-9
+ moin = 5.1
+ bgidl = 2320000000.0
+ nigc = 3.083
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ noff = 2.7195
+ dmcgt = 0
+ noia = 3.11e+42
+ noib = 1.22e+22
+ pkvth0we = -1.3e-19
+ noic = 45200000.0
+ tpbswg = 0.0009
+ tcjsw = 0.000357
+ ntox = 1.0
+ pcit = 1.2000000000000001e-17
+ pclm = 1.5094578
+ vfbsdoff = 0.02
+ bigsd = 0.00125
+ ptvoff = 0
+ phin = 0.15
+ waigsd = 3.1112026e-12
+ wvoff = 1.3365577e-8
+ pkt1 = -1.76e-16
+ paramchk = 1
+ diomod = 1
+ wvsat = -0.0028059037
+ wvth0 = -1.5368414000000002e-8
+ njtsswg = 9
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 2.9779200000000003e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.9779200000000003e-10
+ waigc = 2.8724444e-11
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ rbdb = 50
+ prwb = 0
+ prwg = 0
+ pub1 = 1.6e-34
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.0047029422
+ rdsw = 100
+ pdiblcb = -0.3
+ ijthdfwd = 0.01
+ mjswgd = 0.85
+ xpart = 1
+ mjswgs = 0.85
+ tcjswg = 0.001
+ egidl = 0.29734
+ pvfbsdoff = 0
+ bigbacc = 0.002588
+ ijthdrev = 0.01
+ rshg = 15.6
+ kvth0we = 0.00018
+ lintnoi = -1.5e-8
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ )

.model nch_sf_26 nmos (
+ level = 54
+ poxedge = 1
+ capmod = 2
+ wku0we = 2e-11
+ binunit = 2
+ mobmod = 0
+ pkvth0we = -1.3e-19
+ tvoff = 0.0019388906
+ vfbsdoff = 0.02
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ laigsd = -2.019482e-16
+ paramchk = 1
+ ku0we = -0.0007
+ beta0 = 13
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ leta0 = -1.6000000000000003e-9
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ ijthdfwd = 0.01
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ keta = -0.091670067
+ dmcgt = 0
+ tcjsw = 0.000357
+ lags = -1.7808411e-7
+ njtsswg = 9
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ ijthdrev = 0.01
+ lcit = 6.7578289e-10
+ kt1l = 0
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ lpdiblc2 = 2.6261368e-8
+ bigsd = 0.00125
+ ckappad = 0.6
+ ckappas = 0.6
+ lint = 6.5375218e-9
+ pdiblc1 = 0
+ pdiblc2 = 0.0017817666
+ toxref = 3e-9
+ pdiblcb = -0.3
+ lkt1 = 8.817275899999999e-9
+ lkt2 = -2.1662043e-8
+ lmax = 8.9991e-6
+ wvoff = 1.3633649999999999e-8
+ lmin = 8.9908e-7
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ wvsat = -0.0028059037
+ wvth0 = -1.5716317e-8
+ minv = -0.3
+ wtvfbsdoff = 0
+ lua1 = -8.9279603e-16
+ lub1 = 6.8784226e-25
+ luc1 = -5.9256432e-18
+ waigc = 2.989874e-11
+ bigbacc = 0.002588
+ ndep = 1e+18
+ lkvth0we = -2e-12
+ lwlc = 0
+ moin = 5.1
+ ltvoff = -1.582327e-9
+ ltvfbsdoff = 0
+ lketa = 6.5795695e-8
+ kvth0we = 0.00018
+ nigc = 3.083
+ xpart = 1
+ lintnoi = -1.5e-8
+ acnqsmod = 0
+ pvfbsdoff = 0
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ egidl = 0.29734
+ vtsswgs = 4.2
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ lku0we = 2.5e-11
+ rbodymod = 0
+ epsrox = 3.9
+ pags = 1.7531187e-13
+ ntox = 1.0
+ pcit = -9.498337e-17
+ pclm = 1.5094578
+ rdsmod = 0
+ ptvfbsdoff = 0
+ igbmod = 1
+ phin = 0.15
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ pbswgd = 0.95
+ pkt1 = -2.7553875e-14
+ pkt2 = -4.4253241e-16
+ pbswgs = 0.95
+ igcmod = 1
+ wpdiblc2 = 5.7318301e-9
+ pvoff = -2.4499792999999998e-15
+ cdscb = 0
+ cdscd = 0
+ rbdb = 50
+ pua1 = 1.9942546e-22
+ prwb = 0
+ prwg = 0
+ pub1 = -1.9923615000000002e-31
+ puc1 = 1.7835157e-23
+ nfactor = 1
+ pvsat = 1.44e-11
+ rbpb = 50
+ rbpd = 50
+ wk2we = 5e-12
+ rbps = 50
+ pvth0 = 3.2476501999999998e-15
+ rbsb = 50
+ pvag = 1.2
+ drout = 0.56
+ rdsw = 100
+ paigc = -1.0556924e-17
+ voffl = 0
+ paigsd = 1.1026372e-22
+ weta0 = -1.1162667e-8
+ wetab = 2.2325333e-8
+ wkvth0we = 2e-12
+ nigbacc = 10
+ permod = 1
+ trnqsmod = 0
+ cgidl = 0.22
+ rshg = 15.6
+ nigbinv = 10
+ pbswd = 0.8
+ pbsws = 0.8
+ voffcv = -0.16942
+ wpemod = 1
+ rgatemod = 0
+ tnjtsswg = 1
+ tnom = 25
+ pdits = 0
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ a0 = 3.8452644
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ cigsd = 0.069865
+ b1 = 0
+ at = -81312.781
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.023323392000000002
+ k3 = -1.8419
+ em = 1000000.0
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ ll = 0
+ lw = 0
+ u0 = 0.01824456
+ w0 = 0
+ fnoimod = 1
+ ua = -1.6436128e-9
+ ub = 2.0158412e-18
+ uc = 5.8736458e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 3.4e-9
+ eigbinv = 1.1
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ tpbswg = 0.0009
+ wags = -7.6969804e-8
+ wcit = 2.6826906e-10
+ tnoia = 0
+ voff = -0.13348839
+ peta0 = 0.0
+ acde = 0.4
+ wketa = 1.8850903e-8
+ vsat = 102889.02
+ ptvoff = 2.7553621e-16
+ wint = 0
+ tpbsw = 0.0019
+ vth0 = 0.38569778
+ cigbacc = 0.32875
+ waigsd = 3.1111904e-12
+ wkt1 = 5.5083105e-9
+ wkt2 = -5.2803902e-9
+ cjswd = 8.6592e-11
+ cjsws = 8.6592e-11
+ wmax = 5.426e-7
+ mjswd = 0.11
+ aigc = 0.011795195
+ mjsws = 0.11
+ wmin = 2.726e-7
+ agidl = 9.41e-8
+ diomod = 1
+ tnoimod = 0
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 2.9779200000000003e-10
+ pku0we = -1.5e-18
+ wua1 = -2.0961923e-16
+ wub1 = 1.3682244e-25
+ cjswgs = 2.9779200000000003e-10
+ wuc1 = -2.9511024e-17
+ cigbinv = 0.006
+ bigc = 0.001442
+ wwlc = 0
+ tvfbsdoff = 0.022
+ cdsc = 0
+ mjswgd = 0.85
+ mjswgs = 0.85
+ scref = 1e-6
+ version = 4.5
+ ijthsfwd = 0.01
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ pigcd = 2.621
+ cgsl = 3.31989e-12
+ tcjswg = 0.001
+ cgso = 4.90562e-11
+ tempmod = 0
+ aigsd = 0.010772818
+ cigc = 0.000625
+ ags = 1.0874158
+ lvoff = -1.1633525e-8
+ cjd = 0.001432992
+ cit = 0.00026829437
+ cjs = 0.001432992
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ aigbacc = 0.02
+ dlc = 9.8024918e-9
+ lvsat = 0.00016
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ lvth0 = 5.1708999e-8
+ ijthsrev = 0.01
+ delta = 0.007595625
+ laigc = -1.416882e-10
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ la0 = -2.722152e-6
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ rnoia = 0
+ rnoib = 0
+ dmdg = 0
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = 0.20207035
+ kt1 = -0.22156452
+ lk2 = -1.3986155e-8
+ kt2 = -0.033027229
+ llc = 0
+ lln = 1
+ lu0 = -2.2825026e-9
+ mjd = 0.26
+ aigbinv = 0.0163
+ lua = -2.9346741e-16
+ mjs = 0.26
+ lub = 5.7165214e-26
+ luc = 2.4824263e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 3.4236885e-13
+ fprout = 300
+ nsd = 1e+20
+ pbd = 0.52
+ pat = -6.367392400000001e-8
+ pbs = 0.52
+ pketa = -2.2733801e-14
+ pk2 = -1.3939214e-15
+ ngate = 8e+20
+ pu0 = 1.6419558e-16
+ xrcrg1 = 12
+ xrcrg2 = 1
+ k2we = 5e-5
+ prt = 0
+ pua = 4.226297e-23
+ pub = -4.4156209e-32
+ puc = -1.0695581e-23
+ pud = 0
+ ngcon = 1
+ wpclm = 9.3989653e-8
+ dsub = 0.75
+ rsh = 17.5
+ tcj = 0.00076
+ dtox = 2.7e-10
+ ua1 = 1.720591e-9
+ ub1 = -9.5473708e-19
+ uc1 = 7.0015137e-11
+ ppdiblc2 = -6.6555967e-15
+ tpb = 0.0014
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ wa0 = -4.9804098e-8
+ gbmin = 1e-12
+ ute = -1
+ wat = 0.078525419
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 2.0146831e-9
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ wtvoff = -3.0649189e-11
+ wlc = 0
+ wln = 1
+ wu0 = -1.2661044e-9
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -1.3568102e-16
+ wub = 1.003525e-25
+ wuc = -1.2660669e-18
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ eta0 = 0.24044444
+ etab = -0.28088889
+ )

.model nch_sf_27 nmos (
+ level = 54
+ ntox = 1.0
+ pcit = -1.0405802e-16
+ pclm = 1.5094578
+ fnoimod = 1
+ phin = 0.15
+ eigbinv = 1.1
+ pbswd = 0.8
+ pbsws = 0.8
+ pkt1 = 4.636844300000001e-15
+ pkt2 = 2.2738921e-15
+ pdits = 0
+ rbdb = 50
+ pua1 = -2.6369043e-23
+ prwb = 0
+ prwg = 0
+ pub1 = 4.8919292e-32
+ cigsd = 0.069865
+ puc1 = 6.8677984e-24
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ dvt0w = 0
+ pvag = 1.2
+ dvt1w = 0
+ dvt2w = 0
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ rdsw = 100
+ ijthsfwd = 0.01
+ cigbacc = 0.32875
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ tnoimod = 0
+ tnoia = 0
+ ijthsrev = 0.01
+ cigbinv = 0.006
+ peta0 = 0.0
+ rshg = 15.6
+ wketa = -2.2122195e-8
+ wtvfbsdoff = 0
+ tpbsw = 0.0019
+ toxref = 3e-9
+ cjswd = 8.6592e-11
+ cjsws = 8.6592e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ version = 4.5
+ ltvfbsdoff = 0
+ tempmod = 0
+ ppdiblc2 = 1.7501102e-15
+ tnom = 25
+ aigbacc = 0.02
+ tvfbsdoff = 0.022
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ ltvoff = 1.3913801e-9
+ ags = 0.41766657
+ scref = 1e-6
+ cjd = 0.001432992
+ cit = 0.00059502911
+ cjs = 0.001432992
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 9.8024918e-9
+ pigcd = 2.621
+ k3b = 1.9326
+ aigsd = 0.010772818
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ ptvfbsdoff = 0
+ aigbinv = 0.0163
+ lvoff = -4.8532203e-10
+ wags = 3.9284036e-7
+ lku0we = 2.5e-11
+ pkvth0we = -1.3e-19
+ la0 = 3.6355951e-7
+ epsrox = 3.9
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.052658453
+ kt1 = -0.19312528
+ lk2 = -1.4722356e-8
+ kt2 = -0.039065148
+ wcit = 2.7846529999999997e-10
+ lvsat = 0.00016
+ llc = 0
+ lln = 1
+ lu0 = -1.7556993e-9
+ mjd = 0.26
+ lvth0 = -7.8158156e-9
+ lua = -1.1159069e-16
+ mjs = 0.26
+ lub = -2.3732546e-26
+ luc = -2.9405776e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ voff = -0.14601446
+ njs = 1.02
+ pa0 = -3.8856002e-13
+ nsd = 1e+20
+ delta = 0.007595625
+ acde = 0.4
+ pbd = 0.52
+ wvfbsdoff = 0
+ pat = -8.392236300000001e-10
+ pbs = 0.52
+ rdsmod = 0
+ pk2 = 1.1847359e-15
+ lvfbsdoff = 0
+ laigc = -3.3762752e-11
+ pu0 = 1.2848191e-16
+ vfbsdoff = 0.02
+ igbmod = 1
+ prt = 0
+ pua = 2.9945529e-23
+ pub = -3.9782718e-32
+ puc = 6.3626704e-24
+ pud = 0
+ vsat = 102889.02
+ wint = 0
+ rnoia = 0
+ rnoib = 0
+ vth0 = 0.45257959
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 6.6639379e-10
+ ub1 = 1.1665789e-19
+ uc1 = 5.9635906e-11
+ wkt1 = -3.0661037e-8
+ wkt2 = -8.3325526e-9
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ tpb = 0.0014
+ wmax = 5.426e-7
+ wa0 = 7.714643e-7
+ aigc = 0.01167393
+ wmin = 2.726e-7
+ ute = -1
+ wat = 0.0079246317
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -8.8268726e-10
+ pbswgd = 0.95
+ pketa = 1.3732256e-14
+ poxedge = 1
+ pbswgs = 0.95
+ ngate = 8e+20
+ wlc = 0
+ wln = 1
+ wu0 = -1.2259767e-9
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -1.218412e-16
+ wub = 9.5438468e-26
+ wuc = -2.0432641e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ ngcon = 1
+ paramchk = 1
+ wpclm = 9.3989653e-8
+ igcmod = 1
+ binunit = 2
+ wua1 = 4.4082452e-17
+ wub1 = -1.420039e-25
+ wuc1 = -1.718815e-17
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ bigc = 0.001442
+ wwlc = 0
+ cdsc = 0
+ ijthdfwd = 0.01
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ permod = 1
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ ijthdrev = 0.01
+ tvoff = -0.0014023534
+ lpdiblc2 = -7.3119259e-9
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ voffcv = -0.16942
+ wpemod = 1
+ k2we = 5e-5
+ ku0we = -0.0007
+ dsub = 0.75
+ dtox = 2.7e-10
+ beta0 = 13
+ leta0 = -1.6000000000000003e-9
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ njtsswg = 9
+ lkvth0we = -2e-12
+ eta0 = 0.24044444
+ etab = -0.28088889
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.039504569
+ pdiblcb = -0.3
+ tpbswg = 0.0009
+ acnqsmod = 0
+ dmcgt = 0
+ tcjsw = 0.000357
+ rbodymod = 0
+ ptvoff = -5.8159511e-16
+ bigbacc = 0.002588
+ waigsd = 3.1113143e-12
+ bigsd = 0.00125
+ a0 = 0.37817284
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 204899.36
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.02415059
+ k3 = -1.8419
+ em = 1000000.0
+ kvth0we = 0.00018
+ diomod = 1
+ ll = 0
+ lw = 0
+ u0 = 0.017652646
+ w0 = 0
+ wvoff = 1.6091259e-8
+ ua = -1.8479686e-9
+ ub = 2.1067376e-18
+ uc = 1.1966909e-10
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 3.4e-9
+ lintnoi = -1.5e-8
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 2.9779200000000003e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.9779200000000003e-10
+ bigbinv = 0.004953
+ wvsat = -0.0028059037
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ wvth0 = -1.8899760999999997e-8
+ wpdiblc2 = -3.7127843e-9
+ waigc = 2.313153e-11
+ mjswgd = 0.85
+ mjswgs = 0.85
+ lketa = -4.8021757e-8
+ tcjswg = 0.001
+ xpart = 1
+ pvfbsdoff = 0
+ keta = 0.03621471
+ egidl = 0.29734
+ wkvth0we = 2e-12
+ lags = 4.1799271e-7
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 3.8498897000000005e-10
+ trnqsmod = 0
+ kt1l = 0
+ nfactor = 1
+ lint = 6.5375218e-9
+ fprout = 300
+ lkt1 = -1.6493643e-8
+ lkt2 = -1.6288295e-8
+ xrcrg1 = 12
+ xrcrg2 = 1
+ lmax = 8.9908e-7
+ lmin = 4.4908e-7
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ rgatemod = 0
+ wtvoff = 9.3241971e-10
+ pvoff = -4.6372513e-15
+ minv = -0.3
+ tnjtsswg = 1
+ lua1 = 4.5439491e-17
+ lub1 = -2.6569927e-25
+ luc1 = 3.3118724e-18
+ cdscb = 0
+ cdscd = 0
+ nigbacc = 10
+ ndep = 1e+18
+ pvsat = 1.44e-11
+ wk2we = 5e-12
+ pvth0 = 6.0809158e-15
+ lwlc = 0
+ drout = 0.56
+ moin = 5.1
+ capmod = 2
+ paigc = -4.5341069e-18
+ nigc = 3.083
+ voffl = 0
+ wku0we = 2e-11
+ nigbinv = 10
+ mobmod = 0
+ weta0 = -1.1162667e-8
+ wetab = 2.2325333e-8
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ pags = -2.4281917e-13
+ cgidl = 0.22
+ )

.model nch_sf_28 nmos (
+ level = 54
+ wuc1 = -1.3268706e-17
+ bigc = 0.001442
+ ppclm = -7.9196439e-14
+ wwlc = 0
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ cdsc = 0
+ bigbacc = 0.002588
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ wtvfbsdoff = 0
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ kvth0we = 0.00018
+ dmcgt = 0
+ tcjsw = 0.000357
+ wkvth0we = 2e-12
+ lintnoi = -1.5e-8
+ ltvfbsdoff = 0
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ trnqsmod = 0
+ toxref = 3e-9
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ bigsd = 0.00125
+ wvoff = 4.8567953e-9
+ k2we = 5e-5
+ dsub = 0.75
+ wvsat = -0.0054199005
+ dtox = 2.7e-10
+ ptvfbsdoff = 0
+ wvth0 = -1.2869543000000001e-9
+ rgatemod = 0
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ tnjtsswg = 1
+ waigc = -1.6608588e-12
+ ltvoff = -7.6859018e-11
+ eta0 = 0.24044444
+ etab = -0.28088889
+ lketa = -5.7215427e-9
+ nfactor = 1
+ xpart = 1
+ pvfbsdoff = 0
+ lku0we = 2.5e-11
+ egidl = 0.29734
+ epsrox = 3.9
+ rdsmod = 0
+ igbmod = 1
+ nigbacc = 10
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ pbswgd = 0.95
+ pbswgs = 0.95
+ igcmod = 1
+ nigbinv = 10
+ pvoff = 3.0591262e-16
+ cdscb = 0
+ cdscd = 0
+ pvsat = 1.1645586000000001e-9
+ wk2we = 5e-12
+ pvth0 = -1.6687192000000002e-15
+ drout = 0.56
+ paigc = 6.374544e-18
+ ijthsfwd = 0.01
+ paigsd = 2.2627557e-23
+ voffl = 0
+ fnoimod = 1
+ eigbinv = 1.1
+ keta = -0.05992214
+ weta0 = -1.1162667e-8
+ wetab = 2.2325333e-8
+ permod = 1
+ lpclm = 1.4504842e-7
+ lags = 5.906061e-7
+ jswd = 1.28e-13
+ ijthsrev = 0.01
+ jsws = 1.28e-13
+ lcit = 1.01365571e-10
+ cgidl = 0.22
+ kt1l = 0
+ lint = 9.7879675e-9
+ voffcv = -0.16942
+ wpemod = 1
+ lkt1 = 8.6203069e-9
+ lkt2 = -2.5638367e-9
+ lmax = 4.4908e-7
+ cigbacc = 0.32875
+ pbswd = 0.8
+ pbsws = 0.8
+ lmin = 2.1577e-7
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ ppdiblc2 = -5.242001e-17
+ tnoimod = 0
+ minv = -0.3
+ lua1 = -4.6794128e-17
+ lub1 = -3.0489654e-26
+ luc1 = -2.1335001e-17
+ pdits = 0
+ ndep = 1e+18
+ cigsd = 0.069865
+ cigbinv = 0.006
+ dvt0w = 0
+ lwlc = 0
+ dvt1w = 0
+ dvt2w = 0
+ moin = 5.1
+ nigc = 3.083
+ tpbswg = 0.0009
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ version = 4.5
+ tempmod = 0
+ pkvth0we = -1.3e-19
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ tnoia = 0
+ pags = 1.2428184e-13
+ peta0 = 0.0
+ ptvoff = -1.5558646e-16
+ aigbacc = 0.02
+ ntox = 1.0
+ pcit = 3.0152771000000005e-18
+ pclm = 1.1798023
+ waigsd = 3.1112628e-12
+ wketa = 2.3981389e-8
+ vfbsdoff = 0.02
+ tpbsw = 0.0019
+ cjswd = 8.6592e-11
+ cjsws = 8.6592e-11
+ diomod = 1
+ mjswd = 0.11
+ phin = 0.15
+ mjsws = 0.11
+ agidl = 9.41e-8
+ pditsd = 0
+ pditsl = 0
+ aigbinv = 0.0163
+ pkt1 = -1.2676052e-14
+ pkt2 = -7.0784646e-16
+ cjswgd = 2.9779200000000003e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.9779200000000003e-10
+ paramchk = 1
+ ags = 0.025363416000000014
+ cjd = 0.001432992
+ tvfbsdoff = 0.022
+ cit = 0.0012396277
+ cjs = 0.001432992
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 1.30529375e-8
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ rbdb = 50
+ pua1 = 1.8291934e-23
+ prwb = 0
+ prwg = 0
+ pub1 = -6.3924188e-33
+ puc1 = 5.143243e-24
+ mjswgd = 0.85
+ mjswgs = 0.85
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ tcjswg = 0.001
+ rdsw = 100
+ scref = 1e-6
+ ijthdfwd = 0.01
+ la0 = -6.0902319e-7
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.014956938
+ kt1 = -0.25020244
+ lk2 = -1.0681005e-8
+ kt2 = -0.070257098
+ pigcd = 2.621
+ llc = -1.18e-13
+ lln = 0.7
+ aigsd = 0.010772818
+ lu0 = -7.0983626e-10
+ mjd = 0.26
+ lua = -1.8564943e-17
+ mjs = 0.26
+ lub = -5.2748233e-26
+ luc = -4.2757753e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 2.2627554e-14
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 2.5781001e-9
+ poxedge = 1
+ pbs = 0.52
+ pk2 = 8.6250113e-16
+ lvoff = -7.1314494000000004e-9
+ a0 = 2.5885881
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ pu0 = 4.9938272000000003e-17
+ at = 119214.09
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.014965692000000001
+ k3 = -1.8419
+ em = 1000000.0
+ prt = 0
+ pua = 5.6394132e-24
+ pub = -7.710339e-34
+ puc = -1.5613012e-24
+ pud = 0
+ ll = -1.18e-13
+ lw = 0
+ u0 = 0.015275684000000001
+ w0 = 0
+ ua = -2.0593908e-9
+ ub = 2.1726824e-18
+ uc = 6.2555449e-11
+ ud = 0
+ wl = 0
+ rsh = 17.5
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 3.4e-9
+ tcj = 0.00076
+ ua1 = 8.7601565e-10
+ lvsat = -0.0040072412
+ ub1 = -4.1790941e-19
+ uc1 = 1.1565153e-10
+ binunit = 2
+ lvth0 = 1.8743980000000003e-9
+ ijthdrev = 0.01
+ tpb = 0.0014
+ wvfbsdoff = 0
+ wa0 = -1.6305293e-7
+ lvfbsdoff = 0
+ ute = -1
+ wat = 0.00015798693
+ delta = 0.007595625
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -1.5033038e-10
+ laigc = -3.7429738e-11
+ wlc = 0
+ wln = 1
+ rshg = 15.6
+ wu0 = -1.0474684e-9
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -6.6600022e-17
+ wub = 6.7755498e-27
+ wuc = -2.4236148e-18
+ wud = 0
+ lpdiblc2 = -4.2799755e-9
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ rnoia = 0
+ rnoib = 0
+ fprout = 300
+ xrcrg1 = 12
+ xrcrg2 = 1
+ pketa = -6.5533207e-15
+ ngate = 8e+20
+ ngcon = 1
+ wpclm = 2.7398156e-7
+ wtvoff = -3.5781771e-11
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ tnom = 25
+ jswgs = 1.28e-13
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ lkvth0we = -2e-12
+ capmod = 2
+ wku0we = 2e-11
+ mobmod = 0
+ acnqsmod = 0
+ wags = -4.4148013e-7
+ wcit = 3.5116891e-11
+ rbodymod = 0
+ voff = -0.13090963
+ acde = 0.4
+ tvoff = 0.0019345538
+ njtsswg = 9
+ vsat = 112360.02
+ wint = 0
+ xjbvd = 1
+ xjbvs = 1
+ vth0 = 0.43055638
+ lk2we = -1.5e-12
+ wkt1 = 8.6864548e-9
+ wkt2 = -1.5558741e-9
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ wmax = 5.426e-7
+ laigsd = -8.1983894e-17
+ aigc = 0.011682264
+ wmin = 2.726e-7
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.032613772
+ pdiblcb = -0.3
+ ku0we = -0.0007
+ beta0 = 13
+ leta0 = -1.6000000000000003e-9
+ wua1 = -5.7419768e-17
+ wpdiblc2 = 3.8387521e-10
+ wub1 = -1.6295463e-26
+ )

.model nch_sf_29 nmos (
+ level = 54
+ keta = 0.0092481698
+ aigbinv = 0.0163
+ tnoia = 0
+ ijthdrev = 0.01
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = -5.537106000000001e-12
+ peta0 = 0.0
+ ptvfbsdoff = 0
+ kt1l = 0
+ wketa = -2.0169501e-8
+ toxref = 3e-9
+ lpdiblc2 = -9.0824285e-10
+ tpbsw = 0.0019
+ ags = 2.8244444
+ cjswd = 8.6592e-11
+ cjsws = 8.6592e-11
+ lint = 9.7879675e-9
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ cjd = 0.001432992
+ cit = 0.0017462755
+ cjs = 0.001432992
+ clc = 1e-7
+ cle = 0.6
+ lkt1 = -2.7662126e-9
+ bvd = 8.7
+ lkt2 = -3.9513595e-9
+ bvs = 8.7
+ lmax = 2.1577e-7
+ dlc = 1.30529375e-8
+ lmin = 9e-8
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ poxedge = 1
+ tvfbsdoff = 0.022
+ la0 = -2.075695e-7
+ minv = -0.3
+ jsd = 6.11e-7
+ ltvoff = 5.8839234e-11
+ jss = 6.11e-7
+ lat = -0.0015137311
+ lua1 = -5.8912951e-18
+ lub1 = -2.6977439000000003e-26
+ luc1 = 7.212716e-18
+ kt1 = -0.1962379
+ lk2 = -3.2022951e-9
+ kt2 = -0.063681161
+ llc = -1.18e-13
+ binunit = 2
+ lln = 0.7
+ lu0 = -2.5951767e-10
+ mjd = 0.26
+ lua = 5.2959027e-17
+ mjs = 0.26
+ lub = -7.97606935e-26
+ luc = -8.8267893e-18
+ lud = 0
+ lwc = 0
+ ndep = 1e+18
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ lkvth0we = -2e-12
+ njs = 1.02
+ pa0 = 1.0407708e-13
+ nsd = 1e+20
+ lwlc = 0
+ pbd = 0.52
+ pat = -3.5721950999999997e-10
+ pbs = 0.52
+ pk2 = -9.7578421e-17
+ moin = 5.1
+ pu0 = 1.7060797e-17
+ prt = 0
+ pua = -7.1102082e-24
+ pub = 9.57267e-33
+ puc = 7.19078e-25
+ pud = 0
+ scref = 1e-6
+ nigc = 3.083
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 6.8216336e-10
+ pigcd = 2.621
+ ub1 = -4.3455498e-19
+ uc1 = -1.9645420999999998e-11
+ aigsd = 0.010772818
+ tpb = 0.0014
+ lku0we = 2.5e-11
+ wa0 = -5.4906963e-7
+ acnqsmod = 0
+ ute = -1
+ wat = 0.014069454
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 4.3998097e-9
+ epsrox = 3.9
+ lvoff = 2.34836653e-9
+ wlc = 0
+ wln = 1
+ wu0 = -8.9165099e-10
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -6.1752756e-18
+ wub = -4.2246744000000004e-26
+ wuc = -1.3231099e-17
+ wud = 0
+ wwc = 0
+ noff = 2.7195
+ wwl = 0
+ wwn = 1
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ lvsat = -0.00029734827
+ rbodymod = 0
+ rdsmod = 0
+ wvfbsdoff = 0
+ lvth0 = -1.1794990599999998e-8
+ lvfbsdoff = 0
+ igbmod = 1
+ delta = 0.007595625
+ laigc = 2.6175146e-12
+ ntox = 1.0
+ pcit = 1.9820824800000002e-17
+ jtsswgd = 2.3e-7
+ pclm = 2.3689724
+ jtsswgs = 2.3e-7
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ rnoia = 0
+ rnoib = 0
+ pbswgd = 0.95
+ pbswgs = 0.95
+ phin = 0.15
+ pketa = 2.762517e-15
+ ngate = 8e+20
+ igcmod = 1
+ ngcon = 1
+ pkt1 = 4.8916645e-16
+ pkt2 = 9.3582987e-16
+ wpclm = -2.0834879e-7
+ wpdiblc2 = 1.3111248e-10
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ rbdb = 50
+ pua1 = 1.9734917e-24
+ prwb = 0
+ prwg = 0
+ pub1 = -5.0622001000000004e-33
+ puc1 = -3.1412237000000002e-24
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ njtsswg = 9
+ paigsd = -9.4615512e-24
+ rdsw = 100
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ permod = 1
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.016633997
+ pdiblcb = -0.3
+ wkvth0we = 2e-12
+ trnqsmod = 0
+ tvoff = 0.0012914341
+ rshg = 15.6
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ voffcv = -0.16942
+ wpemod = 1
+ bigbacc = 0.002588
+ ku0we = -0.0007
+ kvth0we = 0.00018
+ beta0 = 13
+ leta0 = -1.6000000000000003e-9
+ rgatemod = 0
+ lintnoi = -1.5e-8
+ tnjtsswg = 1
+ tnom = 25
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ ppclm = 2.2575265e-14
+ vtsswgs = 4.2
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ tpbswg = 0.0009
+ dmcgt = 0
+ wags = 1.4753332999999998e-7
+ tcjsw = 0.000357
+ wcit = -4.4530253800000005e-11
+ ptvoff = 2.7225835e-17
+ voff = -0.175837897
+ waigsd = 3.1114149e-12
+ acde = 0.4
+ vsat = 94777.65030000001
+ wint = 0
+ bigsd = 0.00125
+ vth0 = 0.49534045399999993
+ diomod = 1
+ wkt1 = -5.3707946e-8
+ wkt2 = -9.3458092e-9
+ wmax = 5.426e-7
+ aigc = 0.011492467
+ wmin = 2.726e-7
+ nfactor = 1
+ pditsd = 0
+ pditsl = 0
+ wvoff = 8.6692167e-9
+ cjswgd = 2.9779200000000003e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.9779200000000003e-10
+ wvsat = -0.0005775380999999999
+ wvth0 = -1.4725728e-8
+ wua1 = 1.991882e-17
+ wub1 = -2.2599817e-26
+ wuc1 = 2.5994103e-17
+ waigc = 3.9031408e-11
+ bigc = 0.001442
+ mjswgd = 0.85
+ mjswgs = 0.85
+ wwlc = 0
+ tcjswg = 0.001
+ nigbacc = 10
+ lketa = -2.0316478e-8
+ cdsc = 0
+ ijthsfwd = 0.01
+ cgbo = 0
+ xpart = 1
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ pvfbsdoff = 0
+ xtid = 3
+ xtis = 3
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ egidl = 0.29734
+ nigbinv = 10
+ ijthsrev = 0.01
+ fprout = 300
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ fnoimod = 1
+ k2we = 5e-5
+ wtvoff = -9.0219076e-10
+ eigbinv = 1.1
+ dsub = 0.75
+ dtox = 2.7e-10
+ ppdiblc2 = 9.1292629e-19
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ pvoff = -4.985090499999997e-16
+ a0 = 0.68596391
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 55502.213
+ cf = 8.15e-11
+ cdscb = 0
+ cdscd = 0
+ ef = 1.0
+ k1 = 0.274
+ k2 = -0.02047843
+ k3 = -1.8419
+ em = 1000000.0
+ ll = -1.18e-13
+ lw = 0
+ u0 = 0.013141473
+ pvsat = 1.4282156000000005e-10
+ w0 = 0
+ ua = -2.398367e-9
+ ub = 2.300703286e-18
+ uc = 8.4124236e-11
+ ud = 0
+ wk2we = 5e-12
+ capmod = 2
+ wl = 0
+ wr = 1
+ pvth0 = 1.1668619999999998e-15
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ eta0 = 0.24044444
+ xw = 3.4e-9
+ drout = 0.56
+ etab = -0.28088889
+ wku0we = 2e-11
+ paigc = -2.2115244e-18
+ mobmod = 0
+ voffl = 0
+ cigbacc = 0.32875
+ weta0 = -1.1162667e-8
+ wetab = 2.2325333e-8
+ pkvth0we = -1.3e-19
+ lpclm = -1.0586647e-7
+ tnoimod = 0
+ cgidl = 0.22
+ vfbsdoff = 0.02
+ cigbinv = 0.006
+ laigsd = 3.4280989e-17
+ pbswd = 0.8
+ pbsws = 0.8
+ paramchk = 1
+ version = 4.5
+ wtvfbsdoff = 0
+ tempmod = 0
+ pdits = 0
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ cigsd = 0.069865
+ ltvfbsdoff = 0
+ dvt0w = 0
+ aigbacc = 0.02
+ dvt1w = 0
+ dvt2w = 0
+ ijthdfwd = 0.01
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ )

.model nch_sf_30 nmos (
+ level = 54
+ keta = -0.29566775
+ aigbinv = 0.0163
+ tnoia = 0
+ ijthdrev = 0.01
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 1.8234428e-10
+ peta0 = -9.3037135e-16
+ ptvfbsdoff = 0
+ petab = -1.2138265e-15
+ kt1l = 0
+ wketa = -4.7865407e-8
+ toxref = 3e-9
+ lpdiblc2 = 8.2379047e-15
+ tpbsw = 0.0019
+ ags = 2.8244444
+ cjswd = 8.6592e-11
+ cjsws = 8.6592e-11
+ lint = 0
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ cjd = 0.001432992
+ cit = -0.00025246267
+ cjs = 0.001432992
+ clc = 1e-7
+ cle = 0.6
+ lkt1 = -8.735083599999999e-9
+ bvd = 8.7
+ lkt2 = 3.8424987e-10
+ bvs = 8.7
+ lmax = 9e-8
+ dlc = 3.26497e-9
+ lmin = 5.4e-8
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ poxedge = 1
+ tvfbsdoff = 0.022
+ la0 = 3.9829889e-7
+ minv = -0.3
+ jsd = 6.11e-7
+ ltvoff = -2.7237524e-10
+ jss = 6.11e-7
+ lat = 0.00536560498
+ lua1 = -1.2736334e-17
+ lub1 = 1.8485594000000001e-26
+ luc1 = 3.67094421e-18
+ kt1 = -0.13273927
+ lk2 = 1.0502722e-9
+ kt2 = -0.10980467
+ llc = 0
+ binunit = 2
+ lln = 1
+ lu0 = -2.0875966000000002e-10
+ mjd = 0.26
+ lua = -7.6887484e-18
+ mjs = 0.26
+ lub = 6.3606825e-27
+ luc = -3.2720592999999998e-18
+ lud = 0
+ lwc = 0
+ ndep = 1e+18
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ lkvth0we = -2e-12
+ njs = 1.02
+ pa0 = -1.1411036e-13
+ nsd = 1e+20
+ lwlc = 0
+ pbd = 0.52
+ pat = -1.7176563e-9
+ pbs = 0.52
+ pk2 = -3.7289588e-16
+ moin = 5.1
+ pu0 = 7.1384501e-17
+ prt = 0
+ pua = 1.3044266e-23
+ pub = -1.13966382e-32
+ puc = 2.3653651e-24
+ pud = 0
+ scref = 1e-6
+ nigc = 3.083
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 7.5498293e-10
+ pigcd = 2.621
+ ub1 = -9.1820427e-19
+ uc1 = 1.8032940999999987e-11
+ aigsd = 0.010772818
+ tpb = 0.0014
+ lku0we = 2.5e-11
+ wa0 = 1.7720733e-6
+ acnqsmod = 0
+ ute = -1
+ wat = 0.028542186400000003
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 7.3287188e-9
+ epsrox = 3.9
+ lvoff = -3.2351799e-9
+ wlc = 0
+ wln = 1
+ wu0 = -1.4695626999999999e-9
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -2.2058458e-16
+ wub = 1.80830997e-25
+ wuc = -3.0744792e-17
+ wud = 0
+ wwc = 0
+ noff = 2.7195
+ wwl = 0
+ wwn = 1
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ lvsat = 0.0037119283000000003
+ rbodymod = 0
+ rdsmod = 0
+ wvfbsdoff = 0
+ lvth0 = 3.989724300000001e-9
+ lvfbsdoff = 0
+ igbmod = 1
+ delta = 0.007595625
+ laigc = -3.0244582e-11
+ ntox = 1.0
+ pcit = -7.457676e-18
+ jtsswgd = 2.3e-7
+ pclm = 1.7776553
+ jtsswgs = 2.3e-7
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ rnoia = 0
+ rnoib = 0
+ pbswgd = 0.95
+ pbswgs = 0.95
+ phin = 0.15
+ pketa = 5.3659323e-15
+ ngate = 8e+20
+ igcmod = 1
+ ngcon = 1
+ pkt1 = 4.9305068e-15
+ pkt2 = -5.9202052e-16
+ wpclm = 4.3365813e-8
+ wpdiblc2 = 1.4083642e-10
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ rbdb = 50
+ pua1 = 4.1884121e-24
+ prwb = 0
+ prwg = 0
+ pub1 = -9.626998799999999e-33
+ puc1 = 1.4280652000000004e-24
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ njtsswg = 9
+ rdsw = 100
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ permod = 1
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.0069717513
+ pdiblcb = -0.3
+ wkvth0we = 2e-12
+ trnqsmod = 0
+ tvoff = 0.0048149924
+ rshg = 15.6
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ voffcv = -0.16942
+ wpemod = 1
+ bigbacc = 0.002588
+ ku0we = -0.0007
+ kvth0we = 0.00018
+ beta0 = 13
+ leta0 = 1.8440248999999998e-8
+ rgatemod = 0
+ letab = -2.6551319e-8
+ lintnoi = -1.5e-8
+ tnjtsswg = 1
+ tnom = 25
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ ppclm = -1.085908e-15
+ vtsswgs = 4.2
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ tpbswg = 0.0009
+ dmcgt = 0
+ wags = 1.4753332999999998e-7
+ tcjsw = 0.000357
+ wcit = 2.4566655999999997e-10
+ ptvoff = 9.0058483e-17
+ voff = -0.116438471
+ waigsd = 3.1113143e-12
+ acde = 0.4
+ vsat = 52125.77300000001
+ wint = 0
+ bigsd = 0.00125
+ vth0 = 0.327417953
+ diomod = 1
+ wkt1 = -1.0095625e-7
+ wkt2 = 6.9079183e-9
+ wmax = 5.426e-7
+ aigc = 0.011842064
+ wmin = 2.726e-7
+ nfactor = 1
+ pditsd = 0
+ pditsl = 0
+ wvoff = 3.9876867999999985e-9
+ cjswgd = 2.9779200000000003e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.9779200000000003e-10
+ wvsat = 0.0060216695
+ wvth0 = -4.325777100000002e-9
+ wua1 = -3.6441631e-18
+ wub1 = 2.5961869999999995e-26
+ wuc1 = -2.2615369999999997e-17
+ waigc = 4.5087747e-12
+ bigc = 0.001442
+ mjswgd = 0.85
+ mjswgs = 0.85
+ wwlc = 0
+ tcjswg = 0.001
+ nigbacc = 10
+ lketa = 8.345618e-9
+ cdsc = 0
+ ijthsfwd = 0.01
+ cgbo = 0
+ xpart = 1
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ pvfbsdoff = 0
+ xtid = 3
+ xtis = 3
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ egidl = 0.29734
+ nigbinv = 10
+ ijthsrev = 0.01
+ fprout = 300
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ fnoimod = 1
+ k2we = 5e-5
+ wtvoff = -1.5706231e-9
+ eigbinv = 1.1
+ dsub = 0.75
+ dtox = 2.7e-10
+ ppdiblc2 = -1.1241984e-21
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ pvoff = -5.844511799999985e-17
+ a0 = -5.7594444
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = -17682.2125
+ cf = 8.15e-11
+ cdscb = 0
+ cdscd = 0
+ ef = 1.0
+ k1 = 0.274
+ k2 = -0.065718509
+ k3 = -1.8419
+ em = 1000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.012601494000000001
+ pvsat = -4.77504e-10
+ w0 = 0
+ ua = -1.7531779e-9
+ ub = 1.3845184050000002e-18
+ uc = 2.5031363e-11
+ ud = 0
+ wk2we = 5e-12
+ capmod = 2
+ wl = 0
+ wr = 1
+ pvth0 = 1.8926666000000022e-16
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ eta0 = 0.027250304
+ xw = 3.4e-9
+ drout = 0.56
+ etab = 0.001571952
+ wku0we = 2e-11
+ paigc = 1.0336032e-18
+ mobmod = 0
+ voffl = 0
+ cigbacc = 0.32875
+ weta0 = -1.2650991e-9
+ wetab = 3.5238381e-8
+ pkvth0we = -1.3e-19
+ lpclm = -5.0282662e-8
+ tnoimod = 0
+ cgidl = 0.22
+ vfbsdoff = 0.02
+ cigbinv = 0.006
+ pbswd = 0.8
+ pbsws = 0.8
+ paramchk = 1
+ version = 4.5
+ wtvfbsdoff = 0
+ tempmod = 0
+ pdits = 0
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ cigsd = 0.069865
+ ltvfbsdoff = 0
+ dvt0w = 0
+ aigbacc = 0.02
+ dvt1w = 0
+ dvt2w = 0
+ ijthdfwd = 0.01
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ )

.model nch_sf_31 nmos (
+ level = 54
+ nigbacc = 10
+ wvoff = 2.2964685300000028e-9
+ wvsat = 0.019777184200000006
+ wvth0 = -2.7887312999999994e-8
+ ltvoff = 2.6647905e-10
+ waigc = 1.8753243e-11
+ tnom = 25
+ nigbinv = 10
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ lketa = -2.3617222e-8
+ pvfbsdoff = 0
+ xpart = 1
+ lku0we = 2.5e-11
+ epsrox = 3.9
+ egidl = 0.29734
+ fnoimod = 1
+ pkvth0we = -1.3e-19
+ wags = 1.4753332999999998e-7
+ rdsmod = 0
+ eigbinv = 1.1
+ wcit = 3.3128934e-10
+ igbmod = 1
+ voff = -0.07382279000000001
+ acde = 0.4
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ vfbsdoff = 0.02
+ vsat = 48765.08000000001
+ pbswgd = 0.95
+ pbswgs = 0.95
+ wint = 0
+ vth0 = 0.34682439000000004
+ wkt1 = -1.4134348999999998e-8
+ wkt2 = -2.0876247e-8
+ wmax = 5.426e-7
+ igcmod = 1
+ aigc = 0.011696193
+ wmin = 2.726e-7
+ paramchk = 1
+ cigbacc = 0.32875
+ wua1 = -1.1132499e-16
+ wub1 = 7.746802000000003e-26
+ wuc1 = 6.392091000000002e-17
+ pvoff = 3.964544000000059e-17
+ bigc = 0.001442
+ cdscb = 0
+ cdscd = 0
+ tnoimod = 0
+ wwlc = 0
+ pvsat = -1.275324e-9
+ wk2we = 5e-12
+ pvth0 = 1.5558357999999996e-15
+ drout = 0.56
+ paigsd = 1.7624612e-23
+ cdsc = 0
+ paigc = 2.0742404e-19
+ cigbinv = 0.006
+ ijthdfwd = 0.01
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ voffl = 0
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ permod = 1
+ weta0 = -1.2005104e-7
+ wetab = 5.6750807e-8
+ lpclm = 5.458214e-8
+ version = 4.5
+ tempmod = 0
+ ijthdrev = 0.01
+ cgidl = 0.22
+ voffcv = -0.16942
+ wpemod = 1
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ aigbacc = 0.02
+ pbswd = 0.8
+ pbsws = 0.8
+ k2we = 5e-5
+ dsub = 0.75
+ dtox = 2.7e-10
+ aigbinv = 0.0163
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ pdits = 0
+ cigsd = 0.069865
+ lkvth0we = -2e-12
+ eta0 = 1.0176617
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ etab = -1.3959412
+ tpbswg = 0.0009
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ acnqsmod = 0
+ tnoia = 0
+ ptvoff = -4.401556e-18
+ poxedge = 1
+ rbodymod = 0
+ ags = 2.8244444
+ waigsd = 3.1110104e-12
+ peta0 = 5.9592132e-15
+ cjd = 0.001432992
+ cit = -0.0053709179
+ cjs = 0.001432992
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ petab = -2.4615472e-15
+ dlc = 3.26497e-9
+ binunit = 2
+ wketa = -5.877032e-8
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ diomod = 1
+ tpbsw = 0.0019
+ cjswd = 8.6592e-11
+ cjsws = 8.6592e-11
+ mjswd = 0.11
+ pditsd = 0
+ pditsl = 0
+ mjsws = 0.11
+ agidl = 9.41e-8
+ cjswgd = 2.9779200000000003e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.9779200000000003e-10
+ la0 = -1.4097724e-8
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.0006394376999999999
+ kt1 = -0.39757001
+ lk2 = 7.4338958e-10
+ kt2 = -0.14677127
+ llc = 0
+ lln = 1
+ lu0 = 5.0370058e-10
+ mjd = 0.26
+ lua = 6.4763643e-17
+ mjs = 0.26
+ lub = -2.3096342000000002e-26
+ luc = -1.0931136000000001e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = -1.7333804e-13
+ nsd = 1e+20
+ pbd = 0.52
+ pat = -4.2349470999999994e-10
+ tvfbsdoff = 0.022
+ pbs = 0.52
+ pk2 = -1.0803308e-16
+ wpdiblc2 = 1.4081704e-10
+ pu0 = -4.7327483e-17
+ prt = 0
+ pua = -2.1774501e-24
+ pub = -5.473259300000002e-33
+ puc = 4.761497700000001e-24
+ pud = 0
+ mjswgd = 0.85
+ mjswgs = 0.85
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 1.4910078e-9
+ ub1 = -1.7286540799999999e-18
+ uc1 = -3.206985999999997e-11
+ tpb = 0.0014
+ tcjswg = 0.001
+ wa0 = 2.7932403e-6
+ ute = -1
+ wat = 0.006229054600000004
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 2.7621189e-9
+ wlc = 0
+ wln = 1
+ wu0 = 5.771956e-10
+ jtsswgd = 2.3e-7
+ xgl = -1.09e-8
+ jtsswgs = 2.3e-7
+ xgw = 0
+ wua = 4.1858808e-17
+ wub = 7.870378029999999e-26
+ wuc = -7.2057435e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ scref = 1e-6
+ pigcd = 2.621
+ aigsd = 0.010772819
+ keta = 0.2554158
+ lvoff = -5.706889800000001e-9
+ wkvth0we = 2e-12
+ wvfbsdoff = 0
+ lvsat = 0.0039068485699999995
+ lvfbsdoff = 0
+ lvth0 = 2.8641506e-9
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 4.792146899999999e-10
+ trnqsmod = 0
+ delta = 0.007595625
+ laigc = -2.1784105e-11
+ kt1l = 0
+ fprout = 300
+ xrcrg1 = 12
+ xrcrg2 = 1
+ rnoia = 0
+ rnoib = 0
+ lint = 0
+ njtsswg = 9
+ lkt1 = 6.6250994e-9
+ lkt2 = 2.528313e-9
+ pketa = 5.998417e-15
+ ngate = 8e+20
+ lmax = 5.4e-8
+ lmin = 4.5e-8
+ wtvoff = 5.799816e-11
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ ngcon = 1
+ wpclm = 2.4669208e-7
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ ckappad = 0.6
+ ckappas = 0.6
+ rgatemod = 0
+ gbmin = 1e-12
+ pdiblc1 = 0
+ pdiblc2 = 0.0069718933
+ pdiblcb = -0.3
+ tnjtsswg = 1
+ minv = -0.3
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ lua1 = -5.5425775e-17
+ lub1 = 6.549168e-26
+ luc1 = 6.576863000000002e-18
+ capmod = 2
+ ndep = 1e+18
+ wku0we = 2e-11
+ lwlc = 0
+ moin = 5.1
+ mobmod = 0
+ nigc = 3.083
+ bigbacc = 0.002588
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ kvth0we = 0.00018
+ wtvfbsdoff = 0
+ lintnoi = -1.5e-8
+ bigbinv = 0.004953
+ tvoff = -0.0044755986
+ ntox = 1.0
+ vtsswgd = 4.2
+ pcit = -1.2423797e-17
+ vtsswgs = 4.2
+ pclm = -0.030358553
+ laigsd = -6.385731e-17
+ xjbvd = 1
+ a0 = 1.350842
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ xjbvs = 1
+ lk2we = -1.5e-12
+ at = 85853.00300000001
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = -0.060427428000000005
+ k3 = -1.8419
+ em = 1000000.0
+ ltvfbsdoff = 0
+ ll = 0
+ lw = 0
+ u0 = 0.00031769704690000003
+ w0 = 0
+ ua = -3.002357e-9
+ ub = 1.89239813e-18
+ uc = 1.5708441000000004e-10
+ ud = 0
+ phin = 0.15
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 3.4e-9
+ pkt1 = -1.0516334e-16
+ pkt2 = 1.019461e-15
+ ku0we = -0.0007
+ beta0 = 13
+ leta0 = -3.9003611e-8
+ letab = 5.4504443e-8
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ ppclm = -1.2878832e-14
+ rbdb = 50
+ pua1 = 1.04339e-23
+ prwb = 0
+ prwg = 0
+ pub1 = -1.2614356e-32
+ puc1 = -3.591008600000001e-24
+ rbpb = 50
+ rbpd = 50
+ dlcig = 2.5e-9
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ bgidl = 2320000000.0
+ ptvfbsdoff = 0
+ rdsw = 100
+ ijthsfwd = 0.01
+ nfactor = 1
+ dmcgt = 0
+ tcjsw = 0.000357
+ ijthsrev = 0.01
+ toxref = 3e-9
+ rshg = 15.6
+ bigsd = 0.00125
+ )

.model nch_sf_32 nmos (
+ level = 54
+ eta0 = -0.25440451
+ etab = -0.81370191
+ scref = 1e-6
+ lku0we = 2.5e-11
+ pigcd = 2.621
+ epsrox = 3.9
+ aigsd = 0.010772817
+ njtsswg = 9
+ lvoff = -7.215689799999999e-9
+ rdsmod = 0
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ igbmod = 1
+ lvsat = -0.0007652195999999999
+ ckappad = 0.6
+ ckappas = 0.6
+ lvth0 = 3.3208689999999967e-10
+ pdiblc1 = 0
+ pdiblc2 = 0.0069718933
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ pdiblcb = -0.3
+ delta = 0.007595625
+ laigc = 9.707156e-12
+ pbswgd = 0.95
+ pbswgs = 0.95
+ rnoia = 0
+ rnoib = 0
+ igcmod = 1
+ pketa = -6.053668000000001e-15
+ ngate = 8e+20
+ ngcon = 1
+ wpclm = 1.6305740000000013e-7
+ bigbacc = 0.002588
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ kvth0we = 0.00018
+ paigsd = -1.2154906e-23
+ lintnoi = -1.5e-8
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ ijthsfwd = 0.01
+ permod = 1
+ keta = -0.59506219
+ ijthsrev = 0.01
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 1.3559100000000003e-10
+ tvoff = 0.0034020192
+ kt1l = 0
+ voffcv = -0.16942
+ wpemod = 1
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ lint = 0
+ lkt1 = -1.8769946e-8
+ lkt2 = 1.0897551e-9
+ lmax = 4.5e-8
+ lmin = 3.6e-8
+ ku0we = -0.0007
+ nfactor = 1
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ beta0 = 13
+ leta0 = 2.33276322e-8
+ letab = 2.5974719e-8
+ minv = -0.3
+ lua1 = 7.6118385e-17
+ lub1 = -1.2550425000000001e-25
+ luc1 = -3.7246273e-17
+ ppclm = -8.780734400000002e-15
+ ndep = 1e+18
+ dlcig = 2.5e-9
+ lwlc = 0
+ tpbswg = 0.0009
+ bgidl = 2320000000.0
+ moin = 5.1
+ nigc = 3.083
+ nigbacc = 10
+ dmcgt = 0
+ pkvth0we = -1.3e-19
+ noff = 2.7195
+ tcjsw = 0.000357
+ ptvoff = -5.392468e-18
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ waigsd = 3.1116181e-12
+ nigbinv = 10
+ diomod = 1
+ ntox = 1.0
+ pcit = 2.5771809e-17
+ vfbsdoff = 0.02
+ pclm = 1.46768105
+ bigsd = 0.00125
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 2.9779200000000003e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.9779200000000003e-10
+ phin = 0.15
+ wvoff = -1.1428948000000006e-8
+ paramchk = 1
+ pkt1 = 5.1950205000000005e-15
+ pkt2 = -4.1883975e-17
+ wvsat = -0.021295046
+ wvth0 = -2.3056159e-8
+ fnoimod = 1
+ mjswgd = 0.85
+ mjswgs = 0.85
+ eigbinv = 1.1
+ waigc = 7.6854687e-11
+ tcjswg = 0.001
+ rbdb = 50
+ pua1 = -2.7889543e-23
+ prwb = 0
+ prwg = 0
+ pub1 = 4.5182459e-32
+ puc1 = 1.2190150800000001e-23
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ pvfbsdoff = 0
+ lketa = 1.80561909e-8
+ ijthdfwd = 0.01
+ rdsw = 100
+ xpart = 1
+ egidl = 0.29734
+ cigbacc = 0.32875
+ ijthdrev = 0.01
+ fprout = 300
+ rshg = 15.6
+ xrcrg1 = 12
+ xrcrg2 = 1
+ tnoimod = 0
+ cigbinv = 0.006
+ wtvoff = 7.822084e-11
+ pvoff = 7.121929600000003e-16
+ version = 4.5
+ capmod = 2
+ tnom = 25
+ cdscb = 0
+ cdscd = 0
+ tempmod = 0
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ pvsat = 7.372158200000001e-10
+ wku0we = 2e-11
+ lkvth0we = -2e-12
+ wk2we = 5e-12
+ pvth0 = 1.31910679e-15
+ drout = 0.56
+ mobmod = 0
+ wtvfbsdoff = 0
+ paigc = -2.6395467e-18
+ aigbacc = 0.02
+ voffl = 0
+ acnqsmod = 0
+ ltvfbsdoff = 0
+ weta0 = 8.5615058e-8
+ wetab = 2.2270081e-8
+ wags = 1.4753332999999998e-7
+ lpclm = -1.8821805999999992e-8
+ wcit = -4.482130999999999e-10
+ rbodymod = 0
+ aigbinv = 0.0163
+ voff = -0.04303087299999998
+ cgidl = 0.22
+ acde = 0.4
+ laigsd = 4.4039511e-17
+ vsat = 144113.422
+ wint = 0
+ vth0 = 0.398499171
+ wkt1 = -1.2230137e-7
+ wkt2 = 7.8385579e-10
+ wmax = 5.426e-7
+ aigc = 0.011053515
+ wmin = 2.726e-7
+ pbswd = 0.8
+ pbsws = 0.8
+ ptvfbsdoff = 0
+ wpdiblc2 = 1.4081704e-10
+ wua1 = 6.7078609e-16
+ wub1 = -1.1020589000000001e-24
+ wuc1 = -2.5814450999999997e-16
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ poxedge = 1
+ bigc = 0.001442
+ pdits = 0
+ wwlc = 0
+ cigsd = 0.069865
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ binunit = 2
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ ags = 2.8244444
+ cgsl = 3.31989e-12
+ pk2we = -1e-19
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ a0 = 10.55945905
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 101543.357
+ cf = 8.15e-11
+ cjd = 0.001432992
+ cit = 0.0016418092000000002
+ cjs = 0.001432992
+ clc = 1e-7
+ ef = 1.0
+ k1 = 0.274
+ cle = 0.6
+ k2 = 0.040727321999999996
+ k3 = -1.8419
+ em = 1000000.0
+ bvd = 8.7
+ bvs = 8.7
+ ll = 0
+ lw = 0
+ dlc = 3.26497e-9
+ u0 = 0.0106083374
+ w0 = 0
+ k3b = 1.9326
+ ua = -1.7148580999999998e-9
+ ub = 1.250859149999999e-18
+ uc = 5.4381728e-10
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ dwb = 0
+ ww = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ xw = 3.4e-9
+ wkvth0we = 2e-12
+ tnoia = 0
+ toxref = 3e-9
+ peta0 = -4.1184253e-15
+ la0 = -4.65319969e-7
+ trnqsmod = 0
+ petab = -7.719916e-16
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.00140826488
+ kt1 = 0.12069622
+ lk2 = -4.2131932e-9
+ kt2 = -0.11741295
+ wketa = 1.87190595e-7
+ llc = 0
+ lln = 1
+ lu0 = -5.407799999999904e-13
+ mjd = 0.26
+ lua = 1.6761980000000137e-18
+ mjs = 0.26
+ lub = 8.339062399999967e-27
+ luc = -2.98810456e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ tpbsw = 0.0019
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 9.065128000000001e-14
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ nsd = 1e+20
+ pbd = 0.52
+ pat = -2.5768428e-10
+ pbs = 0.52
+ pk2 = 5.9540883e-16
+ cjswd = 8.6592e-11
+ cjsws = 8.6592e-11
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ pu0 = -5.643113e-17
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ prt = 0
+ pua = -1.6092489999999997e-23
+ pub = 1.5276544400000003e-32
+ puc = 5.518326299999999e-24
+ pud = 0
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = -1.1935669e-9
+ ub1 = 2.1692222300000005e-18
+ uc1 = 8.622799700000001e-10
+ tpb = 0.0014
+ k2we = 5e-5
+ wa0 = -2.59429679e-6
+ tvfbsdoff = 0.022
+ ute = -1
+ wat = 0.0028451685
+ dsub = 0.75
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -1.1593839e-8
+ ltvoff = -1.1952424e-10
+ dtox = 2.7e-10
+ wlc = 0
+ wln = 1
+ rgatemod = 0
+ wu0 = 7.629837000000001e-10
+ xgl = -1.09e-8
+ xgw = 0
+ wua = 3.2583921000000013e-16
+ wub = -3.447615700000002e-25
+ wuc = -8.750290400000002e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ tnjtsswg = 1
+ )

.model nch_sf_33 nmos (
+ level = 54
+ rbodymod = 0
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ version = 4.5
+ pbswgd = 0.95
+ pbswgs = 0.95
+ ntox = 1.0
+ pcit = 1.2000000000000001e-17
+ pclm = 1.8851852
+ tempmod = 0
+ igcmod = 1
+ phin = 0.15
+ aigbacc = 0.02
+ pkt1 = -1.76e-16
+ wpdiblc2 = -2.9834e-10
+ pvoff = -4e-17
+ cdscb = 0
+ cdscd = 0
+ pvsat = 1.44e-11
+ aigbinv = 0.0163
+ rbdb = 50
+ prwb = 0
+ prwg = 0
+ pub1 = 1.6e-34
+ wk2we = 5e-12
+ pvth0 = 1.2e-16
+ drout = 0.56
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ rdsw = 100
+ permod = 1
+ voffl = 0
+ weta0 = 0
+ wkvth0we = 2e-12
+ cgidl = 0.22
+ trnqsmod = 0
+ voffcv = -0.16942
+ wpemod = 1
+ poxedge = 1
+ rshg = 15.6
+ binunit = 2
+ pbswd = 0.8
+ pbsws = 0.8
+ rgatemod = 0
+ tnjtsswg = 1
+ tnom = 25
+ pdits = 0
+ ags = 0.76882593
+ cigsd = 0.069865
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ tpbswg = 0.0009
+ cjd = 0.001432992
+ dvt0w = 0
+ cit = 0.002342713
+ dvt1w = 0
+ cjs = 0.001432992
+ clc = 1e-7
+ cle = 0.6
+ dvt2w = 0
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 9.8024918e-9
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ jtsswgd = 2.3e-7
+ pk2we = -1e-19
+ jtsswgs = 2.3e-7
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ la0 = 0
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = 8e-5
+ kt1 = -0.21767878
+ kt2 = -0.055117852
+ ptvoff = 0
+ llc = 0
+ lln = 1
+ lu0 = -4e-12
+ wags = 2.4994444e-8
+ mjd = 0.26
+ mjs = 0.26
+ lub = 0
+ lud = 0
+ lwc = 0
+ waigsd = 3.1789128e-12
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 0
+ tnoia = 0
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 1.44e-11
+ wcit = -2.9566928e-10
+ pbs = 0.52
+ pu0 = -1.2e-18
+ prt = 0
+ pub = 0
+ pud = 0
+ peta0 = 0.0
+ diomod = 1
+ voff = -0.095952978
+ acde = 0.4
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 9.5347726e-10
+ wketa = -1.1490089e-9
+ ub1 = -5.3850981e-19
+ uc1 = -6.0041111e-11
+ tpb = 0.0014
+ tpbsw = 0.0019
+ pditsd = 0
+ pditsl = 0
+ vsat = 84306.193
+ wa0 = 0
+ cjswgd = 2.9779200000000003e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.9779200000000003e-10
+ wint = 0
+ ute = -1
+ wat = 0
+ vth0 = 0.33989411
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 3.0219344e-9
+ cjswd = 8.6592e-11
+ cjsws = 8.6592e-11
+ wlc = 0
+ wln = 1
+ wu0 = 5.930666700000001e-11
+ wkt1 = 1.6685417500000003e-9
+ wkt2 = 1.0235511e-10
+ xgl = -1.09e-8
+ mjswd = 0.11
+ xgw = 0
+ mjsws = 0.11
+ wua = -1.6467997e-17
+ wub = 3.619626e-26
+ wuc = -1.4955111e-18
+ wud = 0
+ agidl = 9.41e-8
+ wmax = 2.726e-7
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ aigc = 0.01181895
+ wmin = 1.08e-7
+ tvfbsdoff = 0.022
+ njtsswg = 9
+ mjswgd = 0.85
+ mjswgs = 0.85
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ wua1 = -3.1223388e-18
+ wub1 = 2.0807554e-26
+ wuc1 = 8.1864667e-18
+ tcjswg = 0.001
+ bigc = 0.001442
+ ckappad = 0.6
+ ckappas = 0.6
+ wwlc = 0
+ pdiblc1 = 0
+ pdiblc2 = 0.023869018
+ pdiblcb = -0.3
+ scref = 1e-6
+ cdsc = 0
+ ijthsfwd = 0.01
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ pigcd = 2.621
+ aigsd = 0.010772573
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ lvoff = 1.6e-11
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ bigbacc = 0.002588
+ lvsat = 0.00016
+ lvth0 = 4.0000000000000007e-10
+ fprout = 300
+ ijthsrev = 0.01
+ delta = 0.007595625
+ xrcrg1 = 12
+ xrcrg2 = 1
+ kvth0we = 0.00018
+ rnoia = 0
+ rnoib = 0
+ lintnoi = -1.5e-8
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ wtvoff = 2.5061202e-10
+ ngate = 8e+20
+ wtvfbsdoff = 0
+ ngcon = 1
+ wpclm = -9.7111111e-9
+ k2we = 5e-5
+ dsub = 0.75
+ dtox = 2.7e-10
+ gbmin = 1e-12
+ capmod = 2
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ ltvfbsdoff = 0
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ wku0we = 2e-11
+ mobmod = 0
+ eta0 = 0.2
+ etab = -0.2
+ pkvth0we = -1.3e-19
+ nfactor = 1
+ ptvfbsdoff = 0
+ tvoff = 0.00085486634
+ vfbsdoff = 0.02
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ paramchk = 1
+ nigbacc = 10
+ ku0we = -0.0007
+ beta0 = 13
+ leta0 = -1.6000000000000003e-9
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ dlcig = 2.5e-9
+ nigbinv = 10
+ bgidl = 2320000000.0
+ ijthdfwd = 0.01
+ keta = -0.021050128
+ dmcgt = 0
+ tcjsw = 0.000357
+ toxref = 3e-9
+ ijthdrev = 0.01
+ fnoimod = 1
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 8e-12
+ eigbinv = 1.1
+ kt1l = 0
+ bigsd = 0.00125
+ lint = 6.5375218e-9
+ lkt1 = -2.4e-10
+ wvoff = 2.6481533e-9
+ lmax = 2.001e-5
+ lmin = 8.9991e-6
+ ltvoff = 0
+ lpe0 = 9.2e-8
+ wvsat = 0.002322956
+ lpeb = 2.5e-7
+ wvth0 = -1.1513739e-9
+ a0 = 3.5
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 200000
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.017556401
+ k3 = -1.8419
+ em = 1000000.0
+ minv = -0.3
+ waigc = 1.7818122e-11
+ ll = 0
+ lw = 0
+ u0 = 0.013255556000000002
+ w0 = 0
+ lub1 = 2.4000000000000004e-27
+ ua = -2.0911548e-9
+ ub = 2.2368542e-18
+ uc = 5.8018519e-11
+ ud = 0
+ cigbacc = 0.32875
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 3.4e-9
+ ndep = 1e+18
+ lkvth0we = -2e-12
+ pvfbsdoff = 0
+ lwlc = 0
+ moin = 5.1
+ lku0we = 2.5e-11
+ tnoimod = 0
+ epsrox = 3.9
+ xpart = 1
+ nigc = 3.083
+ cigbinv = 0.006
+ acnqsmod = 0
+ rdsmod = 0
+ egidl = 0.29734
+ igbmod = 1
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ )

.model nch_sf_34 nmos (
+ level = 54
+ paramchk = 1
+ wpclm = -9.7111111e-9
+ gbmin = 1e-12
+ wua1 = -1.7574281e-19
+ wub1 = 1.7597088e-26
+ wuc1 = 8.3134424e-18
+ jswgd = 1.28e-13
+ nfactor = 1
+ jswgs = 1.28e-13
+ paigsd = -3.8370159e-23
+ bigc = 0.001442
+ wwlc = 0
+ permod = 1
+ cdsc = 0
+ ijthdfwd = 0.01
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ nigbacc = 10
+ ijthdrev = 0.01
+ voffcv = -0.16942
+ wpemod = 1
+ tvoff = 0.00082419905
+ lpdiblc2 = -9.2950492e-9
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ nigbinv = 10
+ k2we = 5e-5
+ ku0we = -0.0007
+ beta0 = 13
+ dsub = 0.75
+ leta0 = -1.6000000000000003e-9
+ dtox = 2.7e-10
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ tpbswg = 0.0009
+ fnoimod = 1
+ lkvth0we = -2e-12
+ eigbinv = 1.1
+ dlcig = 2.5e-9
+ eta0 = 0.2
+ bgidl = 2320000000.0
+ etab = -0.2
+ acnqsmod = 0
+ ptvoff = -2.3727895e-16
+ waigsd = 3.1789171e-12
+ dmcgt = 0
+ tcjsw = 0.000357
+ rbodymod = 0
+ diomod = 1
+ cigbacc = 0.32875
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 2.9779200000000003e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.9779200000000003e-10
+ bigsd = 0.00125
+ tnoimod = 0
+ wvoff = 2.821381e-9
+ mjswgd = 0.85
+ mjswgs = 0.85
+ cigbinv = 0.006
+ wvsat = 0.002322956
+ wvth0 = -1.3363659000000004e-9
+ wpdiblc2 = -6.4961636e-10
+ tcjswg = 0.001
+ waigc = 1.8291238e-11
+ pvfbsdoff = 0
+ version = 4.5
+ lketa = -2.7750915e-8
+ tempmod = 0
+ xpart = 1
+ egidl = 0.29734
+ aigbacc = 0.02
+ keta = -0.017963263
+ wkvth0we = 2e-12
+ wtvfbsdoff = 0
+ fprout = 300
+ lags = 4.3821463e-7
+ xrcrg1 = 12
+ xrcrg2 = 1
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = -1.2651054999999995e-12
+ trnqsmod = 0
+ kt1l = 0
+ ltvfbsdoff = 0
+ aigbinv = 0.0163
+ wtvoff = 2.7700567e-10
+ lint = 6.5375218e-9
+ lkt1 = -8.905846799999999e-8
+ lkt2 = -1.6837724e-8
+ lmax = 8.9991e-6
+ lmin = 8.9908e-7
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ capmod = 2
+ rgatemod = 0
+ pvoff = -1.5973172e-15
+ tnjtsswg = 1
+ wku0we = 2e-11
+ minv = -0.3
+ lua1 = -7.4262143e-17
+ lub1 = -1.3918035e-25
+ luc1 = 6.2830403e-17
+ cdscb = 0
+ cdscd = 0
+ mobmod = 0
+ pvsat = 1.44e-11
+ ndep = 1e+18
+ wk2we = 5e-12
+ pvth0 = 1.7830782e-15
+ ptvfbsdoff = 0
+ drout = 0.56
+ lwlc = 0
+ poxedge = 1
+ moin = 5.1
+ paigc = -4.2533129e-18
+ nigc = 3.083
+ voffl = 0
+ binunit = 2
+ weta0 = 0
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ laigsd = 3.3658034e-16
+ pags = 5.2134206e-15
+ cgidl = 0.22
+ ntox = 1.0
+ pcit = 9.1881874e-17
+ pclm = 1.8851852
+ phin = 0.15
+ pbswd = 0.8
+ pbsws = 0.8
+ ags = 0.72008125
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ pkt1 = -5.4016964e-16
+ pkt2 = -1.7740443e-15
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ cjd = 0.001432992
+ cit = 0.0023437436
+ cjs = 0.001432992
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 9.8024918e-9
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ pdits = 0
+ cigsd = 0.069865
+ rbdb = 50
+ pua1 = -2.6489898e-23
+ prwb = 0
+ prwg = 0
+ pub1 = 2.902209e-32
+ puc1 = -1.1415122e-24
+ dvt0w = 0
+ la0 = -1.6207075e-6
+ dvt1w = 0
+ dvt2w = 0
+ rbpb = 50
+ rbpd = 50
+ jsd = 6.11e-7
+ rbps = 50
+ jss = 6.11e-7
+ lat = -0.043142769000000004
+ rbsb = 50
+ pvag = 1.2
+ kt1 = -0.20779908
+ lk2 = -1.5849432e-8
+ kt2 = -0.053244913
+ llc = 0
+ lln = 1
+ lu0 = -1.6832432e-9
+ mjd = 0.26
+ lua = -1.2813977e-16
+ mjs = 0.26
+ lub = -8.5009677e-26
+ luc = -2.2547224e-17
+ lud = 0
+ ijthsfwd = 0.01
+ lwc = 0
+ lwl = 0
+ rdsw = 100
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 3.8370159e-14
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 4.0048965e-9
+ pbs = 0.52
+ pk2 = -8.7965669e-16
+ pk2we = -1e-19
+ pu0 = -1.2000000000016282e-18
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ prt = 0
+ pua = -3.3674591e-24
+ pub = -4.9159389e-33
+ puc = 2.3789498e-24
+ pud = 0
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 9.6173779e-10
+ ub1 = -5.2276116e-19
+ uc1 = -6.7030033e-11
+ njtsswg = 9
+ tpb = 0.0014
+ toxref = 3e-9
+ wa0 = -4.2680933e-9
+ tnoia = 0
+ ute = -1
+ wat = -0.0004438817
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 3.1197827e-9
+ wlc = 0
+ wln = 1
+ wu0 = 5.930666700000001e-11
+ ijthsrev = 0.01
+ xgl = -1.09e-8
+ xtsswgd = 0.18
+ xgw = 0
+ xtsswgs = 0.18
+ wua = -1.6093419e-17
+ wub = 3.6743083e-26
+ wuc = -1.7601329e-18
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ peta0 = 0.0
+ wketa = -1.4921751e-9
+ ckappad = 0.6
+ ckappas = 0.6
+ rshg = 15.6
+ pdiblc1 = 0
+ pdiblc2 = 0.02490295
+ tpbsw = 0.0019
+ pdiblcb = -0.3
+ cjswd = 8.6592e-11
+ cjsws = 8.6592e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ tvfbsdoff = 0.022
+ ltvoff = 2.7569894e-10
+ ppdiblc2 = 3.1579745e-15
+ bigbacc = 0.002588
+ tnom = 25
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ kvth0we = 0.00018
+ lku0we = 2.5e-11
+ epsrox = 3.9
+ scref = 1e-6
+ lintnoi = -1.5e-8
+ pigcd = 2.621
+ bigbinv = 0.004953
+ aigsd = 0.010772573
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ rdsmod = 0
+ wvfbsdoff = 0
+ igbmod = 1
+ lvoff = -1.4722881e-8
+ lvfbsdoff = 0
+ pkvth0we = -1.3e-19
+ wags = 2.4414531000000003e-8
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ lvsat = 0.00016
+ wcit = -3.0455491e-10
+ lvth0 = 5.701542e-8
+ pbswgd = 0.95
+ pbswgs = 0.95
+ voff = -0.094313503
+ delta = 0.007595625
+ laigc = -1.6452737e-10
+ acde = 0.4
+ a0 = 3.6802789
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ vfbsdoff = 0.02
+ igcmod = 1
+ at = 204807.87
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.019319408
+ k3 = -1.8419
+ em = 1000000.0
+ rnoia = 0
+ rnoib = 0
+ ll = 0
+ lw = 0
+ vsat = 84306.193
+ u0 = 0.013442346
+ w0 = 0
+ wint = 0
+ ua = -2.0769012e-9
+ ub = 2.2463102e-18
+ uc = 6.0526552e-11
+ ud = 0
+ vth0 = 0.33359651
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 3.4e-9
+ wkt1 = 1.7090500500000002e-9
+ wkt2 = 2.996904e-10
+ wmax = 2.726e-7
+ aigc = 0.011837251
+ wmin = 1.08e-7
+ pketa = 3.0850638e-15
+ ngate = 8e+20
+ ngcon = 1
+ )

.model nch_sf_35 nmos (
+ level = 54
+ a0 = 2.7573663
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ voffl = 0
+ at = 225908.74
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.012837040000000001
+ k3 = -1.8419
+ em = 1000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.01303229
+ w0 = 0
+ ua = -2.2251639e-9
+ ub = 2.3450974e-18
+ uc = 3.6825844e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 3.4e-9
+ weta0 = 0
+ keta = -0.063873893
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ voffcv = -0.16942
+ wpemod = 1
+ lags = -4.2829945e-7
+ ijthsrev = 0.01
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ cgidl = 0.22
+ lcit = -6.1090204e-10
+ kt1l = 0
+ ags = 1.6936926
+ cjd = 0.001432992
+ cit = 0.0030287289
+ cjs = 0.001432992
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 9.8024918e-9
+ k3b = 1.9326
+ lint = 6.5375218e-9
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ lkt1 = 4.8811427e-8
+ lkt2 = -1.4519819e-8
+ pbswd = 0.8
+ pbsws = 0.8
+ lmax = 8.9908e-7
+ lmin = 4.4908e-7
+ lpe0 = 9.2e-8
+ la0 = -7.9931523e-7
+ lpeb = 2.5e-7
+ jsd = 6.11e-7
+ ppdiblc2 = -1.3141262e-15
+ jss = 6.11e-7
+ lat = -0.061922545
+ kt1 = -0.36270908
+ lk2 = -1.00801338e-8
+ kt2 = -0.0558493
+ llc = 0
+ lln = 1
+ lu0 = -1.3182934e-9
+ njtsswg = 9
+ mjd = 0.26
+ lua = 3.8140531e-18
+ mjs = 0.26
+ lub = -1.7293024e-25
+ luc = -1.4535934e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ tpbswg = 0.0009
+ njd = 1.02
+ minv = -0.3
+ njs = 1.02
+ pa0 = -6.7606598e-14
+ lua1 = -1.6437259e-16
+ lub1 = 2.5218043e-26
+ nsd = 1e+20
+ pdits = 0
+ luc1 = 5.6450349e-17
+ pbd = 0.52
+ pat = 1.7176657e-9
+ pbs = 0.52
+ pk2 = -9.651779000000002e-17
+ cigsd = 0.069865
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ pu0 = 7.7578742e-18
+ prt = 0
+ ndep = 1e+18
+ pua = -1.9061799e-24
+ pub = 1.3958464e-33
+ puc = -1.352132e-24
+ pud = 0
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ lwlc = 0
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 1.0629855e-9
+ ckappad = 0.6
+ ub1 = -7.0747845e-19
+ moin = 5.1
+ uc1 = -5.9861432e-11
+ ckappas = 0.6
+ tpb = 0.0014
+ pdiblc1 = 0
+ pdiblc2 = 0.01020022
+ pdiblcb = -0.3
+ wa0 = 1.1480691e-7
+ ute = -1
+ nigc = 3.083
+ wat = 0.0021260405
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 2.2398522999999998e-9
+ wlc = 0
+ pk2we = -1e-19
+ ptvoff = -4.8469984e-16
+ wln = 1
+ wu0 = 4.9241640000000006e-11
+ xgl = -1.09e-8
+ dvtp0 = 4e-7
+ xgw = 0
+ dvtp1 = 0.01
+ wua = -1.7735306e-17
+ wub = 2.9651178e-26
+ wuc = 2.4320938e-18
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ waigsd = 3.178874e-12
+ pkvth0we = -1.3e-19
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ tnoia = 0
+ diomod = 1
+ bigbacc = 0.002588
+ peta0 = 0.0
+ pags = -9.2425378e-15
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 2.9779200000000003e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.9779200000000003e-10
+ wketa = 5.5022601e-9
+ vfbsdoff = 0.02
+ ntox = 1.0
+ pcit = 1.708079e-16
+ pclm = 1.8851852
+ tpbsw = 0.0019
+ kvth0we = 0.00018
+ cjswd = 8.6592e-11
+ cjsws = 8.6592e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ phin = 0.15
+ tvfbsdoff = 0.022
+ lintnoi = -1.5e-8
+ bigbinv = 0.004953
+ mjswgd = 0.85
+ mjswgs = 0.85
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ paramchk = 1
+ pkt1 = -1.3387355e-14
+ pkt2 = 1.7857928e-15
+ tcjswg = 0.001
+ wtvfbsdoff = 0
+ rbdb = 50
+ pua1 = 3.1539092e-23
+ prwb = 0
+ prwg = 0
+ pub1 = -3.1373886e-32
+ puc1 = -7.798421e-24
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ scref = 1e-6
+ ijthdfwd = 0.01
+ rdsw = 100
+ pigcd = 2.621
+ aigsd = 0.010772573
+ ltvfbsdoff = 0
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ lvoff = -2.8440354e-8
+ fprout = 300
+ lvsat = 0.00016
+ xrcrg1 = 12
+ xrcrg2 = 1
+ lvth0 = 1.9154806e-8
+ ijthdrev = 0.01
+ delta = 0.007595625
+ nfactor = 1
+ laigc = -6.1235169e-11
+ lpdiblc2 = 3.7903799e-9
+ rshg = 15.6
+ rnoia = 0
+ rnoib = 0
+ wtvoff = 5.5500668e-10
+ ptvfbsdoff = 0
+ pketa = -3.1399835e-15
+ ngate = 8e+20
+ ngcon = 1
+ wpclm = -9.7111111e-9
+ capmod = 2
+ wku0we = 2e-11
+ gbmin = 1e-12
+ nigbacc = 10
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ mobmod = 0
+ tnom = 25
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ lkvth0we = -2e-12
+ nigbinv = 10
+ acnqsmod = 0
+ wags = 4.0657181e-8
+ rbodymod = 0
+ wcit = -3.9323584e-10
+ voff = -0.078900611
+ tvoff = -3.4914836e-5
+ acde = 0.4
+ fnoimod = 1
+ xjbvd = 1
+ xjbvs = 1
+ vsat = 84306.193
+ lk2we = -1.5e-12
+ eigbinv = 1.1
+ wint = 0
+ vth0 = 0.37613652
+ wkt1 = 1.614409e-8
+ wkt2 = -3.7001265e-9
+ wmax = 2.726e-7
+ aigc = 0.011721192
+ wmin = 1.08e-7
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ ku0we = -0.0007
+ beta0 = 13
+ leta0 = -1.6000000000000003e-9
+ wpdiblc2 = 4.3752159e-9
+ wua1 = -6.5376855e-17
+ wub1 = 8.5457734e-26
+ wuc1 = 1.5793115e-17
+ bigc = 0.001442
+ wwlc = 0
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ cigbacc = 0.32875
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ tnoimod = 0
+ cigc = 0.000625
+ toxref = 3e-9
+ dmcgt = 0
+ tcjsw = 0.000357
+ wkvth0we = 2e-12
+ cigbinv = 0.006
+ trnqsmod = 0
+ bigsd = 0.00125
+ version = 4.5
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ tempmod = 0
+ ltvoff = 1.0403103e-9
+ wvoff = -2.4321636000000003e-9
+ k2we = 5e-5
+ wvsat = 0.002322956
+ aigbacc = 0.02
+ dsub = 0.75
+ wvth0 = 2.1985258999999998e-9
+ dtox = 2.7e-10
+ rgatemod = 0
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ tnjtsswg = 1
+ waigc = 1.00872e-11
+ pvfbsdoff = 0
+ lku0we = 2.5e-11
+ epsrox = 3.9
+ eta0 = 0.2
+ etab = -0.2
+ lketa = 1.3109546e-8
+ aigbinv = 0.0163
+ xpart = 1
+ rdsmod = 0
+ igbmod = 1
+ egidl = 0.29734
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ pbswgd = 0.95
+ pbswgs = 0.95
+ igcmod = 1
+ poxedge = 1
+ binunit = 2
+ pvoff = 3.0783375000000003e-15
+ cdscb = 0
+ cdscd = 0
+ pvsat = 1.44e-11
+ wk2we = 5e-12
+ pvth0 = -1.3629756000000001e-15
+ drout = 0.56
+ permod = 1
+ paigc = 3.0482801e-18
+ ijthsfwd = 0.01
+ )

.model nch_sf_36 nmos (
+ level = 54
+ rshg = 15.6
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ cigbacc = 0.32875
+ tnoimod = 0
+ ku0we = -0.0007
+ a0 = 2.8517872
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ beta0 = 13
+ at = 72186.119
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.0046985251
+ k3 = -1.8419
+ em = 1000000.0
+ leta0 = -1.6000000000000003e-9
+ rgatemod = 0
+ ll = -1.18e-13
+ lw = 0
+ u0 = 0.011248434000000002
+ tpbswg = 0.0009
+ w0 = 0
+ ua = -2.2247872e-9
+ ub = 2.0937783e-18
+ uc = 7.1203963e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ tnjtsswg = 1
+ ww = 0
+ xw = 3.4e-9
+ cigbinv = 0.006
+ tnom = 25
+ ppclm = 2.75592e-14
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ ptvoff = 2.8225911e-16
+ version = 4.5
+ waigsd = 3.178874e-12
+ tempmod = 0
+ dmcgt = 0
+ tcjsw = 0.000357
+ diomod = 1
+ wags = 2.5408180000000003e-7
+ aigbacc = 0.02
+ wcit = 1.4683634000000001e-10
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 2.9779200000000003e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.9779200000000003e-10
+ voff = -0.13810998
+ acde = 0.4
+ bigsd = 0.00125
+ vsat = 84306.193
+ wint = 0
+ vth0 = 0.43875442
+ wtvfbsdoff = 0
+ wkt1 = -3.6010623e-8
+ wkt2 = -4.3121065e-11
+ aigbinv = 0.0163
+ wmax = 2.726e-7
+ mjswgd = 0.85
+ mjswgs = 0.85
+ aigc = 0.011581706
+ wmin = 1.08e-7
+ wvoff = 6.8440927000000005e-9
+ tcjswg = 0.001
+ wvsat = 0.002322956
+ ltvfbsdoff = 0
+ wvth0 = -3.5496131000000003e-9
+ wua1 = 2.3276683e-17
+ wub1 = 1.5603072e-26
+ wuc1 = -5.1034561e-18
+ waigc = 2.6093343e-11
+ pvfbsdoff = 0
+ bigc = 0.001442
+ wwlc = 0
+ lketa = -3.8407777e-8
+ ijthsfwd = 0.01
+ cdsc = 0
+ xpart = 1
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ poxedge = 1
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ egidl = 0.29734
+ fprout = 300
+ ptvfbsdoff = 0
+ binunit = 2
+ xrcrg1 = 12
+ xrcrg2 = 1
+ ijthsrev = 0.01
+ wtvoff = -1.1880818e-9
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ capmod = 2
+ k2we = 5e-5
+ wku0we = 2e-11
+ ppdiblc2 = 3.3310302e-16
+ dsub = 0.75
+ dtox = 2.7e-10
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ pvoff = -1.00321526e-15
+ mobmod = 0
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ cdscb = 0
+ cdscd = 0
+ pvsat = 1.44e-11
+ wk2we = 5e-12
+ pvth0 = 1.1662056e-15
+ drout = 0.56
+ eta0 = 0.2
+ etab = -0.2
+ paigc = -3.9944226e-18
+ voffl = 0
+ weta0 = 0
+ pkvth0we = -1.3e-19
+ ags = -2.4947885
+ lpclm = -2.4174737e-7
+ cjd = 0.001432992
+ cit = 0.00083484714
+ cjs = 0.001432992
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 1.30529375e-8
+ k3b = 1.9326
+ njtsswg = 9
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ cgidl = 0.22
+ vfbsdoff = 0.02
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ la0 = -8.4086042e-7
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = 0.0057154098000000006
+ kt1 = -0.088256509
+ lk2 = -6.4991688e-9
+ kt2 = -0.075738087
+ ckappad = 0.6
+ ckappas = 0.6
+ llc = -1.18e-13
+ lln = 0.7
+ lu0 = -5.3339671e-10
+ mjd = 0.26
+ pdiblc1 = 0
+ pdiblc2 = 0.031716534
+ lua = 3.6483177e-18
+ mjs = 0.26
+ lub = -6.2349821e-26
+ luc = -1.6579966e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ pdiblcb = -0.3
+ njd = 1.02
+ njs = 1.02
+ pa0 = 8.661463e-14
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ pbswd = 0.8
+ pbsws = 0.8
+ nsd = 1e+20
+ pbd = 0.52
+ pat = -3.1274679000000003e-9
+ pbs = 0.52
+ pk2 = -2.9168571e-16
+ paramchk = 1
+ pu0 = 1.2409578e-18
+ prt = 0
+ pua = -4.9144669e-25
+ pub = 1.8790045e-33
+ puc = 1.8346553e-24
+ pud = 0
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 5.8363721e-10
+ ub1 = -5.3348382e-19
+ uc1 = 8.6067289e-11
+ tpb = 0.0014
+ wa0 = -2.3569588e-7
+ ute = -1
+ wat = 0.013137708
+ pdits = 0
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 2.6834067999999997e-9
+ wlc = 0
+ wln = 1
+ cigsd = 0.069865
+ wu0 = 6.4052813e-11
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -2.0950609e-17
+ wub = 2.8553091e-26
+ wuc = -4.8106046e-18
+ wud = 0
+ wwc = 0
+ bigbacc = 0.002588
+ wwl = 0
+ wwn = 1
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ ijthdfwd = 0.01
+ kvth0we = 0.00018
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ toxref = 3e-9
+ lintnoi = -1.5e-8
+ keta = 0.053210932
+ bigbinv = 0.004953
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ tnoia = 0
+ lags = 1.4146322e-6
+ ijthdrev = 0.01
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ peta0 = 0.0
+ lcit = 3.5440592000000004e-10
+ wketa = -7.2433388e-9
+ kt1l = 0
+ lpdiblc2 = -5.676798e-9
+ tpbsw = 0.0019
+ cjswd = 8.6592e-11
+ cjsws = 8.6592e-11
+ mjswd = 0.11
+ tvfbsdoff = 0.022
+ mjsws = 0.11
+ ltvoff = -1.663256e-9
+ agidl = 9.41e-8
+ lint = 9.7879675e-9
+ lkt1 = -7.1947703e-8
+ lkt2 = -5.7687528e-9
+ lmax = 4.4908e-7
+ lmin = 2.1577e-7
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ minv = -0.3
+ lku0we = 2.5e-11
+ lua1 = 4.6540649e-17
+ lub1 = -5.1339597e-26
+ luc1 = -7.7582888e-18
+ epsrox = 3.9
+ lkvth0we = -2e-12
+ ndep = 1e+18
+ nfactor = 1
+ lwlc = 0
+ moin = 5.1
+ scref = 1e-6
+ rdsmod = 0
+ pigcd = 2.621
+ nigc = 3.083
+ igbmod = 1
+ aigsd = 0.010772573
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ acnqsmod = 0
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ lvoff = -2.3882325e-9
+ pbswgd = 0.95
+ noff = 2.7195
+ pbswgs = 0.95
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ lvsat = 0.00016
+ rbodymod = 0
+ lvth0 = -8.3970687e-9
+ igcmod = 1
+ nigbacc = 10
+ delta = 0.007595625
+ pags = -1.0314937e-13
+ laigc = 1.3898222e-13
+ ntox = 1.0
+ pcit = -6.682386e-17
+ pclm = 2.434611
+ rnoia = 0
+ rnoib = 0
+ phin = 0.15
+ pketa = 2.46808e-15
+ ngate = 8e+20
+ nigbinv = 10
+ ngcon = 1
+ wpclm = -7.2345657e-8
+ pkt1 = 9.5607187e-15
+ pkt2 = 1.7671038e-16
+ wpdiblc2 = 6.3151306e-10
+ gbmin = 1e-12
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ permod = 1
+ rbdb = 50
+ pua1 = -7.4684646e-24
+ prwb = 0
+ prwg = 0
+ pub1 = -6.378346e-34
+ puc1 = 1.3960704e-24
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ fnoimod = 1
+ rdsw = 100
+ eigbinv = 1.1
+ wkvth0we = 2e-12
+ voffcv = -0.16942
+ wpemod = 1
+ trnqsmod = 0
+ tvoff = 0.006109554
+ )

.model nch_sf_37 nmos (
+ level = 54
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ pdits = 0
+ cigsd = 0.069865
+ lkvth0we = -2e-12
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ eta0 = 0.2
+ etab = -0.2
+ ptvoff = -1.8615536e-17
+ waigsd = 3.178874e-12
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ acnqsmod = 0
+ diomod = 1
+ wtvfbsdoff = 0
+ tnoia = 0
+ pditsd = 0
+ pditsl = 0
+ rbodymod = 0
+ cjswgd = 2.9779200000000003e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.9779200000000003e-10
+ a0 = -2.4455841
+ a1 = 0
+ a2 = 1
+ peta0 = 0.0
+ b0 = 0
+ b1 = 0
+ ltvfbsdoff = 0
+ at = 121458.51
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = -0.003797302
+ k3 = -1.8419
+ em = 1000000.0
+ ll = -1.18e-13
+ wketa = 1.2169685000000001e-8
+ lw = 0
+ u0 = 0.009644213
+ w0 = 0
+ ua = -2.2679307e-9
+ ub = 1.903479518e-18
+ uc = 2.5998306e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 3.4e-9
+ tpbsw = 0.0019
+ nfactor = 1
+ tvfbsdoff = 0.022
+ cjswd = 8.6592e-11
+ cjsws = 8.6592e-11
+ mjswgd = 0.85
+ mjswd = 0.11
+ mjswgs = 0.85
+ mjsws = 0.11
+ agidl = 9.41e-8
+ tcjswg = 0.001
+ wpdiblc2 = 2.0871493e-9
+ ptvfbsdoff = 0
+ nigbacc = 10
+ scref = 1e-6
+ wvfbsdoff = 0
+ pigcd = 2.621
+ lvfbsdoff = 0
+ aigsd = 0.010772573
+ fprout = 300
+ lvoff = 8.051419999999985e-11
+ nigbinv = 10
+ keta = -0.10792277
+ xrcrg1 = 12
+ xrcrg2 = 1
+ wkvth0we = 2e-12
+ lvsat = -0.00022927429499999992
+ lvth0 = -7.461937700000001e-9
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ trnqsmod = 0
+ delta = 0.007595625
+ lcit = -3.1333293000000004e-11
+ wtvoff = 2.3786433e-10
+ laigc = -6.7426314e-12
+ kt1l = 0
+ rnoia = 0
+ rnoib = 0
+ fnoimod = 1
+ lint = 9.7879675e-9
+ pketa = -1.6280779999999998e-15
+ ngate = 8e+20
+ capmod = 2
+ eigbinv = 1.1
+ lkt1 = 3.1879381e-10
+ lkt2 = 1.6714521e-10
+ lmax = 2.1577e-7
+ ngcon = 1
+ lmin = 9e-8
+ wpclm = 1.5314007e-7
+ wku0we = 2e-11
+ lpe0 = 9.2e-8
+ lpeb = 2.5e-7
+ mobmod = 0
+ rgatemod = 0
+ gbmin = 1e-12
+ tnjtsswg = 1
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ minv = -0.3
+ lua1 = -6.7367772e-18
+ lub1 = -3.5961216e-26
+ luc1 = -1.0970607e-17
+ ndep = 1e+18
+ lwlc = 0
+ moin = 5.1
+ nigc = 3.083
+ cigbacc = 0.32875
+ tnoimod = 0
+ noff = 2.7195
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ cigbinv = 0.006
+ tvoff = -0.0028392003
+ ntox = 1.0
+ pcit = 2.6940572e-17
+ pclm = 1.0592301
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ phin = 0.15
+ version = 4.5
+ tempmod = 0
+ pkt1 = -3.6229533e-16
+ pkt2 = -2.0087744e-16
+ ku0we = -0.0007
+ beta0 = 13
+ leta0 = -1.6000000000000003e-9
+ ppclm = -2.0018289e-14
+ aigbacc = 0.02
+ rbdb = 50
+ pua1 = 2.2068447e-24
+ prwb = 0
+ prwg = 0
+ pub1 = -2.5826774e-33
+ puc1 = 1.8773731e-24
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ ijthsfwd = 0.01
+ rdsw = 100
+ toxref = 3e-9
+ aigbinv = 0.0163
+ dmcgt = 0
+ tcjsw = 0.000357
+ ijthsrev = 0.01
+ rshg = 15.6
+ bigsd = 0.00125
+ ltvoff = 2.2493116e-10
+ wvoff = 1.4856166000000002e-9
+ poxedge = 1
+ wvsat = 0.00180338308
+ ppdiblc2 = 2.596377e-17
+ wvth0 = 2.1151897e-9
+ binunit = 2
+ pvfbsdoff = 0
+ lku0we = 2.5e-11
+ waigc = 5.3999849e-12
+ tnom = 25
+ epsrox = 3.9
+ toxe = 2.43e-9
+ toxm = 2.43e-9
+ rdsmod = 0
+ lketa = -4.408530899999999e-9
+ igbmod = 1
+ xpart = 1
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ egidl = 0.29734
+ pbswgd = 0.95
+ pbswgs = 0.95
+ pkvth0we = -1.3e-19
+ wags = -2.3477778e-7
+ igcmod = 1
+ wcit = -2.9754486000000003e-10
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ voff = -0.149810363
+ acde = 0.4
+ vfbsdoff = 0.02
+ vsat = 86151.12359999999
+ wint = 0
+ vth0 = 0.434322633
+ wkt1 = 1.10178791e-8
+ wkt2 = 1.7463947e-9
+ wmax = 2.726e-7
+ aigc = 0.01161432
+ wmin = 1.08e-7
+ paramchk = 1
+ pvoff = 1.2741821999999993e-16
+ wua1 = -2.2577864e-17
+ wub1 = 2.4820337e-26
+ wuc1 = -7.3845115e-18
+ cdscb = 0
+ cdscd = 0
+ bigc = 0.001442
+ permod = 1
+ pvsat = 1.2403312000000008e-10
+ wwlc = 0
+ njtsswg = 9
+ wk2we = 5e-12
+ pvth0 = -2.906062000000001e-17
+ drout = 0.56
+ ags = 4.2096296
+ paigc = 3.7187593e-19
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ ijthdfwd = 0.01
+ cdsc = 0
+ cjd = 0.001432992
+ cit = 0.0026629951
+ cgbo = 0
+ cjs = 0.001432992
+ clc = 1e-7
+ cle = 0.6
+ voffl = 0
+ cgdl = 3.31989e-12
+ bvd = 8.7
+ cgdo = 4.90562e-11
+ xtid = 3
+ bvs = 8.7
+ xtis = 3
+ dlc = 1.30529375e-8
+ ckappad = 0.6
+ ckappas = 0.6
+ k3b = 1.9326
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ cigc = 0.000625
+ pdiblc1 = 0
+ pdiblc2 = 0.0095469071
+ pdiblcb = -0.3
+ weta0 = 0
+ voffcv = -0.16942
+ wpemod = 1
+ lpclm = 4.8457997e-8
+ la0 = 2.768849e-7
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.0046810641
+ kt1 = -0.43075175
+ lk2 = -4.7065454e-9
+ kt2 = -0.10387031
+ ijthdrev = 0.01
+ llc = -1.18e-13
+ lln = 0.7
+ lu0 = -1.9490617e-10
+ mjd = 0.26
+ mjs = 0.26
+ lua = 1.2751594e-17
+ lub = -2.21968369e-26
+ cgidl = 0.22
+ luc = -7.0415723e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = -2.9632335e-14
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 5.169644e-10
+ pbs = 0.52
+ pk2 = 3.1759465e-16
+ lpdiblc2 = -9.9900678e-10
+ pu0 = -7.7197738e-19
+ bigbacc = 0.002588
+ prt = 0
+ pua = 3.9870432e-24
+ pub = -6.31495433e-33
+ puc = 2.2635812e-25
+ pud = 0
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 8.3613685e-10
+ ub1 = -6.0636714e-19
+ uc1 = 1.0129155e-10
+ tpb = 0.0014
+ wa0 = 3.1523761e-7
+ kvth0we = 0.00018
+ pbswd = 0.8
+ pbsws = 0.8
+ ute = -1
+ wat = -0.0041344832
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -2.0418175e-10
+ wlc = 0
+ wln = 1
+ wu0 = 7.359279e-11
+ xgl = -1.09e-8
+ xgw = 0
+ wua = -4.2175679e-17
+ wub = 6.73870221e-26
+ wuc = 2.8116572e-18
+ wud = 0
+ k2we = 5e-5
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ lintnoi = -1.5e-8
+ tpbswg = 0.0009
+ dsub = 0.75
+ bigbinv = 0.004953
+ dtox = 2.7e-10
+ vtsswgd = 4.2
+ vtsswgs = 4.2
+ )

.model nch_sf_38 nmos (
+ level = 54
+ dmcgt = 0
+ poxedge = 1
+ pkvth0we = -1.3e-19
+ tcjsw = 0.000357
+ pditsd = 0
+ pditsl = 0
+ noff = 2.7195
+ cjswgd = 2.9779200000000003e-10
+ pku0we = -1.5e-18
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ cjswgs = 2.9779200000000003e-10
+ binunit = 2
+ vfbsdoff = 0.02
+ ntox = 1.0
+ pcit = 1.07254761e-17
+ pclm = 2.2357699
+ bigsd = 0.00125
+ ptvfbsdoff = 0
+ mjswgd = 0.85
+ mjswgs = 0.85
+ tcjswg = 0.001
+ phin = 0.15
+ wvoff = 4.554463324000001e-9
+ paramchk = 1
+ pkt1 = -2.6265624e-15
+ pkt2 = 3.9546557e-16
+ wvsat = 0.0013518940999999985
+ wvth0 = 4.419156600000002e-9
+ pvfbsdoff = 0
+ waigc = -1.2918923e-11
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ rbdb = 50
+ pua1 = -4.7371604e-25
+ prwb = 0
+ pub1 = 5.4790487999999994e-33
+ prwg = 0
+ puc1 = -4.218097e-24
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 1.2
+ lketa = 3.7750018e-8
+ a0 = 0.7744856
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ ijthdfwd = 0.01
+ at = 111412.77840000001
+ cf = 8.15e-11
+ xpart = 1
+ ef = 1.0
+ k1 = 0.274
+ k2 = -0.041738197000000005
+ k3 = -1.8419
+ em = 1000000.0
+ rdsw = 100
+ ll = 0
+ lw = 0
+ u0 = 0.0054412099
+ w0 = 0
+ ua = -2.6695158e-9
+ ub = 2.0926996330000003e-18
+ uc = -9.6044814e-11
+ ud = 0
+ fprout = 300
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 3.4e-9
+ xrcrg1 = 12
+ xrcrg2 = 1
+ egidl = 0.29734
+ ijthdrev = 0.01
+ wtvoff = 2.7545299e-10
+ lpdiblc2 = 4.9724259e-14
+ rshg = 15.6
+ njtsswg = 9
+ capmod = 2
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ wku0we = 2e-11
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = -0.0010813536
+ mobmod = 0
+ pdiblcb = -0.3
+ ags = 4.2096296
+ pvoff = -1.610533700000001e-16
+ cjd = 0.001432992
+ cit = 0.001090691
+ cjs = 0.001432992
+ clc = 1e-7
+ cle = 0.6
+ cdscb = 0
+ cdscd = 0
+ bvd = 8.7
+ tnom = 25
+ bvs = 8.7
+ dlc = 3.26497e-9
+ pvsat = 1.664725e-10
+ k3b = 1.9326
+ lkvth0we = -2e-12
+ wk2we = 5e-12
+ toxe = 2.43e-9
+ dwb = 0
+ dwc = 0
+ toxm = 2.43e-9
+ dwg = 0
+ dwj = 0
+ pvth0 = -2.4563349999999997e-16
+ drout = 0.56
+ paigc = 2.0938533e-18
+ bigbacc = 0.002588
+ la0 = -2.5801646e-8
+ voffl = 0
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.00373676425
+ kt1 = -0.62571779
+ kt2 = -0.068117715
+ lk2 = -1.1401013e-9
+ llc = 0
+ lln = 1
+ lu0 = 2.0017611999999998e-10
+ mjd = 0.26
+ acnqsmod = 0
+ mjs = 0.26
+ lua = 5.0500592e-17
+ lub = -3.9983527e-26
+ luc = 4.4304811e-18
+ lud = 0
+ laigsd = 1.06572e-17
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ kvth0we = 0.00018
+ weta0 = 4.2794074e-8
+ pa0 = 2.9413877e-15
+ wetab = -1.5859302e-8
+ nsd = 1e+20
+ pbd = 0.52
+ pat = 7.9459749e-10
+ pbs = 0.52
+ pk2 = 2.316472e-16
+ lpclm = -6.2136744e-8
+ pu0 = -4.1481775e-17
+ wags = -2.3477778e-7
+ prt = 0
+ pua = -3.0159915e-24
+ pub = 1.3943639e-33
+ puc = 2.394639e-25
+ pud = 0
+ lintnoi = -1.5e-8
+ rbodymod = 0
+ wcit = -1.25043837e-10
+ bigbinv = 0.004953
+ rsh = 17.5
+ tcj = 0.00076
+ ua1 = 7.2026227e-10
+ vtsswgd = 4.2
+ ub1 = -6.033332e-19
+ vtsswgs = 4.2
+ uc1 = -2.7209866e-10
+ cgidl = 0.22
+ tpb = 0.0014
+ wa0 = -3.1291358e-8
+ voff = -0.11849200800000002
+ ute = -1
+ wat = -0.00708802596
+ acde = 0.4
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 7.1015279e-10
+ wlc = 0
+ wln = 1
+ wu0 = 5.0667574e-10
+ xgl = -1.09e-8
+ xgw = 0
+ wua = 3.2324691e-17
+ wub = -1.4627000299999995e-26
+ wuc = 2.6722336e-18
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ vsat = 69045.23300000001
+ wint = 0
+ vth0 = 0.29573340800000003
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ wkt1 = 3.5105826e-8
+ wkt2 = -4.5976799e-9
+ wmax = 2.726e-7
+ aigc = 0.011905208
+ wmin = 1.08e-7
+ pbswd = 0.8
+ pbsws = 0.8
+ wpdiblc2 = 2.3634934e-9
+ wua1 = 5.9387403e-18
+ wub1 = -6.0942626e-26
+ wuc1 = 5.7460914e-17
+ pdits = 0
+ bigc = 0.001442
+ cigsd = 0.069865
+ wwlc = 0
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ cdsc = 0
+ nfactor = 1
+ toxref = 3e-9
+ cgbo = 0
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ pk2we = -1e-19
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ wkvth0we = 2e-12
+ tnoia = 0
+ peta0 = -4.0226429e-15
+ trnqsmod = 0
+ petab = 1.4907744e-15
+ wketa = 2.4101615e-8
+ tpbsw = 0.0019
+ ltvoff = 1.3417313e-10
+ nigbacc = 10
+ tvfbsdoff = 0.022
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ cjswd = 8.6592e-11
+ cjsws = 8.6592e-11
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ k2we = 5e-5
+ nigbinv = 10
+ dsub = 0.75
+ rgatemod = 0
+ lku0we = 2.5e-11
+ dtox = 2.7e-10
+ tnjtsswg = 1
+ epsrox = 3.9
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ rdsmod = 0
+ eta0 = -0.13238438
+ etab = 0.18670848
+ igbmod = 1
+ scref = 1e-6
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ pigcd = 2.621
+ aigsd = 0.010772573
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ fnoimod = 1
+ pbswgd = 0.95
+ pbswgs = 0.95
+ eigbinv = 1.1
+ lvoff = -2.8634111999999997e-9
+ igcmod = 1
+ lvsat = 0.00137867915
+ lvth0 = 5.5654495e-9
+ delta = 0.007595625
+ laigc = -3.4086068e-11
+ rnoia = 0
+ rnoib = 0
+ pketa = -2.74968201e-15
+ ngate = 8e+20
+ paigsd = -2.9413875e-24
+ ngcon = 1
+ cigbacc = 0.32875
+ wpclm = -8.3073835e-8
+ gbmin = 1e-12
+ tnoimod = 0
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ permod = 1
+ cigbinv = 0.006
+ ijthsfwd = 0.01
+ voffcv = -0.16942
+ wpemod = 1
+ version = 4.5
+ keta = -0.55641828
+ tempmod = 0
+ ijthsrev = 0.01
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 1.164633e-10
+ tvoff = -0.0018736893
+ aigbacc = 0.02
+ kt1l = 0
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ lint = 0
+ lkt1 = 1.8645602e-8
+ lkt2 = -3.1935983e-9
+ lmax = 9e-8
+ lmin = 5.4e-8
+ tpbswg = 0.0009
+ ku0we = -0.0007
+ aigbinv = 0.0163
+ beta0 = 13
+ lpe0 = 9.2e-8
+ ppdiblc2 = -1.2574432e-20
+ lpeb = 2.5e-7
+ leta0 = 2.9644132e-8
+ letab = -3.6350598e-8
+ wtvfbsdoff = 0
+ minv = -0.3
+ ppclm = 2.1858187e-15
+ lua1 = 4.1554342e-18
+ lub1 = -3.6246403e-26
+ luc1 = 2.4128073e-17
+ ndep = 1e+18
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ ptvoff = -2.2148869e-17
+ lwlc = 0
+ moin = 5.1
+ ltvfbsdoff = 0
+ waigsd = 3.1789053e-12
+ nigc = 3.083
+ diomod = 1
+ )

.model nch_sf_39 nmos (
+ level = 54
+ wkt1 = 8.520945e-9
+ wkt2 = 1.1625249e-8
+ wmax = 2.726e-7
+ aigc = 0.011615807
+ wmin = 1.08e-7
+ fnoimod = 1
+ eigbinv = 1.1
+ wua1 = -1.0774777e-16
+ wub1 = 2.3670019e-25
+ wuc1 = 1.606153e-17
+ bigc = 0.001442
+ wwlc = 0
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ scref = 1e-6
+ ijthsfwd = 0.01
+ cdsc = 0
+ fprout = 300
+ pigcd = 2.621
+ cgbo = 0
+ aigsd = 0.010772573
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ xrcrg1 = 12
+ xrcrg2 = 1
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ lvoff = -6.472439900000001e-9
+ cigbacc = 0.32875
+ lvsat = -0.0009854400999999998
+ wtvoff = 7.91509e-11
+ lvth0 = 8.3107327e-9
+ ijthsrev = 0.01
+ tnoimod = 0
+ delta = 0.007595625
+ laigc = -1.730084e-11
+ rnoia = 0
+ rnoib = 0
+ cigbinv = 0.006
+ dmcg = 3.1e-8
+ capmod = 2
+ dmci = 3.1e-8
+ dmdg = 0
+ wku0we = 2e-11
+ pketa = 4.904375999999999e-15
+ ngate = 8e+20
+ a0 = 19.191807
+ a1 = 0
+ a2 = 1
+ ngcon = 1
+ b0 = 0
+ b1 = 0
+ mobmod = 0
+ wpclm = -5.2664346e-8
+ at = 96903.002
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = -0.056113829000000004
+ k3 = -1.8419
+ em = 1000000.0
+ k2we = 5e-5
+ ll = 0
+ lw = 0
+ u0 = 0.0024707365
+ w0 = 0
+ ua = -2.3710013e-9
+ ub = 1.4550579529999998e-18
+ uc = -1.4785261e-10
+ ud = 0
+ version = 4.5
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 3.4e-9
+ dsub = 0.75
+ dtox = 2.7e-10
+ gbmin = 1e-12
+ tempmod = 0
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ eta0 = 1.1504337
+ aigbacc = 0.02
+ etab = -1.3364008
+ pkvth0we = -1.3e-19
+ aigbinv = 0.0163
+ tvoff = -0.0045522389
+ vfbsdoff = 0.02
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ paramchk = 1
+ ku0we = -0.0007
+ beta0 = 13
+ leta0 = -4.4759315e-8
+ poxedge = 1
+ letab = 5.198974e-8
+ ppclm = 4.2206835e-16
+ binunit = 2
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ ijthdfwd = 0.01
+ toxref = 3e-9
+ dmcgt = 0
+ keta = 0.43329502999999997
+ tcjsw = 0.000357
+ ijthdrev = 0.01
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 4.6979023e-10
+ ltvoff = 2.8952901e-10
+ kt1l = 0
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ bigsd = 0.00125
+ lint = 0
+ wvoff = -2.548824599999999e-9
+ lkt1 = 1.0173925000000002e-8
+ lkt2 = 8.1983323e-9
+ lmax = 5.4e-8
+ lmin = 4.5e-8
+ wvsat = 0.002929912199999998
+ lku0we = 2.5e-11
+ pvfbsdoff = 0
+ lpe0 = 9.2e-8
+ wvth0 = -7.224421000000017e-10
+ lpeb = 2.5e-7
+ epsrox = 3.9
+ waigc = 4.0939876e-11
+ minv = -0.3
+ lua1 = -3.9796071e-17
+ lub1 = 6.2484051e-26
+ luc1 = 1.4911728e-19
+ rdsmod = 0
+ lkvth0we = -2e-12
+ ndep = 1e+18
+ igbmod = 1
+ lwlc = 0
+ lketa = -1.96532807e-8
+ moin = 5.1
+ njtsswg = 9
+ xpart = 1
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ nigc = 3.083
+ pbswgd = 0.95
+ pbswgs = 0.95
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ acnqsmod = 0
+ egidl = 0.29734
+ igcmod = 1
+ ckappad = 0.6
+ ckappas = 0.6
+ noff = 2.7195
+ pdiblc1 = 0
+ pdiblc2 = -0.0010804963
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ pdiblcb = -0.3
+ rbodymod = 0
+ ntox = 1.0
+ pcit = -9.822646999999999e-18
+ pclm = 1.0542662
+ ags = 4.2096296
+ bigbacc = 0.002588
+ phin = 0.15
+ cjd = 0.001432992
+ cit = -0.0050011527
+ cjs = 0.001432992
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 3.26497e-9
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ pkt1 = -1.08463924e-15
+ pkt2 = -5.454643e-16
+ dwg = 0
+ dwj = 0
+ kvth0we = 0.00018
+ wpdiblc2 = 2.3632766e-9
+ permod = 1
+ pvoff = 2.5093735e-16
+ lintnoi = -1.5e-8
+ la0 = -1.0940063e-6
+ cdscb = 0
+ cdscd = 0
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.00289519958
+ bigbinv = 0.004953
+ kt1 = -0.47965441
+ kt2 = -0.26453031
+ lk2 = -3.0631458e-10
+ vtsswgd = 4.2
+ pvsat = 7.49481800000001e-11
+ vtsswgs = 4.2
+ llc = 0
+ lln = 1
+ lu0 = 3.7246358e-10
+ wk2we = 5e-12
+ pvth0 = 5.2579253999999975e-17
+ mjd = 0.26
+ mjs = 0.26
+ lua = 3.3186753e-17
+ lub = -3.0003129999999985e-27
+ luc = 7.435334e-18
+ lud = 0
+ rbdb = 50
+ pua1 = 6.1201017e-24
+ prwb = 0
+ lwc = 0
+ pub1 = -1.17842519e-32
+ prwg = 0
+ drout = 0.56
+ lwl = 0
+ puc1 = -1.8169327e-24
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 1.2471671e-13
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ nsd = 1e+20
+ pvag = 1.2
+ pbd = 0.52
+ pat = 1.9909584e-10
+ pbs = 0.52
+ pk2 = 1.8168527e-16
+ paigc = -1.0299571e-18
+ pu0 = -1.1106070399999999e-17
+ prt = 0
+ pua = 6.5377716e-24
+ pub = -1.101976303e-32
+ rdsw = 100
+ puc = -3.076481e-25
+ pud = 0
+ voffl = 0
+ rsh = 17.5
+ tcj = 0.00076
+ voffcv = -0.16942
+ wpemod = 1
+ ua1 = 1.4780468e-9
+ ub1 = -2.3055828999999997e-18
+ uc1 = 1.4133161e-10
+ tpb = 0.0014
+ wa0 = -2.130866e-6
+ weta0 = -1.5669611e-7
+ ute = -1
+ wetab = 4.0317659e-8
+ wat = 0.003179234299999999
+ web = 6843.8
+ wec = -25529.0
+ wk2 = 1.5715655e-9
+ wlc = 0
+ wln = 1
+ wu0 = -1.7043296999999997e-11
+ lpclm = 6.3904735e-9
+ xgl = -1.09e-8
+ wkvth0we = 2e-12
+ xgw = 0
+ wua = -1.3239536e-16
+ wub = 1.9940967600000001e-25
+ wuc = 1.2105201e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ cgidl = 0.22
+ trnqsmod = 0
+ rshg = 15.6
+ wtvfbsdoff = 0
+ nfactor = 1
+ pbswd = 0.8
+ pbsws = 0.8
+ tpbswg = 0.0009
+ ltvfbsdoff = 0
+ rgatemod = 0
+ tnjtsswg = 1
+ pdits = 0
+ tnom = 25
+ cigsd = 0.069865
+ toxe = 2.43e-9
+ ptvoff = -1.0763348e-17
+ toxm = 2.43e-9
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ waigsd = 3.1788545e-12
+ nigbacc = 10
+ pk2we = -1e-19
+ diomod = 1
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ ptvfbsdoff = 0
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 2.9779200000000003e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.9779200000000003e-10
+ wags = -2.3477778e-7
+ tnoia = 0
+ nigbinv = 10
+ wcit = 2.2923413999999998e-10
+ peta0 = 7.5477876e-15
+ petab = -1.7674893e-15
+ voff = -0.056267378999999965
+ wketa = -1.07864979e-7
+ acde = 0.4
+ tvfbsdoff = 0.022
+ tpbsw = 0.0019
+ mjswgd = 0.85
+ mjswgs = 0.85
+ vsat = 109805.91299999997
+ wint = 0
+ cjswd = 8.6592e-11
+ cjsws = 8.6592e-11
+ vth0 = 0.24840093900000004
+ tcjswg = 0.001
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ )

.model nch_sf_40 nmos (
+ level = 54
+ wkt1 = -2.3678067e-8
+ wkt2 = -1.1473225e-8
+ wmax = 2.726e-7
+ aigc = 0.011144932
+ wmin = 1.08e-7
+ fnoimod = 1
+ eigbinv = 1.1
+ wua1 = 1.9140234e-16
+ wub1 = -2.6574903999999996e-25
+ wuc1 = 2.7994334999999996e-17
+ bigc = 0.001442
+ wwlc = 0
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ scref = 1e-6
+ ijthsfwd = 0.01
+ cdsc = 0
+ fprout = 300
+ pigcd = 2.621
+ cgbo = 0
+ aigsd = 0.010772574
+ cgdl = 3.31989e-12
+ cgdo = 4.90562e-11
+ xtid = 3
+ xtis = 3
+ xrcrg1 = 12
+ xrcrg2 = 1
+ cgsl = 3.31989e-12
+ cgso = 4.90562e-11
+ cigc = 0.000625
+ lvoff = -1.8479393000000007e-9
+ cigbacc = 0.32875
+ lvsat = 0.00502537152
+ wtvoff = -7.2128996e-10
+ lvth0 = 3.330764800000001e-9
+ ijthsrev = 0.01
+ tnoimod = 0
+ delta = 0.007595625
+ laigc = 5.7720314e-12
+ rnoia = 0
+ rnoib = 0
+ cigbinv = 0.006
+ dmcg = 3.1e-8
+ capmod = 2
+ dmci = 3.1e-8
+ dmdg = 0
+ wku0we = 2e-11
+ pketa = -8.4677334e-15
+ ngate = 8e+20
+ a0 = -5.925916599999999
+ a1 = 0
+ a2 = 1
+ ngcon = 1
+ b0 = 0
+ b1 = 0
+ mobmod = 0
+ wpclm = -7.2101286e-7
+ at = 114373.142
+ cf = 8.15e-11
+ ef = 1.0
+ k1 = 0.274
+ k2 = 0.017123130999999993
+ k3 = -1.8419
+ em = 1000000.0
+ k2we = 5e-5
+ ll = 0
+ lw = 0
+ u0 = 0.01403564272
+ w0 = 0
+ ua = -5.589164400000002e-10
+ ub = -4.454503999999649e-21
+ uc = 3.789344e-10
+ ud = 0
+ version = 4.5
+ wl = 0
+ wr = 1
+ xj = 8.6e-8
+ xl = 4e-9
+ ww = 0
+ xw = 3.4e-9
+ dsub = 0.75
+ dtox = 2.7e-10
+ gbmin = 1e-12
+ tempmod = 0
+ jswgd = 1.28e-13
+ jswgs = 1.28e-13
+ dvt0 = 3.2
+ dvt1 = 0.5
+ dvt2 = -0.35
+ eta0 = -0.288265897
+ aigbacc = 0.02
+ etab = -0.74723747
+ laigsd = -1.5325105e-17
+ pkvth0we = -1.3e-19
+ aigbinv = 0.0163
+ tvoff = 0.0062987975
+ vfbsdoff = 0.02
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = -1.5e-12
+ alpha0 = 2e-10
+ alpha1 = 3.6
+ paramchk = 1
+ ku0we = -0.0007
+ beta0 = 13
+ leta0 = 2.5736964e-8
+ poxedge = 1
+ letab = 2.3120738e-8
+ ppclm = 3.3171145e-14
+ binunit = 2
+ dlcig = 2.5e-9
+ bgidl = 2320000000.0
+ ijthdfwd = 0.01
+ toxref = 3e-9
+ dmcgt = 0
+ keta = -0.51478944
+ tcjsw = 0.000357
+ ijthdrev = 0.01
+ jswd = 1.28e-13
+ jsws = 1.28e-13
+ lcit = 1.910268e-10
+ ltvoff = -2.4217179e-10
+ kt1l = 0
+ jtsswgd = 2.3e-7
+ jtsswgs = 2.3e-7
+ bigsd = 0.00125
+ lint = 0
+ wvoff = 1.82724831e-8
+ lkt1 = -1.7340467e-9
+ lkt2 = -1.1864945e-9
+ lmax = 4.5e-8
+ lmin = 3.6e-8
+ wvsat = 0.022030641400000002
+ lku0we = 2.5e-11
+ pvfbsdoff = 0
+ lpe0 = 9.2e-8
+ wvth0 = -9.679447000000004e-9
+ lpeb = 2.5e-7
+ epsrox = 3.9
+ waigc = 5.1623453e-11
+ minv = -0.3
+ lua1 = 6.0050187e-18
+ lub1 = -8.3060953e-27
+ luc1 = 1.56225695e-17
+ rdsmod = 0
+ lkvth0we = -2e-12
+ ndep = 1e+18
+ igbmod = 1
+ lwlc = 0
+ lketa = 2.6802806000000003e-8
+ moin = 5.1
+ njtsswg = 9
+ xpart = 1
+ pscbe1 = 1000000000.0
+ pscbe2 = 1e-20
+ nigc = 3.083
+ pbswgd = 0.95
+ pbswgs = 0.95
+ xtsswgd = 0.18
+ xtsswgs = 0.18
+ acnqsmod = 0
+ egidl = 0.29734
+ igcmod = 1
+ ckappad = 0.6
+ ckappas = 0.6
+ noff = 2.7195
+ pdiblc1 = 0
+ pdiblc2 = -0.0010804963
+ noia = 3.11e+42
+ noib = 1.22e+22
+ noic = 45200000.0
+ pdiblcb = -0.3
+ rbodymod = 0
+ ntox = 1.0
+ pcit = 1.0471520000000003e-17
+ pclm = 4.6708343
+ ags = 4.2096296
+ bigbacc = 0.002588
+ phin = 0.15
+ paigsd = 4.2297301e-24
+ cjd = 0.001432992
+ cit = 0.0006878963
+ cjs = 0.001432992
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.7
+ bvs = 8.7
+ dlc = 3.26497e-9
+ k3b = 1.9326
+ dwb = 0
+ dwc = 0
+ pkt1 = 4.9311236e-16
+ pkt2 = 5.863609e-16
+ dwg = 0
+ dwj = 0
+ kvth0we = 0.00018
+ wpdiblc2 = 2.3632766e-9
+ permod = 1
+ pvoff = -7.6930684e-16
+ lintnoi = -1.5e-8
+ la0 = 1.3676219000000002e-7
+ cdscb = 0
+ cdscd = 0
+ jsd = 6.11e-7
+ jss = 6.11e-7
+ lat = -0.0037512333199999997
+ bigbinv = 0.004953
+ kt1 = -0.23663458
+ kt2 = -0.073003235
+ lk2 = -3.894925700000001e-9
+ vtsswgd = 4.2
+ pvsat = -8.609877599999999e-10
+ vtsswgs = 4.2
+ llc = 0
+ lln = 1
+ lu0 = -1.9421681300000002e-10
+ wk2we = 5e-12
+ pvth0 = 4.914723899999999e-16
+ mjd = 0.26
+ mjs = 0.26
+ lua = -5.56054081e-17
+ lub = 6.85157957e-26
+ luc = -1.83772219e-17
+ lud = 0
+ rbdb = 50
+ pua1 = -8.5382538e-24
+ prwb = 0
+ lwc = 0
+ pub1 = 1.2835769e-32
+ prwg = 0
+ drout = 0.56
+ lwl = 0
+ puc1 = -2.4016428e-24
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = -7.5523402e-14
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ nsd = 1e+20
+ pvag = 1.2
+ pbd = 0.52
+ pat = 3.8897647999999997e-10
+ pbs = 0.52
+ pk2 = 5.0756697e-16
+ paigc = -1.5534524e-18
+ pu0 = -2.9764861999999995e-18
+ prt = 0
+ pua = -2.8276596999999977e-25
+ pub = -1.3322338800000025e-33
+ rdsw = 100
+ puc = 2.3432717e-24
+ pud = 0
+ voffl = 0
+ rsh = 17.5
+ tcj = 0.00076
+ voffcv = -0.16942
+ wpemod = 1
+ ua1 = 5.4333072e-10
+ ub1 = -8.6088544e-19
+ uc1 = -1.7445285e-10
+ tpb = 0.0014
+ wa0 = 1.9556670799999998e-6
+ weta0 = 9.4960797e-8
+ ute = -1
+ wetab = 3.9258957e-9
+ wat = -0.0006958275000000002
+ web = 6843.8
+ wec = -25529.0
+ wk2 = -5.0790816e-9
+ wlc = 0
+ wln = 1
+ wu0 = -1.8295357e-10
+ lpclm = -1.70821362e-7
+ xgl = -1.09e-8
+ wkvth0we = 2e-12
+ xgw = 0
+ wua = 6.799270000000015e-18
+ wub = 1.704964999999993e-27
+ wuc = -4.1995115e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ cgidl = 0.22
+ trnqsmod = 0
+ rshg = 15.6
+ wtvfbsdoff = 0
+ nfactor = 1
+ pbswd = 0.8
+ pbsws = 0.8
+ tpbswg = 0.0009
+ ltvfbsdoff = 0
+ rgatemod = 0
+ tnjtsswg = 1
+ pdits = 0
+ tnom = 25
+ cigsd = 0.069865
+ toxe = 2.43e-9
+ ptvoff = 2.8458255e-17
+ toxm = 2.43e-9
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ waigsd = 3.1787682e-12
+ nigbacc = 10
+ pk2we = -1e-19
+ diomod = 1
+ dvtp0 = 4e-7
+ dvtp1 = 0.01
+ ptvfbsdoff = 0
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 2.9779200000000003e-10
+ pku0we = -1.5e-18
+ cjswgs = 2.9779200000000003e-10
+ wags = -2.3477778e-7
+ tnoia = 0
+ nigbinv = 10
+ wcit = -1.8493278000000003e-10
+ peta0 = -4.7834008e-15
+ petab = 1.5707054e-17
+ voff = -0.150644936
+ wketa = 1.65035329e-7
+ acde = 0.4
+ tvfbsdoff = 0.022
+ tpbsw = 0.0019
+ mjswgd = 0.85
+ mjswgs = 0.85
+ vsat = -12863.757999999987
+ wint = 0
+ cjswd = 8.6592e-11
+ cjsws = 8.6592e-11
+ vth0 = 0.350032947
+ tcjswg = 0.001
+ mjswd = 0.11
+ mjsws = 0.11
+ agidl = 9.41e-8
+ )

.model pch_ss_1 pmos (
+ level = 54
+ ppclm = 0
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ bigbacc = 0.0054401
+ wpdiblc2 = 0
+ tnom = 25
+ kvth0we = -0.00022
+ tvfbsdoff = 0.1
+ dmcgt = 0
+ toxe = 2.71e-9
+ toxm = 2.67e-9
+ tcjsw = 9.34e-5
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ toxref = 3e-9
+ bigsd = 0.0003327
+ wkvth0we = 0.0
+ wvoff = 0
+ trnqsmod = 0
+ voff = -0.11110337
+ acde = 0.5
+ wvsat = 0
+ wvfbsdoff = 0
+ wvth0 = -2.8e-9
+ lvfbsdoff = 0
+ vsat = 120000
+ wint = 0
+ vth0 = -0.40313527
+ ltvoff = 0
+ wmax = 0.00090001
+ aigc = 0.0068307507
+ wmin = 9.0026e-6
+ a0 = 2.531
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 72000
+ cf = 7.598099999999999e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.00077592763
+ k3 = -2.5823
+ em = 20000000.0
+ lketa = 0
+ ll = 0
+ lw = 0
+ u0 = 0.010075
+ w0 = 0
+ rgatemod = 0
+ ua = 1.297e-10
+ ub = 1.182572e-18
+ uc = 2.014e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 5.6700000000000005e-9
+ ww = 0
+ xpart = 1
+ xw = 3.4e-9
+ nfactor = 1
+ tnjtsswg = 1
+ lku0we = 1.8e-11
+ bigc = 0.0012521
+ egidl = 0.001
+ wwlc = 0
+ epsrox = 3.9
+ cdsc = 0
+ rdsmod = 0
+ cgbo = 0
+ cgdl = 2.799765e-11
+ cgdo = 2.4628259999999997e-11
+ xtid = 3
+ xtis = 3
+ igbmod = 1
+ cgsl = 2.799765e-11
+ cgso = 2.4628259999999997e-11
+ cigc = 0.15259
+ nigbacc = 10
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ pbswgd = 0.8
+ pbswgs = 0.8
+ igcmod = 1
+ nigbinv = 2.171
+ pvoff = 2.5e-17
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ cdscb = 0
+ cdscd = 0
+ pvsat = -5e-11
+ wk2we = 0.0
+ pvth0 = -7e-17
+ drout = 0.56
+ k2we = 5e-5
+ dsub = 0.5
+ dtox = 3.91e-10
+ voffl = 0
+ fnoimod = 1
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ eigbinv = 1.1
+ weta0 = -2e-10
+ permod = 1
+ lpclm = 0
+ eta0 = 0.1672
+ etab = -0.23
+ ijthsfwd = 0.01
+ cgidl = 1
+ voffcv = -0.125
+ wpemod = 1
+ ijthsrev = 0.01
+ pbswd = 0.9
+ pbsws = 0.9
+ cigbacc = 0.245
+ tnoimod = 0
+ pdits = 0
+ cigsd = 0.013281
+ cigbinv = 0.006
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ ppdiblc2 = 0
+ tpbswg = 0.001
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ version = 4.5
+ tempmod = 0
+ tnoia = 0
+ peta0 = -1.5e-17
+ ptvoff = 0
+ aigbacc = 0.012071
+ tpbsw = 0.0025
+ pkvth0we = 0.0
+ pvfbsdoff = 0
+ keta = -0.042350111
+ cjswd = 5.457e-11
+ cjsws = 5.457e-11
+ diomod = 1
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ pditsd = 0
+ pditsl = 0
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ cjswgd = 1.9367000000000001e-10
+ pku0we = 0.0
+ cjswgs = 1.9367000000000001e-10
+ lcit = 0
+ aigbinv = 0.009974
+ vfbsdoff = 0.01
+ wtvfbsdoff = 0
+ kt1l = 0
+ lint = 6.5375218e-9
+ ltvfbsdoff = 0
+ mjswgd = 0.95
+ mjswgs = 0.95
+ lkt1 = -1e-9
+ paramchk = 1
+ lmax = 2.001e-5
+ lmin = 8.99743e-6
+ tcjswg = 0.00128
+ scref = 1e-6
+ lpe0 = 6.44e-8
+ lpeb = 0
+ pigcd = 2.572
+ aigsd = 0.0063636
+ minv = -0.33
+ lvoff = 0
+ poxedge = 1
+ ndep = 1e+18
+ lwlc = 0
+ ijthdfwd = 0.01
+ lvsat = 0.00024
+ moin = 5.5538
+ lvth0 = -6e-10
+ binunit = 2
+ ptvfbsdoff = 0
+ nigc = 2.291
+ delta = 0.018814
+ rnoia = 0
+ rnoib = 0
+ fprout = 200
+ noff = 2.2684
+ ags = 0.8379228
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ ijthdrev = 0.01
+ ngate = 1.7e+20
+ cjd = 0.00144022
+ cit = 5e-6
+ cjs = 0.00144022
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 1.0572421799999999e-8
+ ngcon = 1
+ k3b = 2.1176
+ wpclm = 0
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ lpdiblc2 = 0
+ ntox = -1.9260000000000002
+ wtvoff = 0
+ pcit = 0
+ pclm = 1.484
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ la0 = 0
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0.001
+ kt1 = -0.17107633
+ lk2 = 4e-10
+ kt2 = -0.04747
+ jtsswgd = 1.75e-7
+ phin = 0.15
+ llc = 0
+ jtsswgs = 1.75e-7
+ lln = 1
+ lu0 = 5e-12
+ mjd = 0.335
+ mjs = 0.335
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 0
+ capmod = 2
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ pk2 = 0
+ pkt1 = 0
+ pu0 = 0
+ prt = 0
+ wku0we = 1.5e-11
+ pud = 0
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 1.1969344e-9
+ ub1 = -1.3666143e-18
+ uc1 = 6.873e-11
+ mobmod = 0
+ tpb = 0.0016
+ wa0 = 0
+ lkvth0we = 3e-12
+ ute = -1
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 0
+ wlc = 0
+ wln = 1
+ rbdb = 50
+ prwb = 0
+ wu0 = 0
+ prwg = 0
+ xgl = -8.2e-9
+ xgw = 0
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ rdsw = 200
+ tvoff = 0.0026155642
+ acnqsmod = 0
+ njtsswg = 6.489
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ xtsswgd = 0.32
+ rbodymod = 0
+ xtsswgs = 0.32
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.0026729629
+ ku0we = -0.0007
+ pdiblcb = 0
+ beta0 = 13.32
+ rshg = 14.1
+ leta0 = -5e-10
+ )

.model pch_ss_2 pmos (
+ level = 54
+ aigbinv = 0.009974
+ eta0 = 0.1672
+ tnoia = 0
+ etab = -0.23
+ ijthdfwd = 0.01
+ peta0 = -1.5e-17
+ toxref = 3e-9
+ pvfbsdoff = 0
+ tpbsw = 0.0025
+ cjswd = 5.457e-11
+ cjsws = 5.457e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ ijthdrev = 0.01
+ lpdiblc2 = 7.1311563e-9
+ poxedge = 1
+ ltvoff = -4.7585658e-10
+ binunit = 2
+ scref = 1e-6
+ pigcd = 2.572
+ aigsd = 0.0063636
+ lku0we = 1.8e-11
+ epsrox = 3.9
+ lkvth0we = 3e-12
+ lvoff = -8.0044387e-9
+ lvsat = 0.00024
+ rdsmod = 0
+ lvth0 = -5.7267628e-9
+ ags = 0.80385259
+ igbmod = 1
+ delta = 0.018814
+ laigc = -4.8397409e-11
+ cjd = 0.00144022
+ cit = 5e-6
+ cjs = 0.00144022
+ clc = 1e-7
+ cle = 0.6
+ acnqsmod = 0
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 1.0572421799999999e-8
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ k3b = 2.1176
+ rnoia = 0
+ rnoib = 0
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ keta = -0.040853613
+ pbswgd = 0.8
+ pbswgs = 0.8
+ rbodymod = 0
+ a0 = 2.5747309
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 72000
+ lags = 3.062912e-7
+ ngate = 1.7e+20
+ cf = 7.598099999999999e-11
+ igcmod = 1
+ la0 = -3.9314047e-7
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.0012551498
+ k3 = -2.5823
+ em = 20000000.0
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0.001
+ ll = 0
+ lw = 0
+ kt1 = -0.16652617
+ kt2 = -0.046491549
+ lk2 = 4.708207500000001e-9
+ u0 = 0.010074890100000001
+ ngcon = 1
+ w0 = 0
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ ua = 1.4083134e-10
+ ub = 1.1675774e-18
+ uc = 1.8373185e-11
+ ud = 0
+ llc = 0
+ wpclm = 0
+ lln = 1
+ lcit = 0
+ wl = 0
+ wr = 1
+ lu0 = 5.98779012e-12
+ xj = 1.1e-7
+ xl = 5.6700000000000005e-9
+ ww = 0
+ xw = 3.4e-9
+ mjd = 0.335
+ mjs = 0.335
+ lua = -1.0007073e-16
+ lub = 1.3480174e-25
+ luc = 1.5883665e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ kt1l = 0
+ njs = 1.02
+ pa0 = 0
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ pk2 = 0
+ gbmin = 1e-12
+ pu0 = 0
+ jswgd = 3.69e-13
+ prt = 0
+ jswgs = 3.69e-13
+ pud = 0
+ lint = 6.5375218e-9
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 1.1817684e-9
+ ub1 = -1.3634053e-18
+ uc1 = 6.7786161e-11
+ tpb = 0.0016
+ lkt1 = -4.1906013000000006e-8
+ lkt2 = -8.7962711e-9
+ wa0 = 0
+ lmax = 8.99743e-6
+ ute = -1
+ lmin = 8.974099999999999e-7
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 0
+ wlc = 0
+ wln = 1
+ wu0 = 0
+ xgl = -8.2e-9
+ xgw = 0
+ njtsswg = 6.489
+ lpe0 = 6.44e-8
+ wud = 0
+ wpdiblc2 = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ lpeb = 0
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ minv = -0.33
+ lua1 = 1.3634229e-16
+ lub1 = -2.8849398e-26
+ luc1 = 8.4851172e-18
+ permod = 1
+ ckappad = 0.6
+ ckappas = 0.6
+ ndep = 1e+18
+ pdiblc1 = 0
+ pdiblc2 = 0.0018797309
+ pdiblcb = 0
+ lwlc = 0
+ moin = 5.5538
+ nigc = 2.291
+ tvoff = 0.002668496
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ wkvth0we = 0.0
+ voffcv = -0.125
+ wpemod = 1
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ bigbacc = 0.0054401
+ trnqsmod = 0
+ ku0we = -0.0007
+ beta0 = 13.32
+ kvth0we = -0.00022
+ ntox = -1.9260000000000002
+ pcit = 0
+ pclm = 1.484
+ leta0 = -5e-10
+ lintnoi = -5e-9
+ ppclm = 0
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ phin = 0.15
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ pkt1 = 0
+ rgatemod = 0
+ tpbswg = 0.001
+ tnjtsswg = 1
+ tvfbsdoff = 0.1
+ dmcgt = 0
+ rbdb = 50
+ tcjsw = 9.34e-5
+ prwb = 0
+ prwg = 0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ ptvoff = 0
+ wtvfbsdoff = 0
+ rdsw = 200
+ bigsd = 0.0003327
+ diomod = 1
+ ltvfbsdoff = 0
+ pditsd = 0
+ pditsl = 0
+ nfactor = 1
+ wvoff = 0
+ cjswgd = 1.9367000000000001e-10
+ pku0we = 0.0
+ cjswgs = 1.9367000000000001e-10
+ wvfbsdoff = 0
+ wvsat = 0
+ lvfbsdoff = 0
+ wvth0 = -2.8e-9
+ rshg = 14.1
+ mjswgd = 0.95
+ mjswgs = 0.95
+ tcjswg = 0.00128
+ lketa = -1.3453518e-8
+ ptvfbsdoff = 0
+ nigbacc = 10
+ xpart = 1
+ tnom = 25
+ egidl = 0.001
+ toxe = 2.71e-9
+ toxm = 2.67e-9
+ ijthsfwd = 0.01
+ nigbinv = 2.171
+ fprout = 200
+ xrcrg1 = 12
+ xrcrg2 = 1
+ ijthsrev = 0.01
+ fnoimod = 1
+ voff = -0.110213
+ wtvoff = 0
+ acde = 0.5
+ eigbinv = 1.1
+ pvoff = 2.5e-17
+ vsat = 120000
+ wint = 0
+ vth0 = -0.402565
+ cdscb = 0
+ cdscd = 0
+ wmax = 0.00090001
+ pvsat = -5e-11
+ aigc = 0.0068361342
+ wmin = 9.0026e-6
+ wk2we = 0.0
+ capmod = 2
+ pvth0 = -7e-17
+ drout = 0.56
+ wku0we = 1.5e-11
+ ppdiblc2 = 0
+ mobmod = 0
+ voffl = 0
+ bigc = 0.0012521
+ weta0 = -2e-10
+ cigbacc = 0.245
+ wwlc = 0
+ lpclm = 0
+ cdsc = 0
+ tnoimod = 0
+ cgbo = 0
+ cgidl = 1
+ cgdl = 2.799765e-11
+ cgdo = 2.4628259999999997e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 2.799765e-11
+ cgso = 2.4628259999999997e-11
+ cigc = 0.15259
+ pkvth0we = 0.0
+ cigbinv = 0.006
+ pbswd = 0.9
+ pbsws = 0.9
+ vfbsdoff = 0.01
+ version = 4.5
+ tempmod = 0
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ pdits = 0
+ cigsd = 0.013281
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ dvt0w = 0
+ paramchk = 1
+ dvt1w = 0
+ dvt2w = 0
+ aigbacc = 0.012071
+ k2we = 5e-5
+ dsub = 0.5
+ dtox = 3.91e-10
+ pk2we = 0.0
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ )

.model pch_ss_3 pmos (
+ level = 54
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ nigbacc = 10
+ ijthsrev = 0.01
+ wvoff = 0
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ wvsat = 0
+ ntox = -1.9260000000000002
+ wvth0 = -2.8e-9
+ pcit = 0
+ pclm = 1.484
+ ltvoff = -2.3123852e-10
+ nigbinv = 2.171
+ phin = 0.15
+ lketa = -1.5940244e-8
+ pkt1 = 0
+ ppdiblc2 = 0
+ xpart = 1
+ lku0we = 1.8e-11
+ epsrox = 3.9
+ egidl = 0.001
+ rbdb = 50
+ fnoimod = 1
+ prwb = 0
+ prwg = 0
+ rdsmod = 0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ eigbinv = 1.1
+ igbmod = 1
+ rdsw = 200
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ pbswgd = 0.8
+ pbswgs = 0.8
+ pkvth0we = 0.0
+ igcmod = 1
+ vfbsdoff = 0.01
+ rshg = 14.1
+ cigbacc = 0.245
+ pvoff = 2.5e-17
+ cdscb = 0
+ cdscd = 0
+ pvsat = -5e-11
+ tnoimod = 0
+ wk2we = 0.0
+ pvth0 = -7e-17
+ paramchk = 1
+ drout = 0.56
+ cigbinv = 0.006
+ voffl = 0
+ permod = 1
+ tnom = 25
+ weta0 = -2e-10
+ toxe = 2.71e-9
+ toxm = 2.67e-9
+ a0 = 2.8917556
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ lpclm = 0
+ at = 72000
+ cf = 7.598099999999999e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = 0.0040664684
+ k3 = -2.5823
+ em = 20000000.0
+ ijthdfwd = 0.01
+ version = 4.5
+ ll = 0
+ lw = 0
+ u0 = 0.010306756
+ w0 = 0
+ ua = 1.1413788e-10
+ ub = 1.1978347e-18
+ uc = 4.3035111e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 5.6700000000000005e-9
+ ww = 0
+ xw = 3.4e-9
+ tempmod = 0
+ cgidl = 1
+ voffcv = -0.125
+ wpemod = 1
+ aigbacc = 0.012071
+ ijthdrev = 0.01
+ pbswd = 0.9
+ pbsws = 0.9
+ voff = -0.10886793
+ lpdiblc2 = 1.7469722e-9
+ acde = 0.5
+ vsat = 120000
+ aigbinv = 0.009974
+ wint = 0
+ vth0 = -0.40518963
+ pdits = 0
+ cigsd = 0.013281
+ wmax = 0.00090001
+ aigc = 0.00683106
+ wmin = 9.0026e-6
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ wtvfbsdoff = 0
+ tpbswg = 0.001
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ ltvfbsdoff = 0
+ lkvth0we = 3e-12
+ bigc = 0.0012521
+ wwlc = 0
+ tnoia = 0
+ ptvoff = 0
+ poxedge = 1
+ cdsc = 0
+ peta0 = -1.5e-17
+ cgbo = 0
+ cgdl = 2.799765e-11
+ cgdo = 2.4628259999999997e-11
+ xtid = 3
+ xtis = 3
+ acnqsmod = 0
+ pvfbsdoff = 0
+ cgsl = 2.799765e-11
+ cgso = 2.4628259999999997e-11
+ cigc = 0.15259
+ binunit = 2
+ diomod = 1
+ tpbsw = 0.0025
+ cjswd = 5.457e-11
+ cjsws = 5.457e-11
+ mjswd = 0.01
+ pditsd = 0
+ mjsws = 0.01
+ pditsl = 0
+ rbodymod = 0
+ agidl = 3.2166e-9
+ cjswgd = 1.9367000000000001e-10
+ pku0we = 0.0
+ cjswgs = 1.9367000000000001e-10
+ ptvfbsdoff = 0
+ dmcg = 3.1e-8
+ mjswgd = 0.95
+ dmci = 3.1e-8
+ dmdg = 0
+ mjswgs = 0.95
+ tcjswg = 0.00128
+ k2we = 5e-5
+ jtsswgd = 1.75e-7
+ scref = 1e-6
+ jtsswgs = 1.75e-7
+ wpdiblc2 = 0
+ dsub = 0.5
+ pigcd = 2.572
+ dtox = 3.91e-10
+ aigsd = 0.0063635603
+ ags = 0.82774541
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ lvoff = -9.201547e-9
+ cjd = 0.00144022
+ cit = -8.7888889e-5
+ cjs = 0.00144022
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 1.0572421799999999e-8
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ eta0 = 0.1672
+ etab = -0.23
+ lvsat = 0.00024
+ lvth0 = -3.3908382999999997e-9
+ delta = 0.018814
+ laigc = -4.3881382e-11
+ la0 = -6.7529244e-7
+ fprout = 200
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0.001
+ kt1 = -0.19559142
+ kt2 = -0.048919444
+ lk2 = -2.8032719999999973e-11
+ llc = 0
+ lln = 1
+ lu0 = -2.0037244e-10
+ rnoia = 0
+ rnoib = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ mjd = 0.335
+ mjs = 0.335
+ lua = -7.6313554e-17
+ lub = 1.0787275e-25
+ luc = -6.0654489e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ wkvth0we = 0.0
+ njs = 1.02
+ pa0 = 0
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ pk2 = 0
+ njtsswg = 6.489
+ pu0 = 0
+ prt = 0
+ pud = 0
+ ngate = 1.7e+20
+ trnqsmod = 0
+ wtvoff = 0
+ ngcon = 1
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 1.2804108e-9
+ ub1 = -1.1625424e-18
+ uc1 = 4.6637333e-11
+ wpclm = 0
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ tpb = 0.0016
+ wa0 = 0
+ ute = -1
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 0
+ ckappad = 0.6
+ ckappas = 0.6
+ gbmin = 1e-12
+ wlc = 0
+ wln = 1
+ wu0 = 0
+ xgl = -8.2e-9
+ xgw = 0
+ pdiblc1 = 0
+ pdiblc2 = 0.0079293759
+ wud = 0
+ jswgd = 3.69e-13
+ wwc = 0
+ jswgs = 3.69e-13
+ wwl = 0
+ wwn = 1
+ pdiblcb = 0
+ capmod = 2
+ wku0we = 1.5e-11
+ rgatemod = 0
+ mobmod = 0
+ tnjtsswg = 1
+ bigbacc = 0.0054401
+ kvth0we = -0.00022
+ lintnoi = -5e-9
+ tvoff = 0.0023936443
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ laigsd = 3.5374533e-14
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ keta = -0.03805954
+ lags = 2.8502658e-7
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 8.2671111e-11
+ ku0we = -0.0007
+ beta0 = 13.32
+ kt1l = 0
+ leta0 = -5e-10
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ ppclm = 0
+ lint = 6.5375218e-9
+ lkt1 = -1.6037938999999998e-8
+ lkt2 = -6.6354444e-9
+ dlcig = 2.5e-9
+ lmax = 8.974099999999999e-7
+ bgidl = 1834800000.0
+ lmin = 4.4741e-7
+ lpe0 = 6.44e-8
+ lpeb = 0
+ tvfbsdoff = 0.1
+ minv = -0.33
+ lua1 = 4.8550568e-17
+ nfactor = 1
+ lub1 = -2.0761736e-25
+ luc1 = 2.7307573e-17
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ ndep = 1e+18
+ lwlc = 0
+ ijthsfwd = 0.01
+ moin = 5.5538
+ nigc = 2.291
+ toxref = 3e-9
+ bigsd = 0.0003327
+ )

.model pch_ss_4 pmos (
+ level = 54
+ aigc = 0.0067884199
+ wmin = 9.0026e-6
+ cjd = 0.00144022
+ cit = -0.00054497817
+ cjs = 0.00144022
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 1.38228675e-8
+ scref = 1e-6
+ k3b = 2.1176
+ rgatemod = 0
+ lku0we = 1.8e-11
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ pigcd = 2.572
+ tnjtsswg = 1
+ epsrox = 3.9
+ aigsd = 0.0063636407
+ njtsswg = 6.489
+ lvoff = -3.8830249e-9
+ bigc = 0.0012521
+ la0 = -4.3379389e-8
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0.001
+ rdsmod = 0
+ kt1 = -0.2000222
+ kt2 = -0.054670852
+ lk2 = 1.7630221e-9
+ wwlc = 0
+ llc = -1.18e-13
+ xtsswgd = 0.32
+ lln = 0.7
+ xtsswgs = 0.32
+ lu0 = -4.782545000000001e-10
+ igbmod = 1
+ mjd = 0.335
+ mjs = 0.335
+ lua = -1.5477844e-16
+ lub = 5.0676856e-26
+ luc = -5.2541764e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ lvsat = 0.00024
+ njd = 1.02
+ njs = 1.02
+ pa0 = 0
+ lvth0 = 3.7404646e-9
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ ckappad = 0.6
+ pk2 = 0
+ ckappas = 0.6
+ cdsc = 0
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ pu0 = 0
+ pdiblc1 = 0
+ pdiblc2 = 0.013802718
+ delta = 0.018814
+ cgbo = 0
+ prt = 0
+ cgdl = 2.799765e-11
+ cgdo = 2.4628259999999997e-11
+ pud = 0
+ pdiblcb = 0
+ xtid = 3
+ xtis = 3
+ laigc = -2.5119727e-11
+ pbswgd = 0.8
+ pbswgs = 0.8
+ cgsl = 2.799765e-11
+ cgso = 2.4628259999999997e-11
+ rsh = 15.2
+ tcj = 0.000832
+ cigc = 0.15259
+ ua1 = 1.2553592e-9
+ ub1 = -1.2671808e-18
+ uc1 = 1.0455371e-10
+ rnoia = 0
+ rnoib = 0
+ tpb = 0.0016
+ wa0 = 0
+ igcmod = 1
+ ute = -1
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 0
+ wlc = 0
+ wln = 1
+ wu0 = 0
+ xgl = -8.2e-9
+ xgw = 0
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ ngate = 1.7e+20
+ ngcon = 1
+ wpclm = 0
+ bigbacc = 0.0054401
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ kvth0we = -0.00022
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ k2we = 5e-5
+ vtsswgs = 1.1
+ dsub = 0.5
+ dtox = 3.91e-10
+ permod = 1
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ eta0 = 0.1672
+ ijthsfwd = 0.01
+ etab = -0.23
+ tvoff = 0.002134918
+ voffcv = -0.125
+ wpemod = 1
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ ijthsrev = 0.01
+ wtvfbsdoff = 0
+ ku0we = -0.0007
+ beta0 = 13.32
+ nfactor = 1
+ leta0 = -5e-10
+ ltvfbsdoff = 0
+ ppclm = 0
+ a0 = 1.4555895
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 72000
+ cf = 7.598099999999999e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -4.1106394e-6
+ k3 = -2.5823
+ em = 20000000.0
+ ll = -1.18e-13
+ dlcig = 2.5e-9
+ lw = 0
+ u0 = 0.010938306
+ w0 = 0
+ tpbswg = 0.001
+ ua = 2.9246716e-10
+ ub = 1.3278253e-18
+ uc = 4.119131e-11
+ ud = 0
+ bgidl = 1834800000.0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 5.6700000000000005e-9
+ ww = 0
+ xw = 3.4e-9
+ ppdiblc2 = 0
+ tvfbsdoff = 0.1
+ nigbacc = 10
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ ptvoff = 0
+ ptvfbsdoff = 0
+ diomod = 1
+ nigbinv = 2.171
+ pkvth0we = 0.0
+ bigsd = 0.0003327
+ keta = -0.029364427
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.9367000000000001e-10
+ pku0we = 0.0
+ cjswgs = 1.9367000000000001e-10
+ wvoff = 0
+ lags = 5.4107004e-7
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 2.8379039e-10
+ vfbsdoff = 0.01
+ wvsat = 0
+ kt1l = 0
+ wvth0 = -2.8e-9
+ mjswgd = 0.95
+ mjswgs = 0.95
+ fnoimod = 1
+ eigbinv = 1.1
+ tcjswg = 0.00128
+ lint = 9.7879675e-9
+ lkt1 = -1.4088393000000001e-8
+ lkt2 = -4.1048253e-9
+ paramchk = 1
+ lmax = 4.4741e-7
+ lmin = 2.1410000000000002e-7
+ lketa = -1.9766093e-8
+ lpe0 = 6.44e-8
+ xpart = 1
+ lpeb = 0
+ minv = -0.33
+ lua1 = 5.9573279e-17
+ lub1 = -1.6157647e-25
+ egidl = 0.001
+ luc1 = 1.8243668e-18
+ ndep = 1e+18
+ lwlc = 0
+ ijthdfwd = 0.01
+ moin = 5.5538
+ cigbacc = 0.245
+ fprout = 200
+ nigc = 2.291
+ xrcrg1 = 12
+ xrcrg2 = 1
+ tnoimod = 0
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ ijthdrev = 0.01
+ cigbinv = 0.006
+ wtvoff = 0
+ lpdiblc2 = -8.3729822e-10
+ ntox = -1.9260000000000002
+ pcit = 0
+ pclm = 1.484
+ pvoff = 2.5e-17
+ capmod = 2
+ version = 4.5
+ cdscb = 0
+ cdscd = 0
+ pvsat = -5e-11
+ phin = 0.15
+ wku0we = 1.5e-11
+ tempmod = 0
+ wk2we = 0.0
+ pvth0 = -7e-17
+ drout = 0.56
+ mobmod = 0
+ pkt1 = 0
+ voffl = 0
+ aigbacc = 0.012071
+ lkvth0we = 3e-12
+ weta0 = -2e-10
+ rbdb = 50
+ prwb = 0
+ prwg = 0
+ lpclm = 0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ rdsw = 200
+ aigbinv = 0.009974
+ cgidl = 1
+ acnqsmod = 0
+ rbodymod = 0
+ pbswd = 0.9
+ pbsws = 0.9
+ rshg = 14.1
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ pdits = 0
+ poxedge = 1
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ binunit = 2
+ wpdiblc2 = 0
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ tnom = 25
+ toxe = 2.71e-9
+ toxm = 2.67e-9
+ tnoia = 0
+ toxref = 3e-9
+ peta0 = -1.5e-17
+ pvfbsdoff = 0
+ tpbsw = 0.0025
+ wkvth0we = 0.0
+ cjswd = 5.457e-11
+ cjsws = 5.457e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ trnqsmod = 0
+ voff = -0.12095548
+ acde = 0.5
+ ltvoff = -1.1739897e-10
+ vsat = 120000
+ wint = 0
+ vth0 = -0.42139717
+ wmax = 0.00090001
+ ags = 0.24582847
+ )

.model pch_ss_5 pmos (
+ level = 54
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ pbswgd = 0.8
+ pbswgs = 0.8
+ acnqsmod = 0
+ version = 4.5
+ tempmod = 0
+ igcmod = 1
+ keta = -0.12863898
+ rbodymod = 0
+ lags = 3.2185083e-8
+ aigbacc = 0.012071
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 1.26802573e-10
+ kt1l = 0
+ pvoff = 2.5e-17
+ cdscb = 0
+ cdscd = 0
+ lint = 9.7879675e-9
+ pvsat = -5e-11
+ wk2we = 0.0
+ pvth0 = -7e-17
+ aigbinv = 0.009974
+ lkt1 = -5.7409966e-9
+ lkt2 = -5.2805906e-10
+ drout = 0.56
+ lmax = 2.1410000000000002e-7
+ lmin = 8.833e-8
+ wpdiblc2 = 0
+ lpe0 = 6.44e-8
+ permod = 1
+ lpeb = 0
+ voffl = 0
+ minv = -0.33
+ lua1 = -1.5051887e-16
+ lub1 = 1.742578e-25
+ luc1 = 7.2216103e-18
+ weta0 = -2e-10
+ ndep = 1e+18
+ lpclm = -1.4239795e-8
+ wtvfbsdoff = 0
+ lwlc = 0
+ moin = 5.5538
+ cgidl = 1
+ voffcv = -0.125
+ wpemod = 1
+ nigc = 2.291
+ ltvfbsdoff = 0
+ poxedge = 1
+ wkvth0we = 0.0
+ noff = 2.2684
+ binunit = 2
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ pbswd = 0.9
+ pbsws = 0.9
+ trnqsmod = 0
+ ntox = -1.9260000000000002
+ pcit = 0.0
+ pclm = 1.5514872
+ pdits = 0
+ cigsd = 0.013281
+ phin = 0.15
+ tpbswg = 0.001
+ ptvfbsdoff = 0
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ pkt1 = 0
+ rgatemod = 0
+ tnjtsswg = 1
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ ptvoff = 0
+ rbdb = 50
+ prwb = 0
+ prwg = 0
+ tnoia = 0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ pvfbsdoff = 0
+ rdsw = 200
+ peta0 = -1.5e-17
+ diomod = 1
+ tpbsw = 0.0025
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.9367000000000001e-10
+ pku0we = 0.0
+ cjswgs = 1.9367000000000001e-10
+ cjswd = 5.457e-11
+ a0 = 1.4508547
+ a1 = 0
+ a2 = 1
+ cjsws = 5.457e-11
+ b0 = 0
+ b1 = 0
+ mjswd = 0.01
+ at = 72000
+ cf = 7.598099999999999e-11
+ mjsws = 0.01
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.013949949
+ k3 = -2.5823
+ agidl = 3.2166e-9
+ em = 20000000.0
+ ll = -1.18e-13
+ lw = 0
+ u0 = 0.009522119700000001
+ w0 = 0
+ ua = -3.1871506e-10
+ ub = 1.6925299e-18
+ uc = 2.1642376e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 5.6700000000000005e-9
+ ww = 0
+ xw = 3.4e-9
+ ags = 2.6576055
+ njtsswg = 6.489
+ mjswgd = 0.95
+ mjswgs = 0.95
+ cjd = 0.00144022
+ cit = 0.00019903638
+ cjs = 0.00144022
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ rshg = 14.1
+ bvs = 8.2
+ dlc = 1.38228675e-8
+ xtsswgd = 0.32
+ k3b = 2.1176
+ xtsswgs = 0.32
+ tcjswg = 0.00128
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.016932267
+ pdiblcb = 0
+ la0 = -4.2380342e-8
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0.001
+ kt1 = -0.23958332
+ kt2 = -0.07162235
+ lk2 = 4.7055939000000005e-9
+ scref = 1e-6
+ llc = -1.18e-13
+ lln = 0.7
+ lu0 = -1.7943925e-10
+ mjd = 0.335
+ mjs = 0.335
+ lua = -2.581899e-17
+ lub = -2.6275812e-26
+ luc = -1.1293514e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ pigcd = 2.572
+ njd = 1.02
+ njs = 1.02
+ aigsd = 0.0063636407
+ pa0 = 0
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ pk2 = 0
+ pu0 = 0
+ prt = 0
+ pud = 0
+ tnom = 25
+ lvoff = -1.3382853e-9
+ rsh = 15.2
+ toxe = 2.71e-9
+ toxm = 2.67e-9
+ tcj = 0.000832
+ ua1 = 2.2510566e-9
+ ub1 = -2.8588123e-18
+ uc1 = 7.8974359e-11
+ bigbacc = 0.0054401
+ tpb = 0.0016
+ lvsat = 0.00210474684
+ ijthsfwd = 0.01
+ wa0 = 0
+ ute = -1
+ lvth0 = 5.7644432e-9
+ web = 6628.3
+ wec = -16935.0
+ fprout = 200
+ wk2 = 0
+ wlc = 0
+ wln = 1
+ wu0 = 0
+ xgl = -8.2e-9
+ xgw = 0
+ delta = 0.018814
+ wud = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ laigc = -2.0986759e-11
+ kvth0we = -0.00022
+ rnoia = 0
+ rnoib = 0
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ wtvoff = 0
+ vtsswgs = 1.1
+ ijthsrev = 0.01
+ ngate = 1.7e+20
+ wcit = 0.0
+ ngcon = 1
+ wpclm = 0
+ voff = -0.13301586
+ acde = 0.5
+ gbmin = 1e-12
+ capmod = 2
+ vsat = 111162.27
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ wint = 0
+ vth0 = -0.43098955
+ wku0we = 1.5e-11
+ wmax = 0.00090001
+ aigc = 0.0067688324
+ wmin = 9.0026e-6
+ mobmod = 0
+ ppdiblc2 = 0
+ bigc = 0.0012521
+ wwlc = 0
+ nfactor = 1
+ cdsc = 0
+ cgbo = 0
+ cgdl = 2.799765e-11
+ cgdo = 2.4628259999999997e-11
+ xtid = 3
+ xtis = 3
+ tvoff = 0.0018930751
+ cgsl = 2.799765e-11
+ cgso = 2.4628259999999997e-11
+ cigc = 0.15259
+ xjbvd = 1
+ xjbvs = 1
+ pkvth0we = 0.0
+ lk2we = 0.0
+ vfbsdoff = 0.01
+ ku0we = -0.0007
+ nigbacc = 10
+ beta0 = 13.32
+ leta0 = -5e-10
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ ppclm = 0
+ paramchk = 1
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ nigbinv = 2.171
+ k2we = 5e-5
+ tvfbsdoff = 0.1
+ dsub = 0.5
+ dtox = 3.91e-10
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ eta0 = 0.1672
+ ijthdfwd = 0.01
+ etab = -0.23
+ toxref = 3e-9
+ fnoimod = 1
+ eigbinv = 1.1
+ bigsd = 0.0003327
+ ijthdrev = 0.01
+ wvfbsdoff = 0
+ wvoff = 0
+ lvfbsdoff = 0
+ ltvoff = -6.6370123e-11
+ lpdiblc2 = -1.4976331e-9
+ wvsat = 0.0
+ wvth0 = -2.8e-9
+ cigbacc = 0.245
+ lku0we = 1.8e-11
+ lketa = 1.1808374e-9
+ tnoimod = 0
+ epsrox = 3.9
+ xpart = 1
+ rdsmod = 0
+ cigbinv = 0.006
+ egidl = 0.001
+ lkvth0we = 3e-12
+ igbmod = 1
+ )

.model pch_ss_6 pmos (
+ level = 54
+ wpclm = 0
+ vfbsdoff = 0.01
+ rshg = 14.1
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ nfactor = 1
+ wtvfbsdoff = 0
+ paramchk = 1
+ permod = 1
+ ltvfbsdoff = 0
+ tnom = 25
+ toxe = 2.71e-9
+ toxm = 2.67e-9
+ nigbacc = 10
+ ijthdfwd = 0.01
+ voffcv = -0.125
+ wpemod = 1
+ tvoff = 0.00091084129
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ nigbinv = 2.171
+ ptvfbsdoff = 0
+ ijthdrev = 0.01
+ wcit = 0.0
+ ku0we = -0.0007
+ lpdiblc2 = 0
+ voff = -0.11896044
+ beta0 = 13.32
+ acde = 0.5
+ leta0 = -1.6141465e-9
+ letab = 2.0255694e-8
+ vsat = 211212.03
+ wint = 0
+ vth0 = -0.34669182000000004
+ ppclm = 0
+ tpbswg = 0.001
+ wmax = 0.00090001
+ fnoimod = 1
+ aigc = 0.0067067782
+ wmin = 9.0026e-6
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ eigbinv = 1.1
+ tvfbsdoff = 0.1
+ ptvoff = 0
+ lkvth0we = 3e-12
+ bigc = 0.0012521
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ wwlc = 0
+ diomod = 1
+ cdsc = 0
+ cgbo = 0
+ cgdl = 2.799765e-11
+ cgdo = 2.4628259999999997e-11
+ xtid = 3
+ xtis = 3
+ acnqsmod = 0
+ pditsd = 0
+ pditsl = 0
+ cgsl = 2.799765e-11
+ cjswgd = 1.9367000000000001e-10
+ pku0we = 0.0
+ cgso = 2.4628259999999997e-11
+ cigbacc = 0.245
+ cjswgs = 1.9367000000000001e-10
+ cigc = 0.15259
+ bigsd = 0.0003327
+ rbodymod = 0
+ wvfbsdoff = 0
+ tnoimod = 0
+ lvfbsdoff = 0
+ wvoff = 0
+ mjswgd = 0.95
+ mjswgs = 0.95
+ wvsat = 0.0
+ cigbinv = 0.006
+ wvth0 = -2.8e-9
+ tcjswg = 0.00128
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ version = 4.5
+ lketa = 8.4925319e-9
+ k2we = 5e-5
+ tempmod = 0
+ wpdiblc2 = 0
+ xpart = 1
+ dsub = 0.5
+ dtox = 3.91e-10
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ egidl = 0.001
+ a0 = 3.4166667
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 140456.11
+ cf = 7.598099999999999e-11
+ aigbacc = 0.012071
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.010241786
+ k3 = -2.5823
+ em = 20000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.0055138889
+ w0 = 0
+ ua = -1.1682959e-9
+ ub = 1.3195554999999999e-18
+ uc = -8.7638e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 5.6700000000000005e-9
+ ww = 0
+ xw = 3.4e-9
+ fprout = 200
+ eta0 = 0.17905262
+ etab = -0.44548611
+ xrcrg1 = 12
+ xrcrg2 = 1
+ aigbinv = 0.009974
+ wkvth0we = 0.0
+ wtvoff = 0
+ trnqsmod = 0
+ capmod = 2
+ pvoff = 2.5e-17
+ wku0we = 1.5e-11
+ cdscb = 0
+ cdscd = 0
+ mobmod = 0
+ pvsat = -5e-11
+ wk2we = 0.0
+ pvth0 = -7e-17
+ drout = 0.56
+ poxedge = 1
+ rgatemod = 0
+ voffl = 0
+ tnjtsswg = 1
+ binunit = 2
+ weta0 = -2e-10
+ lpclm = -9.8438889e-8
+ cgidl = 1
+ keta = -0.20642296
+ pbswd = 0.9
+ pbsws = 0.9
+ lags = -2.8753242e-8
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ lcit = 2.4609714e-10
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ kt1l = 0
+ pdits = 0
+ cigsd = 0.013281
+ lint = 0
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ lkt1 = -2.23119e-9
+ lkt2 = 1.5220167e-10
+ lmax = 8.833e-8
+ lmin = 5.233e-8
+ lpe0 = 6.44e-8
+ lpeb = 0
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ minv = -0.33
+ lua1 = -7.3062676e-18
+ lub1 = 1.0038041e-26
+ luc1 = 7.6176556e-18
+ ndep = 1e+18
+ toxref = 3e-9
+ njtsswg = 6.489
+ tnoia = 0
+ ijthsfwd = 0.01
+ lwlc = 0
+ pvfbsdoff = 0
+ moin = 5.5538
+ xtsswgd = 0.32
+ peta0 = -1.5e-17
+ xtsswgs = 0.32
+ nigc = 2.291
+ ckappad = 0.6
+ ckappas = 0.6
+ tpbsw = 0.0025
+ ags = 3.3058856
+ pdiblc1 = 0
+ pdiblc2 = 0.001
+ pdiblcb = 0
+ cjswd = 5.457e-11
+ cjd = 0.00144022
+ cjsws = 5.457e-11
+ cit = -0.00107005811
+ cjs = 0.00144022
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ dlc = 4.0349e-9
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ k3b = 2.1176
+ ijthsrev = 0.01
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ ltvoff = 2.5959859e-11
+ la0 = -2.2716667e-7
+ ntox = -1.9260000000000002
+ pcit = 0.0
+ jsd = 1.5e-7
+ pclm = 2.4472222
+ jss = 1.5e-7
+ lat = -0.0054348744
+ kt1 = -0.27692169
+ kt2 = -0.078859167
+ lk2 = 4.3570266e-9
+ llc = 0
+ lln = 1
+ lu0 = 1.9733444e-10
+ mjd = 0.335
+ bigbacc = 0.0054401
+ mjs = 0.335
+ lua = 5.4041604e-17
+ lub = 8.783782e-27
+ luc = 9.143004e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 0
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ pk2 = 0
+ phin = 0.15
+ pu0 = 0
+ lku0we = 1.8e-11
+ prt = 0
+ pub = 0.0
+ pud = 0
+ kvth0we = -0.00022
+ epsrox = 3.9
+ ppdiblc2 = 0
+ rsh = 15.2
+ scref = 1e-6
+ pkt1 = 0
+ tcj = 0.000832
+ ua1 = 7.2751825e-10
+ ub1 = -1.1117937e-18
+ uc1 = 7.4761111e-11
+ tpb = 0.0016
+ pigcd = 2.572
+ lintnoi = -5e-9
+ wa0 = 0
+ aigsd = 0.0063636407
+ ute = -1
+ web = 6628.3
+ wec = -16935.0
+ bigbinv = 0.00149
+ wk2 = 0
+ rdsmod = 0
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ wlc = 0
+ wln = 1
+ wu0 = 0
+ xgl = -8.2e-9
+ xgw = 0
+ wub = 0.0
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ igbmod = 1
+ lvoff = -2.6594942e-9
+ rbdb = 50
+ prwb = 0
+ prwg = 0
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ rbpb = 50
+ rbpd = 50
+ lvsat = -0.0072999309
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ lvth0 = -2.159537e-9
+ pbswgd = 0.8
+ pbswgs = 0.8
+ rdsw = 200
+ delta = 0.018814
+ laigc = -1.5153664e-11
+ igcmod = 1
+ rnoia = 0
+ rnoib = 0
+ pkvth0we = 0.0
+ ngate = 1.7e+20
+ ngcon = 1
+ )

.model pch_ss_7 pmos (
+ level = 54
+ voffl = 0
+ dsub = 0.5
+ dtox = 3.91e-10
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ weta0 = -2e-10
+ ptvfbsdoff = 0
+ lpclm = -4.4240467e-8
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ eta0 = 0.18948293
+ ijthsfwd = 0.01
+ voffcv = -0.125
+ wpemod = 1
+ etab = -0.27185615
+ cgidl = 1
+ ijthsrev = 0.01
+ pbswd = 0.9
+ pbsws = 0.9
+ njtsswg = 6.489
+ tpbswg = 0.001
+ pdits = 0
+ cigsd = 0.013281
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ ppdiblc2 = 0
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.001
+ pdiblcb = 0
+ pk2we = 0.0
+ ptvoff = 0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ ags = 2.81014
+ pvfbsdoff = 0
+ tnoia = 0
+ diomod = 1
+ cjd = 0.00144022
+ cit = -0.0040245511999999995
+ cjs = 0.00144022
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 4.0349e-9
+ peta0 = -1.5e-17
+ k3b = 2.1176
+ pditsd = 0
+ pditsl = 0
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ bigbacc = 0.0054401
+ dwj = 0
+ cjswgd = 1.9367000000000001e-10
+ pku0we = 0.0
+ cjswgs = 1.9367000000000001e-10
+ tpbsw = 0.0025
+ pkvth0we = 0.0
+ keta = 0.048888889
+ cjswd = 5.457e-11
+ kvth0we = -0.00022
+ cjsws = 5.457e-11
+ la0 = -1.5788889e-7
+ jsd = 1.5e-7
+ mjswd = 0.01
+ jss = 1.5e-7
+ lat = 0.0052661578
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ kt1 = -0.090229195
+ kt2 = -0.087042222
+ lk2 = 4.7353879e-9
+ llc = 0
+ lln = 1
+ lu0 = -6.7628889e-11
+ mjd = 0.335
+ mjs = 0.335
+ lua = -4.5270917e-17
+ lub = -3.5537642e-26
+ luc = -2.161341e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ lintnoi = -5e-9
+ njd = 1.02
+ mjswgd = 0.95
+ njs = 1.02
+ mjswgs = 0.95
+ pa0 = 0
+ bigbinv = 0.00149
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ jswd = 3.69e-13
+ vtsswgd = 1.1
+ pk2 = 0
+ jsws = 3.69e-13
+ vtsswgs = 1.1
+ vfbsdoff = 0.01
+ lcit = 4.1745849e-10
+ pu0 = 0
+ tcjswg = 0.00128
+ prt = 0
+ pub = 0.0
+ pud = 0
+ kt1l = 0
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 1.0031266e-9
+ ub1 = -2.5489021e-18
+ uc1 = 1.9738889e-10
+ tpb = 0.0016
+ wa0 = 0
+ ute = -1
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 0
+ lint = 0
+ wlc = 0
+ wln = 1
+ wu0 = 0
+ xgl = -8.2e-9
+ xgw = 0
+ paramchk = 1
+ wub = 0.0
+ wud = 0
+ wwc = 0
+ lkt1 = -1.3059355e-8
+ lkt2 = 6.2681889e-10
+ wwl = 0
+ wwn = 1
+ lmax = 5.233e-8
+ lmin = 4.333e-8
+ scref = 1e-6
+ lpe0 = 6.44e-8
+ lpeb = 0
+ pigcd = 2.572
+ aigsd = 0.0063636407
+ minv = -0.33
+ lvoff = -4.1866651e-9
+ lua1 = -2.3291554e-17
+ lub1 = 9.339033e-26
+ luc1 = 5.0524444e-19
+ fprout = 200
+ ndep = 1e+18
+ lvsat = 0.00262611572
+ ijthdfwd = 0.01
+ xrcrg1 = 12
+ xrcrg2 = 1
+ lwlc = 0
+ lvth0 = -4.1797439e-9
+ moin = 5.5538
+ delta = 0.018814
+ laigc = -9.9932362e-12
+ nigc = 2.291
+ nfactor = 1
+ rnoia = 0
+ rnoib = 0
+ wtvoff = 0
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ ijthdrev = 0.01
+ ngate = 1.7e+20
+ ngcon = 1
+ wpclm = 0
+ lpdiblc2 = 0
+ capmod = 2
+ ntox = -1.9260000000000002
+ pcit = 0.0
+ wku0we = 1.5e-11
+ pclm = 1.5127667
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ nigbacc = 10
+ a0 = 2.2222222
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = -44044.444
+ mobmod = 0
+ cf = 7.598099999999999e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.016765256
+ k3 = -2.5823
+ em = 20000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.010082222200000001
+ w0 = 0
+ ua = 5.4398899e-10
+ ub = 2.0837185999999998e-18
+ uc = 4.42645e-10
+ ud = 0
+ phin = 0.15
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 5.6700000000000005e-9
+ ww = 0
+ xw = 3.4e-9
+ pkt1 = 0
+ nigbinv = 2.171
+ lkvth0we = 3e-12
+ rbdb = 50
+ prwb = 0
+ prwg = 0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ rdsw = 200
+ tvoff = 0.0051729841
+ acnqsmod = 0
+ fnoimod = 1
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ eigbinv = 1.1
+ rbodymod = 0
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = -2.2191043e-9
+ rshg = 14.1
+ letab = 1.0185157e-8
+ ppclm = 0
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ tvfbsdoff = 0.1
+ cigbacc = 0.245
+ wpdiblc2 = 0
+ tnoimod = 0
+ tnom = 25
+ dmcgt = 0
+ toxref = 3e-9
+ tcjsw = 9.34e-5
+ toxe = 2.71e-9
+ toxm = 2.67e-9
+ cigbinv = 0.006
+ bigsd = 0.0003327
+ wkvth0we = 0.0
+ version = 4.5
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ tempmod = 0
+ ltvoff = -2.2124443e-10
+ wvoff = 0
+ wcit = 0.0
+ trnqsmod = 0
+ voff = -0.092629909
+ wvsat = 0.0
+ acde = 0.5
+ wvth0 = -2.8e-9
+ aigbacc = 0.012071
+ vsat = 40073.291
+ wint = 0
+ vth0 = -0.31186069000000005
+ lku0we = 1.8e-11
+ wmax = 0.00090001
+ aigc = 0.0066178053
+ wmin = 9.0026e-6
+ epsrox = 3.9
+ lketa = -6.3155556e-9
+ rgatemod = 0
+ xpart = 1
+ aigbinv = 0.009974
+ tnjtsswg = 1
+ rdsmod = 0
+ igbmod = 1
+ egidl = 0.001
+ bigc = 0.0012521
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ wwlc = 0
+ pbswgd = 0.8
+ pbswgs = 0.8
+ cdsc = 0
+ cgbo = 0
+ igcmod = 1
+ cgdl = 2.799765e-11
+ cgdo = 2.4628259999999997e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 2.799765e-11
+ cgso = 2.4628259999999997e-11
+ cigc = 0.15259
+ wtvfbsdoff = 0
+ poxedge = 1
+ binunit = 2
+ ltvfbsdoff = 0
+ pvoff = 2.5e-17
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ cdscb = 0
+ cdscd = 0
+ pvsat = -5e-11
+ wk2we = 0.0
+ pvth0 = -7e-17
+ drout = 0.56
+ permod = 1
+ k2we = 5e-5
+ )

.model pch_ss_8 pmos (
+ level = 54
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ wkvth0we = 0.0
+ cigbacc = 0.245
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ trnqsmod = 0
+ ku0we = -0.0007
+ tnoimod = 0
+ beta0 = 13.32
+ leta0 = 1.6323128000000002e-9
+ ntox = -1.9260000000000002
+ letab = 3.9337702e-9
+ pcit = 0.0
+ pclm = 1.0208333
+ tpbswg = 0.001
+ cigbinv = 0.006
+ ppclm = 0
+ phin = 0.15
+ dlcig = 2.5e-9
+ tvfbsdoff = 0.1
+ bgidl = 1834800000.0
+ pkt1 = 0.0
+ rgatemod = 0
+ ptvoff = 0
+ tnjtsswg = 1
+ version = 4.5
+ tempmod = 0
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ diomod = 1
+ rbdb = 50
+ prwb = 0
+ prwg = 0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ aigbacc = 0.012071
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.9367000000000001e-10
+ pku0we = 0.0
+ cjswgs = 1.9367000000000001e-10
+ rdsw = 200
+ bigsd = 0.0003327
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ mjswgd = 0.95
+ mjswgs = 0.95
+ wvoff = 0
+ aigbinv = 0.009974
+ tcjswg = 0.00128
+ wvsat = 0.0
+ wvth0 = -2.8e-9
+ rshg = 14.1
+ lketa = 8.0381778e-9
+ xpart = 1
+ poxedge = 1
+ egidl = 0.001
+ tnom = 25
+ fprout = 200
+ toxe = 2.71e-9
+ toxm = 2.67e-9
+ xrcrg1 = 12
+ xrcrg2 = 1
+ binunit = 2
+ ijthsfwd = 0.01
+ wtvoff = 0
+ ijthsrev = 0.01
+ wcit = 0.0
+ capmod = 2
+ voff = -0.10032114
+ wku0we = 1.5e-11
+ acde = 0.5
+ pvoff = 2.5e-17
+ mobmod = 0
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ vsat = 142298.12
+ wint = 0
+ vth0 = -0.38882998
+ cdscb = 0
+ cdscd = 0
+ wkt1 = 0.0
+ pvsat = -5e-11
+ wmax = 0.00090001
+ wk2we = 0.0
+ pvth0 = -7e-17
+ aigc = 0.0065563017
+ wmin = 9.0026e-6
+ drout = 0.56
+ ppdiblc2 = 0
+ voffl = 0
+ weta0 = -2e-10
+ wetab = 0
+ bigc = 0.0012521
+ wwlc = 0
+ lpclm = -2.0135733e-8
+ laigsd = -2.1777787e-18
+ cdsc = 0
+ cgidl = 1
+ njtsswg = 6.489
+ cgbo = 0
+ cgdl = 2.799765e-11
+ cgdo = 2.4628259999999997e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 2.799765e-11
+ cgso = 2.4628259999999997e-11
+ cigc = 0.15259
+ a0 = -0.19555556
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ xtsswgd = 0.32
+ pkvth0we = 0.0
+ xtsswgs = 0.32
+ at = 76220.0
+ cf = 7.598099999999999e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.012217534
+ k3 = -2.5823
+ em = 20000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.0055777778
+ w0 = 0
+ ua = -1.1794951e-9
+ ub = 1.1293934e-18
+ uc = 5.0701667e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 5.6700000000000005e-9
+ ww = 0
+ xw = 3.4e-9
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.001
+ pbswd = 0.9
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ pbsws = 0.9
+ pdiblcb = 0
+ vfbsdoff = 0.01
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ pdits = 0
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ paramchk = 1
+ bigbacc = 0.0054401
+ k2we = 5e-5
+ ags = 1.0774289
+ dsub = 0.5
+ kvth0we = -0.00022
+ dtox = 3.91e-10
+ cjd = 0.00144022
+ cit = 0.00447277333
+ pk2we = 0.0
+ cjs = 0.00144022
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ dlc = 4.0349e-9
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ k3b = 2.1176
+ toxref = 3e-9
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ pvfbsdoff = 0
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ tnoia = 0
+ ijthdfwd = 0.01
+ eta0 = 0.11088258
+ etab = -0.14427684
+ la0 = -3.9417778e-8
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = -0.0006268000000000001
+ kt1 = -0.30391077
+ kt2 = -0.08425
+ lk2 = 4.5125495e-9
+ peta0 = -1.5e-17
+ llc = 0
+ lln = 1
+ lu0 = 1.5308889e-10
+ petab = 0
+ mjd = 0.335
+ mjs = 0.335
+ lua = 3.9179804e-17
+ lub = 1.1224222200000001e-26
+ luc = -2.4081867e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 0
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0.0
+ pbs = 0.75
+ tpbsw = 0.0025
+ pk2 = 0
+ pu0 = 0
+ prt = 0
+ pub = 0.0
+ pud = 0
+ cjswd = 5.457e-11
+ cjsws = 5.457e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ ltvoff = -2.4936809e-11
+ agidl = 3.2166e-9
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 1.4917512e-9
+ ub1 = -1.5908843e-18
+ uc1 = 1.6325556e-10
+ ijthdrev = 0.01
+ tpb = 0.0016
+ wa0 = 0
+ ute = -1
+ wat = 0.0
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 0
+ wlc = 0
+ wln = 1
+ lpdiblc2 = 0
+ wu0 = 0
+ xgl = -8.2e-9
+ xgw = 0
+ wub = 0.0
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ lku0we = 1.8e-11
+ epsrox = 3.9
+ nfactor = 1
+ scref = 1e-6
+ rdsmod = 0
+ pigcd = 2.572
+ aigsd = 0.0063636407
+ igbmod = 1
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ wtvfbsdoff = 0
+ lvoff = -3.8097951e-9
+ lkvth0we = 3e-12
+ pbswgd = 0.8
+ pbswgs = 0.8
+ lvsat = -0.0023829014
+ lvth0 = -4.08253058e-10
+ igcmod = 1
+ ltvfbsdoff = 0
+ delta = 0.018814
+ nigbacc = 10
+ laigc = -6.97956e-12
+ acnqsmod = 0
+ rnoia = 0
+ rnoib = 0
+ keta = -0.24404444
+ rbodymod = 0
+ ngate = 1.7e+20
+ lags = 8.4902844e-8
+ ngcon = 1
+ nigbinv = 2.171
+ wpclm = 0
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 1.088669999999988e-12
+ kt1l = 0
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ ptvfbsdoff = 0
+ lint = 0
+ permod = 1
+ lkt1 = -2.5889574e-9
+ lkt2 = 4.9e-10
+ lmax = 4.333e-8
+ lmin = 3.6e-8
+ fnoimod = 1
+ wpdiblc2 = 0
+ lpe0 = 6.44e-8
+ lpeb = 0
+ eigbinv = 1.1
+ minv = -0.33
+ lua1 = -4.7234158e-17
+ lub1 = 4.6447457e-26
+ luc1 = 2.1777778e-18
+ voffcv = -0.125
+ wpemod = 1
+ ndep = 1e+18
+ lwlc = 0
+ moin = 5.5538
+ tvoff = 0.0011667062
+ nigc = 2.291
+ )

.model pch_ss_9 pmos (
+ level = 54
+ vtsswgs = 1.1
+ ags = 0.82538676
+ vsat = 121084.96
+ wint = 0
+ vth0 = -0.40247063000000005
+ pdits = 0
+ cjd = 0.00144022
+ cit = 5e-6
+ cjs = 0.00144022
+ clc = 1e-7
+ cle = 0.6
+ cigsd = 0.013281
+ bvd = 8.2
+ bvs = 8.2
+ wkt1 = -1.0361455e-8
+ wkt2 = -3.8769913e-9
+ dlc = 1.0572421799999999e-8
+ wmax = 9.0026e-6
+ dvt0w = 0
+ k3b = 2.1176
+ dvt1w = 0
+ aigc = 0.0068303602
+ dvt2w = 0
+ wmin = 9.025999999999999e-7
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ ptvoff = 0
+ waigsd = 1.9139418e-12
+ la0 = 0
+ pk2we = 0.0
+ jsd = 1.5e-7
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ jss = 1.5e-7
+ lat = 0.001
+ wua1 = -3.2799159e-16
+ kt1 = -0.16992583
+ lk2 = 4e-10
+ kt2 = -0.04703951
+ wub1 = 5.9231251e-25
+ wuc1 = -8.7396626e-17
+ llc = 0
+ lln = 1
+ lu0 = 5e-12
+ mjd = 0.335
+ mjs = 0.335
+ lkvth0we = 3e-12
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ diomod = 1
+ pvfbsdoff = 0
+ njd = 1.02
+ bigc = 0.0012521
+ njs = 1.02
+ wute = -7.8572347e-8
+ pa0 = 0
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ wwlc = 0
+ pk2 = 0
+ tnoia = 0
+ pu0 = 0
+ pditsd = 0
+ pditsl = 0
+ prt = 0
+ pud = 0
+ cjswgd = 1.9367000000000001e-10
+ pku0we = 0.0
+ cjswgs = 1.9367000000000001e-10
+ rsh = 15.2
+ tcj = 0.000832
+ peta0 = -1.5e-17
+ cdsc = 0
+ ua1 = 1.2333536e-9
+ ub1 = -1.432383e-18
+ uc1 = 7.8434267e-11
+ cgbo = 0
+ tpb = 0.0016
+ cgdl = 2.799765e-11
+ cgdo = 2.4628259999999997e-11
+ acnqsmod = 0
+ xtid = 3
+ xtis = 3
+ wketa = 2.2362589e-8
+ wa0 = 3.3745816e-7
+ ute = -0.99127556
+ web = 6628.3
+ wec = -16935.0
+ cgsl = 2.799765e-11
+ cgso = 2.4628259999999997e-11
+ wk2 = -2.287053e-9
+ tpbsw = 0.0025
+ cigc = 0.15259
+ wlc = 0
+ wln = 1
+ wu0 = -8.6631049e-11
+ xgl = -8.2e-9
+ xgw = 0
+ wua = -1.124189e-16
+ wub = -6.7100784e-26
+ wuc = -2.319496e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ cjswd = 5.457e-11
+ nfactor = 1
+ cjsws = 5.457e-11
+ mjswd = 0.01
+ mjswgd = 0.95
+ mjsws = 0.01
+ mjswgs = 0.95
+ agidl = 3.2166e-9
+ rbodymod = 0
+ tcjswg = 0.00128
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ nigbacc = 10
+ scref = 1e-6
+ k2we = 5e-5
+ wpdiblc2 = 3.6469361e-10
+ pigcd = 2.572
+ dsub = 0.5
+ aigsd = 0.0063633875
+ dtox = 3.91e-10
+ fprout = 200
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ lvoff = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ nigbinv = 2.171
+ lvsat = 0.00024
+ eta0 = 0.16744607
+ etab = -0.23671111
+ lvth0 = -6e-10
+ delta = 0.018814
+ wtvoff = -9.8925647e-11
+ rnoia = 0
+ rnoib = 0
+ wkvth0we = 0.0
+ fnoimod = 1
+ ngate = 1.7e+20
+ capmod = 2
+ trnqsmod = 0
+ eigbinv = 1.1
+ ngcon = 1
+ wpclm = -3.01194e-7
+ wku0we = 1.5e-11
+ mobmod = 0
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ rgatemod = 0
+ tnjtsswg = 1
+ cigbacc = 0.245
+ tnoimod = 0
+ tvoff = 0.0026265487
+ cigbinv = 0.006
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ keta = -0.044833188
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ version = 4.5
+ jswd = 3.69e-13
+ ku0we = -0.0007
+ jsws = 3.69e-13
+ lcit = 0
+ tempmod = 0
+ beta0 = 13.32
+ leta0 = -5e-10
+ kt1l = 0
+ ppclm = 0
+ aigbacc = 0.012071
+ lint = 6.5375218e-9
+ tvfbsdoff = 0.1
+ dlcig = 2.5e-9
+ lkt1 = -1e-9
+ bgidl = 1834800000.0
+ lmax = 2.001e-5
+ lmin = 8.99743e-6
+ lpe0 = 6.44e-8
+ lpeb = 0
+ a0 = 2.4935296
+ a1 = 0
+ a2 = 1
+ toxref = 3e-9
+ b0 = 0
+ b1 = 0
+ at = 72000
+ cf = 7.598099999999999e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.00052197993
+ k3 = -2.5823
+ em = 20000000.0
+ aigbinv = 0.009974
+ minv = -0.33
+ ll = 0
+ lw = 0
+ u0 = 0.0100846193
+ w0 = 0
+ ua = 1.4218267e-10
+ ub = 1.1900227e-18
+ uc = 2.2715501e-11
+ ud = 0
+ dmcgt = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 5.6700000000000005e-9
+ ww = 0
+ xw = 3.4e-9
+ tcjsw = 9.34e-5
+ ndep = 1e+18
+ ijthsfwd = 0.01
+ lwlc = 0
+ moin = 5.5538
+ nigc = 2.291
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ bigsd = 0.0003327
+ ltvoff = 0
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ ijthsrev = 0.01
+ wvoff = 5.5905393e-9
+ poxedge = 1
+ wvsat = -0.0097711764
+ wvth0 = -8.785454e-9
+ ntox = -1.9260000000000002
+ pcit = 0
+ pclm = 1.5174437
+ binunit = 2
+ lku0we = 1.8e-11
+ wtvfbsdoff = 0
+ waigc = 3.5172206e-12
+ epsrox = 3.9
+ phin = 0.15
+ lketa = 0
+ rdsmod = 0
+ ltvfbsdoff = 0
+ ppdiblc2 = 0
+ pkt1 = 0
+ xpart = 1
+ igbmod = 1
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ egidl = 0.001
+ pbswgd = 0.8
+ pbswgs = 0.8
+ rbdb = 50
+ prwb = 0
+ prwg = 0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ igcmod = 1
+ rbsb = 50
+ pvag = 2.1
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ rdsw = 200
+ ptvfbsdoff = 0
+ pkvth0we = 0.0
+ vfbsdoff = 0.01
+ rshg = 14.1
+ pvoff = 2.5e-17
+ cdscb = 0
+ cdscd = 0
+ permod = 1
+ pvsat = -5e-11
+ wk2we = 0.0
+ pvth0 = -7e-17
+ paramchk = 1
+ njtsswg = 6.489
+ drout = 0.56
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ voffl = 0
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.0026324684
+ weta0 = -2.4161431e-9
+ tnom = 25
+ pdiblcb = 0
+ wetab = 6.0440267e-8
+ voffcv = -0.125
+ wpemod = 1
+ lpclm = 0
+ toxe = 2.71e-9
+ toxm = 2.67e-9
+ ijthdfwd = 0.01
+ cgidl = 1
+ bigbacc = 0.0054401
+ wags = 1.128996e-7
+ ijthdrev = 0.01
+ pbswd = 0.9
+ pbsws = 0.9
+ kvth0we = -0.00022
+ lpdiblc2 = 0
+ voff = -0.11172412
+ tpbswg = 0.001
+ acde = 0.5
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ )

.model pch_ss_10 pmos (
+ level = 54
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ lags = 3.1017116e-7
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 0
+ nfactor = 1
+ kt1l = 0
+ paramchk = 1
+ scref = 1e-6
+ pigcd = 2.572
+ aigsd = 0.0063633879
+ lint = 6.5375218e-9
+ lkt1 = -4.2907452e-8
+ lkt2 = -8.3161855e-9
+ lmax = 8.99743e-6
+ lvoff = -7.1040424e-9
+ lmin = 8.974099999999999e-7
+ lpe0 = 6.44e-8
+ lpeb = 0
+ lvsat = 0.00024
+ lvth0 = -5.0817542e-9
+ ijthdfwd = 0.01
+ toxref = 3e-9
+ nigbacc = 10
+ minv = -0.33
+ delta = 0.018814
+ lua1 = 2.9697696e-17
+ lub1 = 1.2607181e-25
+ luc1 = -4.744495e-18
+ laigc = -4.752933e-11
+ wtvfbsdoff = 0
+ ndep = 1e+18
+ rnoia = 0
+ rnoib = 0
+ lute = -8.6179201e-9
+ lwlc = 0
+ tvfbsdoff = 0.1
+ moin = 5.5538
+ ltvfbsdoff = 0
+ pketa = -2.2807538e-14
+ nigc = 2.291
+ ngate = 1.7e+20
+ ijthdrev = 0.01
+ nigbinv = 2.171
+ ngcon = 1
+ wpclm = -3.01194e-7
+ lpdiblc2 = 7.3300428e-9
+ ltvoff = -4.2514859e-10
+ gbmin = 1e-12
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ pags = -3.4942959e-14
+ ntox = -1.9260000000000002
+ pcit = 0
+ pclm = 1.5174437
+ fnoimod = 1
+ wvfbsdoff = 0
+ lku0we = 1.8e-11
+ ptvfbsdoff = 0
+ eigbinv = 1.1
+ lvfbsdoff = 0
+ epsrox = 3.9
+ phin = 0.15
+ lkvth0we = 3e-12
+ pkt1 = 9.0189586e-15
+ pkt2 = -4.3236504e-15
+ rdsmod = 0
+ igbmod = 1
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ tvoff = 0.0026738399
+ pbswgd = 0.8
+ acnqsmod = 0
+ pbswgs = 0.8
+ rbdb = 50
+ pua1 = 9.6044121e-22
+ prwb = 0
+ pub1 = -1.3952204e-30
+ prwg = 0
+ puc1 = 1.1914589e-22
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ pute = 7.7612988e-14
+ igcmod = 1
+ cigbacc = 0.245
+ rdsw = 200
+ rbodymod = 0
+ tnoimod = 0
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = -5e-10
+ cigbinv = 0.006
+ ppclm = 0
+ paigsd = 3.3403436e-20
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ rshg = 14.1
+ version = 4.5
+ wpdiblc2 = 5.6393415e-10
+ permod = 1
+ tempmod = 0
+ ags = 0.79088496
+ dmcgt = 0
+ cjd = 0.00144022
+ cit = 5e-6
+ cjs = 0.00144022
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ tcjsw = 9.34e-5
+ dlc = 1.0572421799999999e-8
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ aigbacc = 0.012071
+ tnom = 25
+ la0 = -3.6651331e-7
+ toxe = 2.71e-9
+ toxm = 2.67e-9
+ jsd = 1.5e-7
+ voffcv = -0.125
+ wpemod = 1
+ jss = 1.5e-7
+ lat = 0.001
+ kt1 = -0.16526426
+ kt2 = -0.046114462
+ lk2 = 4.9045048e-9
+ llc = 0
+ lln = 1
+ bigsd = 0.0003327
+ lu0 = -1.1444212000000002e-10
+ mjd = 0.335
+ mjs = 0.335
+ lua = -1.1601528e-16
+ lub = 1.1870612e-25
+ luc = 1.7407612e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = -2.3980423e-13
+ wkvth0we = 0.0
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ pk2 = -1.7678537e-15
+ aigbinv = 0.009974
+ wvoff = 6.4925381e-9
+ pu0 = 1.0845918e-15
+ prt = 0
+ pua = 1.4359661e-22
+ pub = 1.4495718e-31
+ puc = -1.3724663e-23
+ pud = 0
+ trnqsmod = 0
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 1.2300502e-9
+ ub1 = -1.4464065e-18
+ uc1 = 7.8962019e-11
+ wvsat = -0.0097711764
+ tpb = 0.0016
+ wvth0 = -8.139308799999998e-9
+ wa0 = 3.6413271e-7
+ ute = -0.99031694
+ wags = 1.1678647e-7
+ web = 6628.3
+ wec = -16935.0
+ wk2 = -2.0904063e-9
+ wlc = 0
+ wln = 1
+ wu0 = -2.0727529e-10
+ xgl = -8.2e-9
+ waigc = 4.3868453e-12
+ xgw = 0
+ wua = -1.2839182e-16
+ wub = -8.3225053e-26
+ wuc = -2.1668301e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ voff = -0.11093391
+ acde = 0.5
+ tpbswg = 0.001
+ lketa = -1.0921036e-8
+ vsat = 121084.96
+ wint = 0
+ xpart = 1
+ vth0 = -0.40197210000000005
+ rgatemod = 0
+ wkt1 = -1.1364676e-8
+ wkt2 = -3.3960513e-9
+ poxedge = 1
+ wmax = 9.0026e-6
+ tnjtsswg = 1
+ aigc = 0.0068356471
+ wmin = 9.025999999999999e-7
+ egidl = 0.001
+ binunit = 2
+ ptvoff = -4.5667618e-16
+ waigsd = 1.9102262e-12
+ wua1 = -4.3482598e-16
+ wub1 = 7.4750944e-25
+ wuc1 = -1.0064978e-16
+ bigc = 0.0012521
+ wute = -8.7205605e-8
+ diomod = 1
+ wwlc = 0
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.9367000000000001e-10
+ pku0we = 0.0
+ cjswgs = 1.9367000000000001e-10
+ cdsc = 0
+ cgbo = 0
+ cgdl = 2.799765e-11
+ cgdo = 2.4628259999999997e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 2.799765e-11
+ cgso = 2.4628259999999997e-11
+ cigc = 0.15259
+ pvoff = -8.0839692e-15
+ jtsswgd = 1.75e-7
+ pvfbsdoff = 0
+ mjswgd = 0.95
+ jtsswgs = 1.75e-7
+ mjswgs = 0.95
+ cdscb = 0
+ cdscd = 0
+ tcjswg = 0.00128
+ pvsat = -5e-11
+ wk2we = 0.0
+ pvth0 = -5.8789325e-15
+ drout = 0.56
+ paigc = -7.8179264e-18
+ a0 = 2.5342986
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 72000
+ cf = 7.598099999999999e-11
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.0010230372
+ k3 = -2.5823
+ em = 20000000.0
+ voffl = 0
+ ll = 0
+ lw = 0
+ u0 = 0.010097905400000001
+ w0 = 0
+ ua = 1.5508759e-10
+ ub = 1.1768184e-18
+ uc = 2.077917e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 5.6700000000000005e-9
+ ww = 0
+ xw = 3.4e-9
+ weta0 = -2.4161431e-9
+ wetab = 6.0440267e-8
+ k2we = 5e-5
+ lpclm = 0
+ dsub = 0.5
+ dtox = 3.91e-10
+ ijthsfwd = 0.01
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ njtsswg = 6.489
+ cgidl = 1
+ fprout = 200
+ xrcrg1 = 12
+ xrcrg2 = 1
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ eta0 = 0.16744607
+ etab = -0.23671111
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.0018171133
+ pdiblcb = 0
+ pbswd = 0.9
+ wtvoff = -4.8127407e-11
+ pbsws = 0.9
+ ijthsrev = 0.01
+ pdits = 0
+ capmod = 2
+ cigsd = 0.013281
+ wku0we = 1.5e-11
+ bigbacc = 0.0054401
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ mobmod = 0
+ ppdiblc2 = -1.7911725e-15
+ kvth0we = -0.00022
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ tnoia = 0
+ peta0 = -1.5e-17
+ wketa = 2.4899578e-8
+ laigsd = -3.7090202e-15
+ tpbsw = 0.0025
+ pkvth0we = 0.0
+ cjswd = 5.457e-11
+ cjsws = 5.457e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ keta = -0.04361839
+ vfbsdoff = 0.01
+ )

.model pch_ss_11 pmos (
+ level = 54
+ egidl = 0.001
+ ltvfbsdoff = 0
+ toxref = 3e-9
+ ijthsfwd = 0.01
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ tnom = 25
+ toxe = 2.71e-9
+ toxm = 2.67e-9
+ ijthsrev = 0.01
+ ptvfbsdoff = 0
+ ltvoff = -2.603747e-10
+ pvfbsdoff = 0
+ wags = -5.7105665e-9
+ pvoff = 6.0760934e-15
+ cdscb = 0
+ cdscd = 0
+ pvsat = -5e-11
+ wk2we = 0.0
+ voff = -0.10782222
+ njtsswg = 6.489
+ pvth0 = 3.1763785e-15
+ drout = 0.56
+ acde = 0.5
+ paigc = 1.0166993e-17
+ lku0we = 1.8e-11
+ xtsswgd = 0.32
+ vsat = 121084.96
+ xtsswgs = 0.32
+ wint = 0
+ ppdiblc2 = 8.932051e-16
+ vth0 = -0.40346699
+ epsrox = 3.9
+ voffl = 0
+ wkt1 = 3.9882501e-9
+ wkt2 = -1.3862366e-8
+ ckappad = 0.6
+ wmax = 9.0026e-6
+ ckappas = 0.6
+ aigc = 0.0068328167
+ wmin = 9.025999999999999e-7
+ pdiblc1 = 0
+ pdiblc2 = 0.0082016634
+ pdiblcb = 0
+ weta0 = -2.4161431e-9
+ rdsmod = 0
+ wetab = 6.0440267e-8
+ igbmod = 1
+ lpclm = 0
+ wua1 = 1.0350058e-15
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ wub1 = -1.41997e-24
+ wuc1 = 5.1522417e-17
+ cgidl = 1
+ pbswgd = 0.8
+ bigc = 0.0012521
+ pbswgs = 0.8
+ wwlc = 0
+ bigbacc = 0.0054401
+ igcmod = 1
+ pkvth0we = 0.0
+ cdsc = 0
+ cgbo = 0
+ cgdl = 2.799765e-11
+ cgdo = 2.4628259999999997e-11
+ xtid = 3
+ xtis = 3
+ pbswd = 0.9
+ pbsws = 0.9
+ kvth0we = -0.00022
+ cgsl = 2.799765e-11
+ cgso = 2.4628259999999997e-11
+ cigc = 0.15259
+ vfbsdoff = 0.01
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ pdits = 0
+ cigsd = 0.013281
+ paigsd = -3.7089273e-20
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ paramchk = 1
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ permod = 1
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ k2we = 5e-5
+ tnoia = 0
+ dsub = 0.5
+ dtox = 3.91e-10
+ ijthdfwd = 0.01
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ peta0 = -1.5e-17
+ voffcv = -0.125
+ wpemod = 1
+ wketa = -2.3248862e-8
+ tpbsw = 0.0025
+ eta0 = 0.16744607
+ nfactor = 1
+ etab = -0.23671111
+ cjswd = 5.457e-11
+ cjsws = 5.457e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ ijthdrev = 0.01
+ lpdiblc2 = 1.6477933e-9
+ nigbacc = 10
+ tpbswg = 0.001
+ scref = 1e-6
+ pigcd = 2.572
+ aigsd = 0.0063633394
+ lvoff = -9.8734428e-9
+ nigbinv = 2.171
+ ptvoff = 2.6240046e-16
+ lkvth0we = 3e-12
+ waigsd = 1.9894315e-12
+ lvsat = 0.00024
+ lvth0 = -3.7513085e-9
+ delta = 0.018814
+ diomod = 1
+ laigc = -4.5010295e-11
+ acnqsmod = 0
+ rnoia = 0
+ rnoib = 0
+ tvfbsdoff = 0.1
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.9367000000000001e-10
+ pku0we = 0.0
+ cjswgs = 1.9367000000000001e-10
+ fnoimod = 1
+ pketa = 2.0044574e-14
+ rbodymod = 0
+ ngate = 1.7e+20
+ eigbinv = 1.1
+ ngcon = 1
+ wpclm = -3.01194e-7
+ keta = -0.035478054
+ mjswgd = 0.95
+ mjswgs = 0.95
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ tcjswg = 0.00128
+ lags = 2.7680102e-7
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 8.2671111e-11
+ kt1l = 0
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ wpdiblc2 = -2.4522204e-9
+ lint = 6.5375218e-9
+ cigbacc = 0.245
+ lkt1 = -1.5522155e-8
+ lkt2 = -7.1896716e-9
+ lmax = 8.974099999999999e-7
+ lmin = 4.4741e-7
+ tnoimod = 0
+ lpe0 = 6.44e-8
+ lpeb = 0
+ fprout = 200
+ minv = -0.33
+ cigbinv = 0.006
+ lua1 = 8.7159171e-17
+ lub1 = -2.6689299e-25
+ luc1 = 2.9116076e-17
+ tvoff = 0.0024887007
+ xrcrg1 = 12
+ xrcrg2 = 1
+ ndep = 1e+18
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ lwlc = 0
+ moin = 5.5538
+ wkvth0we = 0.0
+ wtvoff = -8.5607868e-10
+ nigc = 2.291
+ version = 4.5
+ a0 = 2.8862723
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ trnqsmod = 0
+ at = 72000
+ cf = 7.598099999999999e-11
+ tempmod = 0
+ ef = 1.15
+ ku0we = -0.0007
+ k1 = 0.30425
+ k2 = 0.0046668319
+ k3 = -2.5823
+ em = 20000000.0
+ ll = 0
+ lw = 0
+ beta0 = 13.32
+ u0 = 0.0100844338
+ w0 = 0
+ ua = 8.4190146e-11
+ ub = 1.1838278e-18
+ uc = 4.9200634e-11
+ ud = 0
+ leta0 = -5e-10
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 5.6700000000000005e-9
+ ww = 0
+ xw = 3.4e-9
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ capmod = 2
+ ppclm = 0
+ aigbacc = 0.012071
+ wku0we = 1.5e-11
+ pags = 7.4079401e-14
+ ags = 0.8283795
+ dlcig = 2.5e-9
+ mobmod = 0
+ bgidl = 1834800000.0
+ ntox = -1.9260000000000002
+ pcit = 0
+ pclm = 1.5174437
+ cjd = 0.00144022
+ cit = -8.7888889e-5
+ cjs = 0.00144022
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 1.0572421799999999e-8
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ rgatemod = 0
+ tnjtsswg = 1
+ phin = 0.15
+ aigbinv = 0.009974
+ dmcgt = 0
+ la0 = -6.797699e-7
+ pkt1 = -4.6451461e-15
+ jsd = 1.5e-7
+ pkt2 = 4.9913693e-15
+ tcjsw = 9.34e-5
+ jss = 1.5e-7
+ lat = 0.001
+ kt1 = -0.19603426
+ kt2 = -0.047380208
+ lk2 = -1.594787e-10
+ llc = 0
+ lln = 1
+ lu0 = -1.0245246e-10
+ mjd = 0.335
+ mjs = 0.335
+ lua = -5.2916554e-17
+ lub = 1.1246778e-25
+ luc = -7.8874906e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 4.0323955e-14
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ pk2 = 1.1838025e-15
+ pu0 = -8.8186737e-16
+ laigsd = 3.9492818e-14
+ prt = 0
+ pua = -2.1071339e-22
+ pub = -4.1382897e-32
+ puc = 1.6409308e-23
+ pud = 0
+ rbdb = 50
+ pua1 = -3.4770908e-22
+ prwb = 0
+ pub1 = 5.3383631e-31
+ prwg = 0
+ rsh = 15.2
+ puc1 = -1.6287371e-23
+ tcj = 0.000832
+ ua1 = 1.1654868e-9
+ ub1 = -1.004873e-18
+ uc1 = 4.0916434e-11
+ bigsd = 0.0003327
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ tpb = 0.0016
+ wa0 = 4.9381936e-8
+ ute = -1
+ web = 6628.3
+ wec = -16935.0
+ wk2 = -5.406874e-9
+ rdsw = 200
+ wlc = 0
+ wln = 1
+ wu0 = 2.0022293e-9
+ xgl = -8.2e-9
+ wvoff = -9.4176445e-9
+ xgw = 0
+ wua = 2.6970929e-16
+ wub = 1.2614582e-25
+ wuc = -5.5526695e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ poxedge = 1
+ wvsat = -0.0097711764
+ wvth0 = -1.83138011e-8
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ binunit = 2
+ waigc = -1.5820929e-11
+ rshg = 14.1
+ lketa = -1.8165935e-8
+ xpart = 1
+ wtvfbsdoff = 0
+ )

.model pch_ss_12 pmos (
+ level = 54
+ wkvth0we = 0.0
+ pketa = 2.9922765e-15
+ ngate = 1.7e+20
+ ngcon = 1
+ cigbacc = 0.245
+ ltvoff = -1.0992228e-10
+ wpclm = -3.01194e-7
+ trnqsmod = 0
+ gbmin = 1e-12
+ tnoimod = 0
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ cigbinv = 0.006
+ lku0we = 1.8e-11
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ epsrox = 3.9
+ rgatemod = 0
+ tnjtsswg = 1
+ rdsmod = 0
+ version = 4.5
+ igbmod = 1
+ tempmod = 0
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ pbswgd = 0.8
+ pbswgs = 0.8
+ tvoff = 0.0021467634
+ aigbacc = 0.012071
+ igcmod = 1
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ ku0we = -0.0007
+ ags = 0.29253015
+ aigbinv = 0.009974
+ beta0 = 13.32
+ keta = -0.031086208
+ leta0 = -5e-10
+ cjd = 0.00144022
+ cit = -0.00056559017
+ cjs = 0.00144022
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 1.38228675e-8
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ lags = 5.1257474e-7
+ ppclm = 0
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 2.9285967e-10
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ kt1l = 0
+ la0 = -1.4357692e-8
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0.001
+ kt1 = -0.19916819
+ kt2 = -0.054700402
+ lk2 = 1.8250990000000001e-9
+ permod = 1
+ llc = -1.18e-13
+ lln = 0.7
+ lu0 = -4.757604500000001e-10
+ mjd = 0.335
+ mjs = 0.335
+ lua = -1.6078561e-16
+ lub = 5.7693033e-26
+ luc = -4.8483261e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ lint = 9.7879675e-9
+ pa0 = -2.613694e-13
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ pk2 = -5.5906497e-16
+ lkt1 = -1.4143224e-8
+ lkt2 = -3.9687861e-9
+ pu0 = -2.2461433e-17
+ lmax = 4.4741e-7
+ prt = 0
+ pua = 5.4100623e-23
+ pub = -6.3187687e-32
+ puc = -3.6550877e-24
+ pud = 0
+ dmcgt = 0
+ lmin = 2.1410000000000002e-7
+ poxedge = 1
+ tcjsw = 9.34e-5
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 1.2176874e-9
+ ub1 = -1.2376668e-18
+ lpe0 = 6.44e-8
+ uc1 = 1.0272662e-10
+ lpeb = 0
+ tpb = 0.0016
+ wa0 = 7.3504866e-7
+ ijthsfwd = 0.01
+ ute = -1
+ web = 6628.3
+ wec = -16935.0
+ wk2 = -1.4458115e-9
+ binunit = 2
+ voffcv = -0.125
+ wpemod = 1
+ wlc = 0
+ wln = 1
+ minv = -0.33
+ wu0 = 4.9034036e-11
+ xgl = -8.2e-9
+ xgw = 0
+ lua1 = 6.4190903e-17
+ lub1 = -1.6446372e-25
+ wua = -3.3214073e-16
+ wub = 1.7570216e-25
+ wuc = -9.9257962e-18
+ wud = 0
+ luc1 = 1.9195943e-18
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ ndep = 1e+18
+ bigsd = 0.0003327
+ lwlc = 0
+ moin = 5.5538
+ wvoff = 6.3544834e-9
+ nigc = 2.291
+ ijthsrev = 0.01
+ wvsat = -0.0097711764
+ wvth0 = -1.145475961e-8
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ waigc = 4.9938134e-12
+ tpbswg = 0.001
+ jtsswgd = 1.75e-7
+ pags = 2.5662868e-13
+ jtsswgs = 1.75e-7
+ ntox = -1.9260000000000002
+ pcit = -8.1677938e-17
+ lketa = -2.0098347e-8
+ pclm = 1.5174437
+ xpart = 1
+ ppdiblc2 = -1.9289508e-16
+ phin = 0.15
+ ptvoff = -6.733506e-17
+ egidl = 0.001
+ waigsd = 1.9051377e-12
+ pkt1 = 4.9381461e-16
+ pkt2 = -1.2251691e-15
+ diomod = 1
+ pditsd = 0
+ pditsl = 0
+ rbdb = 50
+ cjswgd = 1.9367000000000001e-10
+ pku0we = 0.0
+ pua1 = -4.1586322e-23
+ prwb = 0
+ pub1 = 2.600258e-32
+ prwg = 0
+ cjswgs = 1.9367000000000001e-10
+ puc1 = -8.5761835e-25
+ njtsswg = 6.489
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ pkvth0we = 0.0
+ rdsw = 200
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ ckappad = 0.6
+ ckappas = 0.6
+ mjswgd = 0.95
+ mjswgs = 0.95
+ pdiblc1 = 0
+ pdiblc2 = 0.01380092
+ pvfbsdoff = 0
+ pdiblcb = 0
+ vfbsdoff = 0.01
+ pvoff = -8.636429e-16
+ tcjswg = 0.00128
+ cdscb = 0
+ cdscd = 0
+ pvsat = -5e-11
+ wk2we = 0.0
+ pvth0 = 1.5840135e-16
+ drout = 0.56
+ paramchk = 1
+ rshg = 14.1
+ paigc = 1.0085061e-18
+ bigbacc = 0.0054401
+ voffl = 0
+ weta0 = -2.4161431e-9
+ kvth0we = -0.00022
+ wetab = 6.0440267e-8
+ lpclm = 0
+ lintnoi = -5e-9
+ fprout = 200
+ ijthdfwd = 0.01
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ xrcrg1 = 12
+ xrcrg2 = 1
+ cgidl = 1
+ tnom = 25
+ toxe = 2.71e-9
+ toxm = 2.67e-9
+ wtvoff = -1.0667978e-10
+ pbswd = 0.9
+ pbsws = 0.9
+ ijthdrev = 0.01
+ lpdiblc2 = -8.1587971e-10
+ capmod = 2
+ wags = -4.2059528e-7
+ wku0we = 1.5e-11
+ wcit = 1.8563168e-10
+ pdits = 0
+ cigsd = 0.013281
+ mobmod = 0
+ voff = -0.12166106
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ acde = 0.5
+ vsat = 121084.96
+ wint = 0
+ vth0 = -0.42043621000000003
+ nfactor = 1
+ pk2we = 0.0
+ wkt1 = -7.6912059e-9
+ wkt2 = 2.6613072e-10
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ wmax = 9.0026e-6
+ aigc = 0.0067878654
+ wmin = 9.025999999999999e-7
+ lkvth0we = 3e-12
+ tnoia = 0
+ a0 = 1.3739719
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 72000
+ wua1 = 3.3927227e-16
+ cf = 7.598099999999999e-11
+ wub1 = -2.6580249e-25
+ wuc1 = 1.6454797e-17
+ ef = 1.15
+ k1 = 0.30425
+ k2 = 0.00015642806
+ k3 = -2.5823
+ em = 20000000.0
+ peta0 = -1.5e-17
+ ll = -1.18e-13
+ lw = 0
+ u0 = 0.010932861
+ w0 = 0
+ ua = 3.293471e-10
+ ub = 1.3083159e-18
+ uc = 4.2293442e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 5.6700000000000005e-9
+ ww = 0
+ bigc = 0.0012521
+ xw = 3.4e-9
+ wketa = 1.5506359e-8
+ wwlc = 0
+ acnqsmod = 0
+ tpbsw = 0.0025
+ nigbacc = 10
+ cjswd = 5.457e-11
+ cjsws = 5.457e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ cdsc = 0
+ cgbo = 0
+ rbodymod = 0
+ cgdl = 2.799765e-11
+ cgdo = 2.4628259999999997e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 2.799765e-11
+ cgso = 2.4628259999999997e-11
+ cigc = 0.15259
+ wtvfbsdoff = 0
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ nigbinv = 2.171
+ ltvfbsdoff = 0
+ scref = 1e-6
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ pigcd = 2.572
+ wpdiblc2 = 1.6189099e-11
+ aigsd = 0.0063634291
+ fnoimod = 1
+ lvoff = -3.7843526e-9
+ eigbinv = 1.1
+ k2we = 5e-5
+ toxref = 3e-9
+ lvsat = 0.00024
+ dsub = 0.5
+ dtox = 3.91e-10
+ lvth0 = 3.7151071000000003e-9
+ ptvfbsdoff = 0
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ delta = 0.018814
+ laigc = -2.5231709e-11
+ tvfbsdoff = 0.1
+ rnoia = 0
+ rnoib = 0
+ eta0 = 0.16744607
+ etab = -0.23671111
+ )

.model pch_ss_13 pmos (
+ level = 54
+ pags = 7.0037917e-14
+ lku0we = 1.8e-11
+ pvth0 = -1.99305891e-15
+ drout = 0.56
+ epsrox = 3.9
+ ntox = -1.9260000000000002
+ pcit = -1.9980153999999996e-17
+ pclm = 1.5924795
+ paigc = -7.3857349e-19
+ voffl = 0
+ rdsmod = 0
+ phin = 0.15
+ igbmod = 1
+ weta0 = -2.4161431e-9
+ wetab = 6.0440267e-8
+ lkvth0we = 3e-12
+ pkt1 = 2.8071967e-16
+ pkt2 = -8.6151083e-16
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ lpclm = -1.5832542e-8
+ pbswgd = 0.8
+ pbswgs = 0.8
+ cgidl = 1
+ igcmod = 1
+ acnqsmod = 0
+ rbdb = 50
+ pua1 = -5.7774504e-23
+ prwb = 0
+ pub1 = 1.0356474e-31
+ prwg = 0
+ puc1 = 6.0450908e-24
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ rdsw = 200
+ rbodymod = 0
+ pbswd = 0.9
+ pbsws = 0.9
+ nfactor = 1
+ pdits = 0
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ permod = 1
+ rshg = 14.1
+ nigbacc = 10
+ wpdiblc2 = -2.9527442e-9
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ tnoia = 0
+ voffcv = -0.125
+ wpemod = 1
+ nigbinv = 2.171
+ peta0 = -1.5e-17
+ tnom = 25
+ wketa = 2.8638443e-8
+ toxe = 2.71e-9
+ toxm = 2.67e-9
+ tpbsw = 0.0025
+ cjswd = 5.457e-11
+ cjsws = 5.457e-11
+ mjswd = 0.01
+ wkvth0we = 0.0
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ trnqsmod = 0
+ fnoimod = 1
+ eigbinv = 1.1
+ wags = 4.6372111e-7
+ tpbswg = 0.001
+ wcit = -1.0677104000000002e-10
+ voff = -0.13366619
+ acde = 0.5
+ scref = 1e-6
+ vsat = 111258.71
+ wint = 0
+ vth0 = -0.43116074000000004
+ rgatemod = 0
+ pigcd = 2.572
+ aigsd = 0.0063634291
+ wkt1 = -6.6812774e-9
+ wkt2 = -1.4573681e-9
+ tnjtsswg = 1
+ ptvoff = -1.8786066e-17
+ wmax = 9.0026e-6
+ aigc = 0.0067673585
+ wmin = 9.025999999999999e-7
+ lvoff = -1.2512704e-9
+ waigsd = 1.9051377e-12
+ cigbacc = 0.245
+ lvsat = 0.00231332323
+ diomod = 1
+ lvth0 = 5.9779736000000005e-9
+ wua1 = 4.1599351e-16
+ wub1 = -6.3339564e-25
+ wuc1 = -1.6259465e-17
+ tnoimod = 0
+ delta = 0.018814
+ laigc = -2.090475e-11
+ pditsd = 0
+ pditsl = 0
+ tvfbsdoff = 0.1
+ bigc = 0.0012521
+ cjswgd = 1.9367000000000001e-10
+ pku0we = 0.0
+ cjswgs = 1.9367000000000001e-10
+ wwlc = 0
+ rnoia = 0
+ rnoib = 0
+ cigbinv = 0.006
+ cdsc = 0
+ pketa = 2.2140676e-16
+ ngate = 1.7e+20
+ cgbo = 0
+ cgdl = 2.799765e-11
+ cgdo = 2.4628259999999997e-11
+ xtid = 3
+ xtis = 3
+ ngcon = 1
+ mjswgd = 0.95
+ cgsl = 2.799765e-11
+ cgso = 2.4628259999999997e-11
+ mjswgs = 0.95
+ wpclm = -3.6917638e-7
+ cigc = 0.15259
+ tcjswg = 0.00128
+ version = 4.5
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ tempmod = 0
+ jswgs = 3.69e-13
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ aigbacc = 0.012071
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ k2we = 5e-5
+ fprout = 200
+ aigbinv = 0.009974
+ dsub = 0.5
+ dtox = 3.91e-10
+ xrcrg1 = 12
+ xrcrg2 = 1
+ ijthsfwd = 0.01
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ tvoff = 0.0019304691
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ ags = 2.6061153
+ wtvoff = -3.3676979e-10
+ eta0 = 0.16744607
+ etab = -0.23671111
+ cjd = 0.00144022
+ cit = 0.00021089184
+ cjs = 0.00144022
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 1.38228675e-8
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ ijthsrev = 0.01
+ ku0we = -0.0007
+ beta0 = 13.32
+ capmod = 2
+ leta0 = -5e-10
+ la0 = -4.2186937e-8
+ poxedge = 1
+ wku0we = 1.5e-11
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0.00128821144
+ kt1 = -0.23884145
+ kt2 = -0.071460529
+ lk2 = 4.7288295e-9
+ llc = -1.18e-13
+ lln = 0.7
+ lu0 = -1.7951509e-10
+ mjd = 0.335
+ ppclm = 1.4344283e-14
+ mjs = 0.335
+ lua = -2.3141614e-17
+ lub = -3.0092793e-26
+ luc = -1.1168748e-18
+ lud = 0
+ lwc = 0
+ mobmod = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = -1.7418058e-15
+ nsd = 1e+20
+ binunit = 2
+ pbd = 0.75
+ pat = -2.5956322e-9
+ pbs = 0.75
+ pk2 = -2.0925962e-16
+ dlcig = 2.5e-9
+ pu0 = 6.8306111e-19
+ bgidl = 1834800000.0
+ prt = 0
+ pua = -2.4112447e-23
+ pub = 3.4375734e-32
+ puc = -1.1236355e-25
+ pud = 0
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 2.2048659e-9
+ ub1 = -2.7884819e-18
+ ppdiblc2 = 4.3354985e-16
+ uc1 = 8.0779763e-11
+ tpb = 0.0016
+ wa0 = -4.9541389e-7
+ ute = -1
+ wat = 0.012301575
+ web = 6628.3
+ wec = -16935.0
+ wk2 = -3.1036812e-9
+ wlc = 0
+ wln = 1
+ wu0 = -6.065551e-11
+ xgl = -8.2e-9
+ xgw = 0
+ wua = 3.8537331e-17
+ wub = -2.8668372e-25
+ wuc = -2.6715958e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ wtvfbsdoff = 0
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ bigsd = 0.0003327
+ ltvfbsdoff = 0
+ pkvth0we = 0.0
+ wvoff = 5.8569161e-9
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ wvsat = -0.0008685858999999997
+ vfbsdoff = 0.01
+ keta = -0.13181891
+ wvth0 = -1.2581604999999999e-9
+ waigc = 1.3273811e-11
+ lags = 2.4408277e-8
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 1.29021159e-10
+ a0 = 1.505864
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ kt1l = 0
+ ptvfbsdoff = 0
+ at = 70634.069
+ paramchk = 1
+ cf = 7.598099999999999e-11
+ lketa = 1.156253e-9
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.013605325
+ k3 = -2.5823
+ em = 20000000.0
+ ll = -1.18e-13
+ lw = 0
+ u0 = 0.0095288547
+ w0 = 0
+ xpart = 1
+ ua = -3.2299413e-10
+ ub = 1.7243624e-18
+ uc = 2.4608838e-11
+ ud = 0
+ njtsswg = 6.489
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 5.6700000000000005e-9
+ ww = 0
+ xw = 3.4e-9
+ lint = 9.7879675e-9
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ lkt1 = -5.7721669e-9
+ lkt2 = -4.3239941e-10
+ egidl = 0.001
+ lmax = 2.1410000000000002e-7
+ lmin = 8.833e-8
+ toxref = 3e-9
+ ckappad = 0.6
+ ckappas = 0.6
+ lpe0 = 6.44e-8
+ pdiblc1 = 0
+ pdiblc2 = 0.017260131
+ lpeb = 0
+ pdiblcb = 0
+ ijthdfwd = 0.01
+ minv = -0.33
+ lua1 = -1.4410376e-16
+ lub1 = 1.6275827e-25
+ luc1 = 6.550381e-18
+ ndep = 1e+18
+ lwlc = 0
+ moin = 5.5538
+ bigbacc = 0.0054401
+ nigc = 2.291
+ ltvoff = -6.4284173e-11
+ ijthdrev = 0.01
+ pvfbsdoff = 0
+ lpdiblc2 = -1.5457732e-9
+ kvth0we = -0.00022
+ pvoff = -7.586562e-16
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ cdscb = 0
+ cdscd = 0
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ pvsat = -1.92842639e-9
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ wk2we = 0.0
+ )

.model pch_ss_14 pmos (
+ level = 54
+ cjd = 0.00144022
+ poxedge = 1
+ cit = -0.00109875246
+ wua1 = -1.4703955e-15
+ cjs = 0.00144022
+ clc = 1e-7
+ cle = 0.6
+ wub1 = 2.631826e-24
+ bvd = 8.2
+ wuc1 = 2.762344e-16
+ bvs = 8.2
+ igcmod = 1
+ dlc = 4.0349e-9
+ k3b = 2.1176
+ tvoff = 0.0011122833
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ bigc = 0.0012521
+ wwlc = 0
+ xjbvd = 1
+ binunit = 2
+ xjbvs = 1
+ lk2we = 0.0
+ pkvth0we = 0.0
+ la0 = -2.3326483e-7
+ jsd = 1.5e-7
+ cdsc = 0
+ jss = 1.5e-7
+ lat = -0.0055502639
+ kt1 = -0.2764195
+ kt2 = -0.075556865
+ lk2 = 4.2809157e-9
+ llc = 0
+ cgbo = 0
+ lln = 1
+ cgdl = 2.799765e-11
+ cgdo = 2.4628259999999997e-11
+ lu0 = 2.1144492000000002e-10
+ xtid = 3
+ xtis = 3
+ mjd = 0.335
+ mjs = 0.335
+ lua = 5.4621428e-17
+ lub = 1.2704216999999999e-26
+ luc = 1.0238844e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ cgsl = 2.799765e-11
+ njs = 1.02
+ cgso = 2.4628259999999997e-11
+ pa0 = 5.4920056e-14
+ cigc = 0.15259
+ ku0we = -0.0007
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 1.0391973e-9
+ pbs = 0.75
+ pk2 = 6.854543e-16
+ beta0 = 13.32
+ vfbsdoff = 0.01
+ pu0 = -1.2707891e-16
+ leta0 = -1.14826039e-9
+ prt = 0
+ pua = -5.2218942e-24
+ pub = -3.5307490999999995e-32
+ puc = -9.869134e-24
+ pud = 0
+ letab = 2.0996791e-8
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 8.9078668e-10
+ ub1 = -1.404024e-18
+ uc1 = 4.4088848e-11
+ ppclm = 7.4853015e-14
+ tpb = 0.0016
+ wa0 = -1.0981997e-6
+ ute = -1
+ wat = -0.026366825
+ web = 6628.3
+ wec = -16935.0
+ wk2 = -1.2621914e-8
+ wlc = 0
+ dlcig = 2.5e-9
+ permod = 1
+ wln = 1
+ wu0 = 1.2985144e-9
+ xgl = -8.2e-9
+ xgw = 0
+ bgidl = 1834800000.0
+ wua = -1.62426e-16
+ wub = 4.546272399999999e-25
+ wuc = 7.7079472e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ paramchk = 1
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ k2we = 5e-5
+ voffcv = -0.125
+ wpemod = 1
+ dsub = 0.5
+ dtox = 3.91e-10
+ ijthdfwd = 0.01
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ bigsd = 0.0003327
+ eta0 = 0.17434246
+ etab = -0.46008122
+ njtsswg = 6.489
+ wvoff = -4.5993296e-9
+ ijthdrev = 0.01
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ wvsat = -0.07177826600000001
+ wvth0 = -4.8319501e-8
+ lpdiblc2 = 0
+ ckappad = 0.6
+ tpbswg = 0.001
+ ckappas = 0.6
+ waigc = -2.1370578e-11
+ pdiblc1 = 0
+ pdiblc2 = 0.00081573526
+ pdiblcb = 0
+ lketa = 9.0137227e-9
+ xpart = 1
+ ptvoff = 1.200911e-16
+ waigsd = 1.9051377e-12
+ bigbacc = 0.0054401
+ egidl = 0.001
+ lkvth0we = 3e-12
+ diomod = 1
+ kvth0we = -0.00022
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.9367000000000001e-10
+ pku0we = 0.0
+ cjswgs = 1.9367000000000001e-10
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ acnqsmod = 0
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ rbodymod = 0
+ mjswgd = 0.95
+ mjswgs = 0.95
+ pvfbsdoff = 0
+ tcjswg = 0.00128
+ keta = -0.21540901
+ pvoff = 2.2423089e-16
+ cdscb = 0
+ cdscd = 0
+ lags = -3.1969346e-8
+ pvsat = 4.7370831e-9
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ wk2we = 0.0
+ pvth0 = 2.4307048999999997e-15
+ lcit = 2.5212768e-10
+ drout = 0.56
+ kt1l = 0
+ paigc = 2.5179991e-18
+ voffl = 0
+ wpdiblc2 = 1.6594883e-9
+ lint = 0
+ lkt1 = -2.2398309e-9
+ lkt2 = -4.7343777e-11
+ weta0 = 4.221971e-8
+ nfactor = 1
+ lmax = 8.833e-8
+ wetab = 1.3144359e-7
+ fprout = 200
+ lmin = 5.233e-8
+ lpclm = -1.0675035e-7
+ xrcrg1 = 12
+ xrcrg2 = 1
+ lpe0 = 6.44e-8
+ lpeb = 0
+ cgidl = 1
+ minv = -0.33
+ lua1 = -2.0580314e-17
+ lub1 = 3.261922e-26
+ luc1 = 9.999327e-18
+ wtvoff = -1.8141864e-9
+ ndep = 1e+18
+ lwlc = 0
+ moin = 5.5538
+ wkvth0we = 0.0
+ nigbacc = 10
+ pbswd = 0.9
+ nigc = 2.291
+ pbsws = 0.9
+ capmod = 2
+ trnqsmod = 0
+ wku0we = 1.5e-11
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ mobmod = 0
+ pdits = 0
+ nigbinv = 2.171
+ cigsd = 0.013281
+ pags = 2.8964227e-14
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ wtvfbsdoff = 0
+ ntox = -1.9260000000000002
+ pcit = -5.430980399999999e-17
+ pclm = 2.5596902
+ rgatemod = 0
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ tnjtsswg = 1
+ ltvfbsdoff = 0
+ phin = 0.15
+ pkt1 = 7.7820041e-17
+ pkt2 = 1.7971063e-15
+ fnoimod = 1
+ tnoia = 0
+ eigbinv = 1.1
+ peta0 = -4.2107701999999996e-15
+ petab = -6.6743123e-15
+ wketa = 8.0928346e-8
+ tpbsw = 0.0025
+ rbdb = 50
+ pua1 = 1.1954606e-22
+ prwb = 0
+ pub1 = -2.033661e-31
+ prwg = 0
+ puc1 = -2.1449333e-23
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ cjswd = 5.457e-11
+ pvag = 2.1
+ cjsws = 5.457e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ rdsw = 200
+ ptvfbsdoff = 0
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ cigbacc = 0.245
+ tnoimod = 0
+ rshg = 14.1
+ scref = 1e-6
+ pigcd = 2.572
+ cigbinv = 0.006
+ aigsd = 0.0063634291
+ lvoff = -2.6816163e-9
+ toxref = 3e-9
+ lvsat = -0.0078314754
+ lvth0 = -2.4372179e-9
+ version = 4.5
+ ijthsfwd = 0.01
+ delta = 0.018814
+ tvfbsdoff = 0.1
+ tempmod = 0
+ laigc = -1.5433256e-11
+ tnom = 25
+ toxe = 2.71e-9
+ toxm = 2.67e-9
+ rnoia = 0
+ rnoib = 0
+ aigbacc = 0.012071
+ ltvoff = 1.2625293e-11
+ pketa = -4.6938441e-15
+ a0 = 3.5386076
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ ngate = 1.7e+20
+ at = 143383.81
+ cf = 7.598099999999999e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.0088402851
+ k3 = -2.5823
+ ijthsrev = 0.01
+ em = 20000000.0
+ ngcon = 1
+ ll = 0
+ lw = 0
+ u0 = 0.0053697056
+ wpclm = -1.0128863e-6
+ w0 = 0
+ ua = -1.1502605e-9
+ ub = 1.2690751e-18
+ uc = -9.619668e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 5.6700000000000005e-9
+ ww = 0
+ xw = 3.4e-9
+ gbmin = 1e-12
+ wags = 9.0067526e-7
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ aigbinv = 0.009974
+ wcit = 2.5843474999999997e-10
+ lku0we = 1.8e-11
+ wvfbsdoff = 0
+ epsrox = 3.9
+ lvfbsdoff = 0
+ voff = -0.11844975
+ acde = 0.5
+ vsat = 219182.19
+ ppdiblc2 = 0
+ rdsmod = 0
+ wint = 0
+ vth0 = -0.34163754
+ igbmod = 1
+ wkt1 = -4.5227706e-9
+ wkt2 = -2.9740529e-8
+ wmax = 9.0026e-6
+ aigc = 0.0067091511
+ wmin = 9.025999999999999e-7
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ pbswgd = 0.8
+ ags = 3.2058772
+ pbswgs = 0.8
+ )

.model pch_ss_15 pmos (
+ level = 54
+ keta = 0.054978601
+ fnoimod = 1
+ pdits = 0
+ eigbinv = 1.1
+ cigsd = 0.013281
+ permod = 1
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 4.182355e-10
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ kt1l = 0
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ lint = 0
+ lkt1 = -1.4608112e-8
+ lkt2 = 1.0752811e-9
+ lmax = 5.233e-8
+ lmin = 4.333e-8
+ voffcv = -0.125
+ wpemod = 1
+ tnoia = 0
+ lpe0 = 6.44e-8
+ lpeb = 0
+ ijthsfwd = 0.01
+ cigbacc = 0.245
+ peta0 = 5.934656900000001e-15
+ petab = -1.9628815e-15
+ minv = -0.33
+ lua1 = -1.9488641e-18
+ lub1 = 6.8003561e-26
+ wketa = -5.4843946e-8
+ luc1 = -2.115524e-18
+ tpbsw = 0.0025
+ ndep = 1e+18
+ tnoimod = 0
+ cjswd = 5.457e-11
+ lwlc = 0
+ cjsws = 5.457e-11
+ moin = 5.5538
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ nigc = 2.291
+ cigbinv = 0.006
+ ijthsrev = 0.01
+ tpbswg = 0.001
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ version = 4.5
+ tempmod = 0
+ ntox = -1.9260000000000002
+ pcit = -6.998464999999996e-18
+ pclm = 1.3082183
+ scref = 1e-6
+ ptvoff = 9.8606268e-17
+ ppdiblc2 = 0
+ pigcd = 2.572
+ aigsd = 0.0063634291
+ waigsd = 1.9051377e-12
+ aigbacc = 0.012071
+ phin = 0.15
+ lvoff = -4.1725981e-9
+ diomod = 1
+ pkt1 = 1.3948109e-14
+ pkt2 = -4.0388508e-15
+ lvsat = 0.00288919592
+ lvth0 = -3.9411155e-9
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.9367000000000001e-10
+ pku0we = 0.0
+ cjswgs = 1.9367000000000001e-10
+ tvfbsdoff = 0.1
+ delta = 0.018814
+ aigbinv = 0.009974
+ laigc = -9.3796225e-12
+ rnoia = 0
+ rnoib = 0
+ rbdb = 50
+ pua1 = -1.9221227e-22
+ prwb = 0
+ pub1 = 2.2863324e-31
+ prwg = 0
+ puc1 = 2.3602641e-23
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ pkvth0we = 0.0
+ rbsb = 50
+ pvag = 2.1
+ mjswgd = 0.95
+ mjswgs = 0.95
+ rdsw = 200
+ pketa = 3.1809489e-15
+ ngate = 1.7e+20
+ ngcon = 1
+ tcjswg = 0.00128
+ wpclm = 1.8421624e-6
+ vfbsdoff = 0.01
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ poxedge = 1
+ paramchk = 1
+ rshg = 14.1
+ binunit = 2
+ ags = 2.6546816
+ cjd = 0.00144022
+ cit = -0.0039626829
+ cjs = 0.00144022
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 4.0349e-9
+ fprout = 200
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ ijthdfwd = 0.01
+ la0 = -1.5436392e-7
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0.0053243403
+ kt1 = -0.063173267
+ kt2 = -0.094912467
+ lk2 = 4.6787193e-9
+ llc = 0
+ tvoff = 0.0053332949
+ lln = 1
+ lu0 = -5.6856188999999995e-11
+ wtvoff = -1.4437583e-9
+ tnom = 25
+ mjd = 0.335
+ mjs = 0.335
+ lua = -3.3837758e-17
+ lub = -4.9508248999999997e-26
+ luc = -2.4014309e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = -3.174587e-14
+ toxe = 2.71e-9
+ toxm = 2.67e-9
+ xjbvd = 1
+ xjbvs = 1
+ nsd = 1e+20
+ pbd = 0.75
+ pat = -5.2399134e-10
+ lk2we = 0.0
+ pbs = 0.75
+ pk2 = 5.1035691e-16
+ pu0 = -9.701894e-17
+ prt = 0
+ pua = -1.0296702e-22
+ pub = 1.2581926e-31
+ puc = 2.16225e-23
+ pud = 0
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ rsh = 15.2
+ wtvfbsdoff = 0
+ tcj = 0.000832
+ ua1 = 5.6955479e-10
+ ub1 = -2.0140988e-18
+ uc1 = 2.5296559e-10
+ ijthdrev = 0.01
+ capmod = 2
+ tpb = 0.0016
+ wa0 = 3.9604044e-7
+ ute = -1
+ wat = 0.00058470362
+ ku0we = -0.0007
+ web = 6628.3
+ wec = -16935.0
+ wk2 = -9.6029938e-9
+ wku0we = 1.5e-11
+ wlc = 0
+ beta0 = 13.32
+ wln = 1
+ wu0 = 7.8023907e-10
+ xgl = -8.2e-9
+ xgw = 0
+ lpdiblc2 = 0
+ wua = 1.5228349e-15
+ wub = -2.3234203999999997e-24
+ leta0 = -2.8797369e-9
+ wuc = -4.6587973e-16
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ letab = 1.0403109e-8
+ ltvfbsdoff = 0
+ mobmod = 0
+ wags = 1.4000585e-6
+ ppclm = -9.0739811e-14
+ wcit = -5.572851699999999e-10
+ voff = -0.092743162
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ acde = 0.5
+ vsat = 34342.667
+ wint = 0
+ vth0 = -0.31570814
+ wkt1 = -2.4366569e-7
+ wkt2 = 7.087942e-8
+ wmax = 9.0026e-6
+ aigc = 0.0066047781
+ wmin = 9.025999999999999e-7
+ njtsswg = 6.489
+ dmcgt = 0
+ lkvth0we = 3e-12
+ tcjsw = 9.34e-5
+ ptvfbsdoff = 0
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ wua1 = 3.9047481e-15
+ wub1 = -4.8164385e-24
+ wuc1 = -5.0052376e-16
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.00081573526
+ pdiblcb = 0
+ bigc = 0.0012521
+ acnqsmod = 0
+ wwlc = 0
+ bigsd = 0.0003327
+ cdsc = 0
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ wvoff = 1.0199556e-9
+ rbodymod = 0
+ cgbo = 0
+ cgdl = 2.799765e-11
+ cgdo = 2.4628259999999997e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 2.799765e-11
+ cgso = 2.4628259999999997e-11
+ cigc = 0.15259
+ wvsat = 0.051609605399999994
+ bigbacc = 0.0054401
+ wvth0 = 3.1849199e-8
+ waigc = 1.173226e-10
+ kvth0we = -0.00022
+ lintnoi = -5e-9
+ lketa = -6.6687589e-9
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ xpart = 1
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ wpdiblc2 = 1.6594883e-9
+ toxref = 3e-9
+ egidl = 0.001
+ k2we = 5e-5
+ dsub = 0.5
+ dtox = 3.91e-10
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ eta0 = 0.2041955
+ etab = -0.27743155
+ ltvoff = -2.3219338e-10
+ wkvth0we = 0.0
+ pvfbsdoff = 0
+ trnqsmod = 0
+ nfactor = 1
+ pvoff = -1.0168765e-16
+ lku0we = 1.8e-11
+ cdscb = 0
+ cdscd = 0
+ epsrox = 3.9
+ pvsat = -2.41941307e-9
+ wk2we = 0.0
+ pvth0 = -2.2190829e-15
+ drout = 0.56
+ paigc = -5.5262052e-18
+ rdsmod = 0
+ igbmod = 1
+ rgatemod = 0
+ voffl = 0
+ tnjtsswg = 1
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ nigbacc = 10
+ weta0 = -1.3270144999999998e-7
+ wetab = 5.0212024e-8
+ pbswgd = 0.8
+ pbswgs = 0.8
+ lpclm = -3.4164983e-8
+ a0 = 2.1782471
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = -44109.368
+ cf = 7.598099999999999e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.015698968
+ k3 = -2.5823
+ em = 20000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.009995586800000001
+ w0 = 0
+ igcmod = 1
+ ua = 3.7489785e-10
+ ub = 2.3417036e-18
+ uc = 4.9437493e-10
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 5.6700000000000005e-9
+ ww = 0
+ xw = 3.4e-9
+ cgidl = 1
+ nigbinv = 2.171
+ pbswd = 0.9
+ pbsws = 0.9
+ )

.model pch_ss_16 pmos (
+ level = 54
+ wpdiblc2 = 1.6594883e-9
+ voffcv = -0.125
+ wpemod = 1
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ bigbacc = 0.0054401
+ tnom = 25
+ kvth0we = -0.00022
+ toxe = 2.71e-9
+ toxm = 2.67e-9
+ bigsd = 0.0003327
+ lintnoi = -5e-9
+ wkvth0we = 0.0
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ wvoff = -9.7608128e-9
+ trnqsmod = 0
+ wvsat = -0.005489889499999999
+ tpbswg = 0.001
+ wvth0 = 1.56900233e-8
+ wags = 3.1454838e-6
+ waigc = -1.1150212e-11
+ wcit = -1.1254199e-9
+ voff = -0.099237323
+ acde = 0.5
+ lketa = 8.2510741e-9
+ ptvoff = -1.3565734e-16
+ xpart = 1
+ waigsd = 2.0479558e-12
+ vsat = 142907.74
+ wint = 0
+ rgatemod = 0
+ vth0 = -0.39088314
+ wkt1 = 3.1251908e-7
+ wkt2 = -1.0928272e-8
+ tnjtsswg = 1
+ wmax = 9.0026e-6
+ aigc = 0.0065575398
+ wmin = 9.025999999999999e-7
+ diomod = 1
+ egidl = 0.001
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.9367000000000001e-10
+ pku0we = 0.0
+ cjswgs = 1.9367000000000001e-10
+ nfactor = 1
+ wua1 = -3.8771176e-15
+ wub1 = 4.6247757e-24
+ wuc1 = 9.3089203e-17
+ bigc = 0.0012521
+ wwlc = 0
+ mjswgd = 0.95
+ mjswgs = 0.95
+ pvfbsdoff = 0
+ cdsc = 0
+ tcjswg = 0.00128
+ cgbo = 0
+ cgdl = 2.799765e-11
+ cgdo = 2.4628259999999997e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 2.799765e-11
+ cgso = 2.4628259999999997e-11
+ cigc = 0.15259
+ nigbacc = 10
+ pvoff = 4.2657e-16
+ cdscb = 0
+ cdscd = 0
+ pvsat = 3.7846031e-10
+ wk2we = 0.0
+ pvth0 = -1.4272744e-15
+ drout = 0.56
+ paigc = 7.6896258e-19
+ nigbinv = 2.171
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ voffl = 0
+ dmdg = 0
+ fprout = 200
+ weta0 = 4.7304045e-9
+ xrcrg1 = 12
+ xrcrg2 = 1
+ wetab = 3.974597e-8
+ wtvfbsdoff = 0
+ lpclm = -2.1829165e-8
+ k2we = 5e-5
+ dsub = 0.5
+ dtox = 3.91e-10
+ ijthsfwd = 0.01
+ wtvoff = 3.3371317e-9
+ cgidl = 1
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ fnoimod = 1
+ ltvfbsdoff = 0
+ eigbinv = 1.1
+ eta0 = 0.11033512
+ etab = -0.14869011
+ capmod = 2
+ pbswd = 0.9
+ pbsws = 0.9
+ ijthsrev = 0.01
+ wku0we = 1.5e-11
+ mobmod = 0
+ pdits = 0
+ cigsd = 0.013281
+ ptvfbsdoff = 0
+ cigbacc = 0.245
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ ppdiblc2 = 0
+ tnoimod = 0
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ laigsd = 7.7486946e-16
+ cigbinv = 0.006
+ tnoia = 0
+ peta0 = -7.995038100000001e-16
+ petab = -1.4500449e-15
+ wketa = 4.9202854e-8
+ version = 4.5
+ tpbsw = 0.0025
+ tempmod = 0
+ cjswd = 5.457e-11
+ pkvth0we = 0.0
+ cjsws = 5.457e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ agidl = 3.2166e-9
+ aigbacc = 0.012071
+ vfbsdoff = 0.01
+ keta = -0.24950779
+ lags = 9.4399385e-8
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = -1.2246200000000013e-12
+ aigbinv = 0.009974
+ kt1l = 0
+ paramchk = 1
+ scref = 1e-6
+ pigcd = 2.572
+ aigsd = 0.0063634133
+ toxref = 3e-9
+ lint = 0
+ lvoff = -3.8543842e-9
+ lkt1 = -1.11161514e-9
+ lkt2 = 4.9336152e-10
+ lmax = 4.333e-8
+ lmin = 3.6e-8
+ lpe0 = 6.44e-8
+ lvsat = -0.0024304684
+ lpeb = 0
+ tvfbsdoff = 0.1
+ lvth0 = -2.57542306e-10
+ ijthdfwd = 0.01
+ delta = 0.018814
+ laigc = -7.0649434e-12
+ minv = -0.33
+ lua1 = -6.8231177e-17
+ lub1 = 7.2428606e-26
+ luc1 = 2.786749e-18
+ poxedge = 1
+ rnoia = 0
+ rnoib = 0
+ ndep = 1e+18
+ ltvoff = -9.8738127e-12
+ lwlc = 0
+ moin = 5.5538
+ binunit = 2
+ pketa = -1.9173443e-15
+ ngate = 1.7e+20
+ nigc = 2.291
+ ijthdrev = 0.01
+ ngcon = 1
+ wpclm = -3.2091624e-7
+ lpdiblc2 = 0
+ gbmin = 1e-12
+ lku0we = 1.8e-11
+ noff = 2.2684
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ epsrox = 3.9
+ ags = 0.72816353
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ cjd = 0.00144022
+ cit = 0.004597740249999999
+ cjs = 0.00144022
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ pags = -8.5525843e-14
+ dlc = 4.0349e-9
+ k3b = 2.1176
+ rdsmod = 0
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ ntox = -1.9260000000000002
+ pcit = 2.0840749999999998e-17
+ pclm = 1.0564669
+ igbmod = 1
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ la0 = -3.7737017e-8
+ jsd = 1.5e-7
+ phin = 0.15
+ jss = 1.5e-7
+ lat = -0.0009151022
+ jtsswgd = 1.75e-7
+ kt1 = -0.33861198
+ kt2 = -0.083036557
+ lk2 = 4.4583258000000006e-9
+ jtsswgs = 1.75e-7
+ llc = 0
+ lln = 1
+ pbswgd = 0.8
+ pbswgs = 0.8
+ lu0 = 1.5817989000000002e-10
+ mjd = 0.335
+ mjs = 0.335
+ lua = 2.9640356e-17
+ lub = 2.9920689e-26
+ luc = -2.5002144e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ lkvth0we = 3e-12
+ njd = 1.02
+ njs = 1.02
+ pa0 = -1.5136929e-14
+ pkt1 = -1.3304944e-14
+ pkt2 = -3.0273858e-17
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 2.5964497e-9
+ pbs = 0.75
+ pk2 = 4.883387e-16
+ igcmod = 1
+ pu0 = -4.5849539e-17
+ prt = 0
+ pua = 8.5912273e-23
+ pub = -1.6837969000000002e-31
+ puc = 8.2880171e-25
+ pud = 0
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 1.9222551e-9
+ ub1 = -2.1044059e-18
+ uc1 = 1.529192e-10
+ tvoff = 0.00079616085
+ tpb = 0.0016
+ wa0 = 5.7082474e-8
+ acnqsmod = 0
+ xjbvd = 1
+ ute = -1
+ wat = -0.063097766
+ xjbvs = 1
+ web = 6628.3
+ wec = -16935.0
+ rbdb = 50
+ wk2 = -9.1536426e-9
+ pua1 = 1.8909915e-22
+ prwb = 0
+ lk2we = 0.0
+ pub1 = -2.3398623999999997e-31
+ prwg = 0
+ puc1 = -5.4843946e-24
+ wlc = 0
+ wln = 1
+ wu0 = -2.6403442e-10
+ xgl = -8.2e-9
+ rbpb = 50
+ rbpd = 50
+ xgw = 0
+ rbps = 50
+ rbsb = 50
+ wua = -2.3318447e-15
+ pvag = 2.1
+ wub = 3.6806403e-24
+ wuc = -4.1518546e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ rdsw = 200
+ rbodymod = 0
+ paigsd = -6.9980875e-21
+ ku0we = -0.0007
+ beta0 = 13.32
+ njtsswg = 6.489
+ leta0 = 1.7194218e-9
+ letab = 4.094779e-9
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ ppclm = 1.5251044e-14
+ permod = 1
+ a0 = -0.20189383
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ ckappad = 0.6
+ at = 83226.192
+ cf = 7.598099999999999e-11
+ ckappas = 0.6
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.01120114
+ k3 = -2.5823
+ em = 20000000.0
+ dlcig = 2.5e-9
+ pdiblc1 = 0
+ pdiblc2 = 0.00081573526
+ ll = 0
+ lw = 0
+ bgidl = 1834800000.0
+ u0 = 0.0056070954
+ w0 = 0
+ pdiblcb = 0
+ ua = -9.2057386e-10
+ ub = 7.207055e-19
+ uc = 5.5311765e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 5.6700000000000005e-9
+ ww = 0
+ xw = 3.4e-9
+ rshg = 14.1
+ )

.model pch_ss_17 pmos (
+ level = 54
+ tpbsw = 0.0025
+ aigbinv = 0.009974
+ eta0 = 0.191845
+ cjswd = 5.457e-11
+ cjsws = 5.457e-11
+ etab = -0.18516667
+ a0 = 2.6112
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ at = 72000
+ cf = 7.598099999999999e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.0045864754
+ k3 = -2.5823
+ em = 20000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.009985966700000001
+ w0 = 0
+ ua = 1.9119717e-10
+ ub = 1.0765761e-18
+ uc = -8.28048e-12
+ ud = 0
+ ijthdrev = 0.01
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 5.6700000000000005e-9
+ ww = 0
+ xw = 3.4e-9
+ tpbswg = 0.001
+ lpdiblc2 = 0
+ ptvoff = 0
+ waigsd = 1.9350626e-12
+ scref = 1e-6
+ poxedge = 1
+ pigcd = 2.572
+ aigsd = 0.0063633642
+ diomod = 1
+ binunit = 2
+ lvoff = 0
+ pditsd = 0
+ lkvth0we = 3e-12
+ pditsl = 0
+ cjswgd = 1.9367000000000001e-10
+ pku0we = 0.0
+ cjswgs = 1.9367000000000001e-10
+ tvfbsdoff = 0.1
+ lvsat = 0.00024
+ lvth0 = -6e-10
+ delta = 0.018814
+ acnqsmod = 0
+ rnoia = 0
+ rnoib = 0
+ mjswgd = 0.95
+ mjswgs = 0.95
+ tcjswg = 0.00128
+ ngate = 1.7e+20
+ rbodymod = 0
+ ags = 0.98525249
+ ngcon = 1
+ wpclm = -5.08417e-8
+ cjd = 0.00144022
+ cit = 5e-6
+ cjs = 0.00144022
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ dlc = 1.0572421799999999e-8
+ k3b = 2.1176
+ dwb = 0
+ keta = -0.016063969
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ gbmin = 1e-12
+ wvfbsdoff = 0
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ lvfbsdoff = 0
+ wtvfbsdoff = 0
+ la0 = 0
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0.001
+ lcit = 0
+ kt1 = -0.18299632
+ lk2 = 4e-10
+ kt2 = -0.042133438
+ llc = 0
+ lln = 1
+ lu0 = 5e-12
+ mjd = 0.335
+ kt1l = 0
+ mjs = 0.335
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 0
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ ltvfbsdoff = 0
+ pk2 = 0
+ wpdiblc2 = -1.7580235e-10
+ fprout = 200
+ pu0 = 0
+ prt = 0
+ pud = 0
+ lint = 6.5375218e-9
+ xrcrg1 = 12
+ xrcrg2 = 1
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 1.45515e-9
+ ub1 = -1.5029257e-18
+ uc1 = -4.3667733e-11
+ lkt1 = -1e-9
+ lmax = 2.001e-5
+ tpb = 0.0016
+ wa0 = 2.308488e-7
+ lmin = 8.99743e-6
+ ute = -0.96728333
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 1.3953799e-9
+ njtsswg = 6.489
+ lpe0 = 6.44e-8
+ wlc = 0
+ wln = 1
+ wu0 = 2.7482e-12
+ xgl = -8.2e-9
+ lpeb = 0
+ xgw = 0
+ wua = -1.5682603e-16
+ wub = 3.5681818e-26
+ wuc = 4.8873989e-18
+ wud = 0
+ wtvoff = -7.2458121e-11
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ tvoff = 0.0025973351
+ minv = -0.33
+ xjbvd = 1
+ xjbvs = 1
+ ckappad = 0.6
+ ckappas = 0.6
+ lk2we = 0.0
+ ndep = 1e+18
+ pdiblc1 = 0
+ pdiblc2 = 0.0032290423
+ pdiblcb = 0
+ lwlc = 0
+ ptvfbsdoff = 0
+ capmod = 2
+ wkvth0we = 0.0
+ moin = 5.5538
+ wku0we = 1.5e-11
+ nigc = 2.291
+ trnqsmod = 0
+ mobmod = 0
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = -5e-10
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ bigbacc = 0.0054401
+ ppclm = 0
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ kvth0we = -0.00022
+ ntox = -1.9260000000000002
+ pcit = 0
+ pclm = 1.2411167
+ rgatemod = 0
+ lintnoi = -5e-9
+ tnjtsswg = 1
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ phin = 0.15
+ vtsswgs = 1.1
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ pkt1 = 0
+ bigsd = 0.0003327
+ rbdb = 50
+ prwb = 0
+ prwg = 0
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ rdsw = 200
+ wvoff = 3.276885e-9
+ wvsat = -0.017628054
+ wvth0 = -1.7405743999999999e-9
+ waigc = -7.2361068e-12
+ nfactor = 1
+ lketa = 0
+ rshg = 14.1
+ xpart = 1
+ toxref = 3e-9
+ egidl = 0.001
+ nigbacc = 10
+ ijthsfwd = 0.01
+ tnom = 25
+ ltvoff = 0
+ toxe = 2.71e-9
+ toxm = 2.67e-9
+ pvfbsdoff = 0
+ nigbinv = 2.171
+ ijthsrev = 0.01
+ lku0we = 1.8e-11
+ pvoff = 2.5e-17
+ epsrox = 3.9
+ wags = -3.1938756e-8
+ cdscb = 0
+ cdscd = 0
+ pvsat = -5e-11
+ wk2we = 0.0
+ rdsmod = 0
+ pvth0 = -7e-17
+ fnoimod = 1
+ drout = 0.56
+ voff = -0.10917042
+ igbmod = 1
+ acde = 0.5
+ eigbinv = 1.1
+ ppdiblc2 = 0
+ vsat = 129757.01
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ wint = 0
+ voffl = 0
+ vth0 = -0.41024647000000003
+ wkt1 = 1.4804073e-9
+ wkt2 = -8.3218931e-9
+ pbswgd = 0.8
+ pbswgs = 0.8
+ wmax = 9.025999999999999e-7
+ aigc = 0.0068422292
+ wmin = 5.426e-7
+ weta0 = -2.4521569999999998e-8
+ wetab = 1.3741e-8
+ igcmod = 1
+ lpclm = 0
+ wua1 = -5.289391e-16
+ wub1 = 6.5622425e-25
+ wuc1 = 2.3227786e-17
+ cgidl = 1
+ bigc = 0.0012521
+ wute = -1.003093e-7
+ cigbacc = 0.245
+ wwlc = 0
+ pkvth0we = 0.0
+ cdsc = 0
+ tnoimod = 0
+ pbswd = 0.9
+ pbsws = 0.9
+ cgbo = 0
+ cgdl = 2.799765e-11
+ cgdo = 2.4628259999999997e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 2.799765e-11
+ cgso = 2.4628259999999997e-11
+ cigc = 0.15259
+ vfbsdoff = 0.01
+ cigbinv = 0.006
+ permod = 1
+ pdits = 0
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ paramchk = 1
+ version = 4.5
+ tempmod = 0
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ voffcv = -0.125
+ wpemod = 1
+ aigbacc = 0.012071
+ k2we = 5e-5
+ tnoia = 0
+ dsub = 0.5
+ dtox = 3.91e-10
+ ijthdfwd = 0.01
+ peta0 = -1.5e-17
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ wketa = -3.7023239e-9
+ )

.model pch_ss_18 pmos (
+ level = 54
+ waigc = -9.2878513e-12
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ nigbacc = 10
+ ptvoff = 6.0745993e-16
+ pags = -1.6587566e-14
+ waigsd = 1.93751e-12
+ lketa = -8.0782883e-8
+ ntox = -1.9260000000000002
+ pcit = 0
+ pclm = 1.2411167
+ xpart = 1
+ ppdiblc2 = 2.0750737e-15
+ diomod = 1
+ nigbinv = 2.171
+ phin = 0.15
+ egidl = 0.001
+ pditsd = 0
+ pditsl = 0
+ a0 = 2.6572474
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ cjswgd = 1.9367000000000001e-10
+ pku0we = 0.0
+ cjswgs = 1.9367000000000001e-10
+ at = 72000
+ cf = 7.598099999999999e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.0050849127
+ k3 = -2.5823
+ em = 20000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.0098657581
+ pkt1 = 7.4878862e-15
+ pkt2 = 7.624365e-15
+ w0 = 0
+ ua = 1.8022848e-10
+ ub = 1.0497212e-18
+ uc = -5.9216956e-12
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 5.6700000000000005e-9
+ ww = 0
+ xw = 3.4e-9
+ mjswgd = 0.95
+ mjswgs = 0.95
+ rbdb = 50
+ pua1 = 3.0135942e-22
+ prwb = 0
+ pub1 = -6.7644414e-31
+ prwg = 0
+ fnoimod = 1
+ puc1 = -4.7294542e-23
+ pvfbsdoff = 0
+ wtvfbsdoff = 0
+ tcjswg = 0.00128
+ pkvth0we = 0.0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ eigbinv = 1.1
+ pute = 3.5290383e-14
+ rdsw = 200
+ ltvfbsdoff = 0
+ vfbsdoff = 0.01
+ pvoff = 8.2387382e-16
+ cdscb = 0
+ cdscd = 0
+ pvsat = -5e-11
+ wk2we = 0.0
+ pvth0 = -1.2364923999999999e-15
+ drout = 0.56
+ paramchk = 1
+ paigc = 1.8445184e-17
+ rshg = 14.1
+ cigbacc = 0.245
+ fprout = 200
+ voffl = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ tnoimod = 0
+ ptvfbsdoff = 0
+ weta0 = -2.4521569999999998e-8
+ wetab = 1.3741e-8
+ lpclm = 0
+ wtvoff = -1.4002875e-10
+ cigbinv = 0.006
+ ijthdfwd = 0.01
+ cgidl = 1
+ tnom = 25
+ toxe = 2.71e-9
+ toxm = 2.67e-9
+ capmod = 2
+ version = 4.5
+ wku0we = 1.5e-11
+ tempmod = 0
+ pbswd = 0.9
+ pbsws = 0.9
+ ijthdrev = 0.01
+ mobmod = 0
+ lpdiblc2 = 3.0626629e-9
+ aigbacc = 0.012071
+ wags = -3.0093643e-8
+ pdits = 0
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ voff = -0.10728654
+ acde = 0.5
+ vsat = 129757.01
+ aigbinv = 0.009974
+ wint = 0
+ vth0 = -0.40917796
+ laigsd = 5.7445099e-14
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ wkt1 = 6.4749443e-10
+ wkt2 = -9.1699871e-9
+ wmax = 9.025999999999999e-7
+ aigc = 0.0068507406
+ wmin = 5.426e-7
+ lkvth0we = 3e-12
+ tnoia = 0
+ peta0 = -1.5e-17
+ wua1 = -5.6246072e-16
+ wub1 = 7.3146831e-25
+ wuc1 = 2.8488581e-17
+ wketa = -8.2059163e-9
+ bigc = 0.0012521
+ wute = -1.0423482e-7
+ acnqsmod = 0
+ tpbsw = 0.0025
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ wwlc = 0
+ cjswd = 5.457e-11
+ cjsws = 5.457e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ poxedge = 1
+ cdsc = 0
+ rbodymod = 0
+ cgbo = 0
+ cgdl = 2.799765e-11
+ cgdo = 2.4628259999999997e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 2.799765e-11
+ cgso = 2.4628259999999997e-11
+ cigc = 0.15259
+ binunit = 2
+ toxref = 3e-9
+ scref = 1e-6
+ pigcd = 2.572
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ wpdiblc2 = -4.0662257e-10
+ aigsd = 0.0063633578
+ dmdg = 0
+ lvoff = -1.6936099e-8
+ tvfbsdoff = 0.1
+ k2we = 5e-5
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ lvsat = 0.00024
+ lvth0 = -1.02058678e-8
+ dsub = 0.5
+ dtox = 3.91e-10
+ delta = 0.018814
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ laigc = -7.651731e-11
+ ltvoff = -1.5996918e-9
+ ags = 0.95300429
+ rnoia = 0
+ rnoib = 0
+ cjd = 0.00144022
+ cit = 5e-6
+ cjs = 0.00144022
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 1.0572421799999999e-8
+ k3b = 2.1176
+ eta0 = 0.191845
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ etab = -0.18516667
+ dwj = 0
+ wkvth0we = 0.0
+ pketa = 4.0487295e-14
+ ngate = 1.7e+20
+ ngcon = 1
+ wpclm = -5.08417e-8
+ trnqsmod = 0
+ la0 = -4.1396638e-7
+ lku0we = 1.8e-11
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0.001
+ kt1 = -0.17852273
+ kt2 = -0.039741464
+ lk2 = 4.8809517e-9
+ llc = 0
+ lln = 1
+ epsrox = 3.9
+ lu0 = 1.0856753e-9
+ mjd = 0.335
+ wvfbsdoff = 0
+ mjs = 0.335
+ lua = 9.8608496e-17
+ lub = 2.4142536e-25
+ luc = -2.1205472e-17
+ lud = 0
+ gbmin = 1e-12
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ lvfbsdoff = 0
+ njd = 1.02
+ njs = 1.02
+ pa0 = -1.9681175e-13
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ pk2 = -1.7465146e-15
+ njtsswg = 6.489
+ pu0 = -2.7146448e-18
+ rdsmod = 0
+ prt = 0
+ pua = -5.0852536e-23
+ pub = 3.3773548e-32
+ puc = 2.1258791e-23
+ pud = 0
+ igbmod = 1
+ xtsswgd = 0.32
+ rsh = 15.2
+ xtsswgs = 0.32
+ tcj = 0.000832
+ ua1 = 1.3709274e-9
+ ub1 = -1.4287011e-18
+ uc1 = -6.3574807e-11
+ tpb = 0.0016
+ wa0 = 2.527411e-7
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ ute = -0.97152091
+ ckappad = 0.6
+ ckappas = 0.6
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 1.5896529e-9
+ wlc = 0
+ rgatemod = 0
+ wln = 1
+ pdiblc1 = 0
+ pdiblc2 = 0.0028883679
+ wu0 = 3.0501627e-12
+ xgl = -8.2e-9
+ xgw = 0
+ pbswgd = 0.8
+ pdiblcb = 0
+ wua = -1.5116947e-16
+ pbswgs = 0.8
+ wub = 3.1925028e-26
+ wuc = 2.5226836e-18
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ tnjtsswg = 1
+ igcmod = 1
+ tvoff = 0.0027752763
+ bigbacc = 0.0054401
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ kvth0we = -0.00022
+ paigsd = -2.2002196e-20
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ ku0we = -0.0007
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ beta0 = 13.32
+ leta0 = -5e-10
+ keta = -0.0070781088
+ permod = 1
+ ppclm = 0
+ lags = 2.8991134e-7
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ dlcig = 2.5e-9
+ lcit = 0
+ bgidl = 1834800000.0
+ kt1l = 0
+ voffcv = -0.125
+ wpemod = 1
+ lint = 6.5375218e-9
+ lkt1 = -4.1217527000000004e-8
+ lkt2 = -2.1503841e-8
+ dmcgt = 0
+ lmax = 8.99743e-6
+ tcjsw = 9.34e-5
+ lmin = 8.974099999999999e-7
+ lpe0 = 6.44e-8
+ lpeb = 0
+ ijthsfwd = 0.01
+ minv = -0.33
+ lua1 = 7.5716104e-16
+ lub1 = -6.6727951e-25
+ luc1 = 1.7896459e-16
+ nfactor = 1
+ bigsd = 0.0003327
+ ndep = 1e+18
+ lute = 3.8095772e-8
+ lwlc = 0
+ moin = 5.5538
+ wvoff = 3.1880225e-9
+ tpbswg = 0.001
+ ijthsrev = 0.01
+ nigc = 2.291
+ wvsat = -0.017628054
+ wvth0 = -1.6108199999999998e-9
+ noff = 2.2684
+ )

.model pch_ss_19 pmos (
+ level = 54
+ cjd = 0.00144022
+ cit = -8.7888889e-5
+ cjs = 0.00144022
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ lvsat = 0.00024
+ dlc = 1.0572421799999999e-8
+ k3b = 2.1176
+ lvth0 = -7.6657388e-10
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ ltvfbsdoff = 0
+ wua1 = -6.1430214e-16
+ wub1 = 1.1920544e-25
+ delta = 0.018814
+ wuc1 = -4.9561039e-17
+ laigc = -1.8208261e-11
+ mjswgd = 0.95
+ mjswgs = 0.95
+ njtsswg = 6.489
+ bigc = 0.0012521
+ wute = -1.2773023e-7
+ rnoia = 0
+ rnoib = 0
+ la0 = -9.6086602e-7
+ wwlc = 0
+ tcjswg = 0.00128
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0.001
+ kt1 = -0.20738899
+ kt2 = -0.065812764
+ lk2 = 1.6919589000000001e-10
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ llc = 0
+ lln = 1
+ lu0 = -1.5232407999999998e-9
+ mjd = 0.335
+ mjs = 0.335
+ lua = -3.205013e-16
+ lub = -3.7552526e-26
+ luc = 5.1848161e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 2.9499704e-13
+ pketa = -2.8529622e-14
+ ckappad = 0.6
+ cdsc = 0
+ ckappas = 0.6
+ ngate = 1.7e+20
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ pk2 = 8.8602334e-16
+ pdiblc1 = 0
+ pdiblc2 = -8.9657994e-6
+ cgbo = 0
+ cgdl = 2.799765e-11
+ cgdo = 2.4628259999999997e-11
+ xtid = 3
+ ngcon = 1
+ xtis = 3
+ pdiblcb = 0
+ pu0 = 4.0536683e-16
+ wpclm = -5.08417e-8
+ prt = 0
+ pua = 3.1718399e-23
+ pub = 9.4535502e-32
+ puc = -3.7711192e-23
+ pud = 0
+ cgsl = 2.799765e-11
+ cgso = 2.4628259999999997e-11
+ cigc = 0.15259
+ rsh = 15.2
+ wvfbsdoff = 0
+ tcj = 0.000832
+ ua1 = 2.985915e-9
+ ub1 = -2.7037422e-18
+ uc1 = 1.5248758e-10
+ lvfbsdoff = 0
+ gbmin = 1e-12
+ tpb = 0.0016
+ wa0 = -2.9985305e-7
+ jswgd = 3.69e-13
+ ptvfbsdoff = 0
+ jswgs = 3.69e-13
+ ute = -0.85901741
+ web = 6628.3
+ wec = -16935.0
+ wk2 = -1.3682549e-9
+ a0 = 3.2717414
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ wlc = 0
+ wln = 1
+ wu0 = -4.5546835e-10
+ at = 72000
+ cf = 7.598099999999999e-11
+ xgl = -8.2e-9
+ ef = 1.15
+ k1 = 0.30425
+ k2 = 0.00020919492
+ xgw = 0
+ k3 = -2.5823
+ em = 20000000.0
+ wua = -2.439458e-16
+ wub = -3.6346832e-26
+ wuc = 6.8781092e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ ll = 0
+ lw = 0
+ u0 = 0.012797124
+ w0 = 0
+ ua = 6.5113837e-10
+ ub = 1.3631795e-18
+ uc = -8.8004429e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 5.6700000000000005e-9
+ ww = 0
+ xw = 3.4e-9
+ bigbacc = 0.0054401
+ fprout = 200
+ xrcrg1 = 12
+ xrcrg2 = 1
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ kvth0we = -0.00022
+ lintnoi = -5e-9
+ wtvoff = 9.9743807e-10
+ bigbinv = 0.00149
+ k2we = 5e-5
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ dsub = 0.5
+ dtox = 3.91e-10
+ ijthsfwd = 0.01
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ tvoff = 0.00044287651
+ capmod = 2
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ wku0we = 1.5e-11
+ eta0 = 0.191845
+ etab = -0.18516667
+ mobmod = 0
+ ijthsrev = 0.01
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = -5e-10
+ ppclm = 0
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ nfactor = 1
+ laigsd = -3.6354984e-15
+ ppdiblc2 = -2.7249029e-15
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ nigbacc = 10
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ bigsd = 0.0003327
+ pkvth0we = 0.0
+ wvoff = 1.2743983e-8
+ nigbinv = 2.171
+ wvsat = -0.017628054
+ vfbsdoff = 0.01
+ wvth0 = -3.53071142e-9
+ keta = -0.13767457
+ waigc = 2.7297355e-11
+ lags = 8.1183869e-8
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 8.2671111e-11
+ toxref = 3e-9
+ paramchk = 1
+ lketa = 3.5447968e-8
+ kt1l = 0
+ xpart = 1
+ fnoimod = 1
+ eigbinv = 1.1
+ lint = 6.5375218e-9
+ egidl = 0.001
+ lkt1 = -1.5526561e-8
+ lkt2 = 1.6996159e-9
+ lmax = 8.974099999999999e-7
+ lmin = 4.4741e-7
+ lpe0 = 6.44e-8
+ lpeb = 0
+ ijthdfwd = 0.01
+ ltvoff = 4.7614406e-10
+ minv = -0.33
+ lua1 = -6.8017788e-16
+ lub1 = 4.6750711e-25
+ luc1 = -1.3330934e-17
+ pvfbsdoff = 0
+ ndep = 1e+18
+ lute = -6.2032341e-8
+ lwlc = 0
+ moin = 5.5538
+ cigbacc = 0.245
+ ijthdrev = 0.01
+ nigc = 2.291
+ lku0we = 1.8e-11
+ epsrox = 3.9
+ tnoimod = 0
+ lpdiblc2 = 5.64129e-9
+ pvoff = -7.6809313e-15
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ rdsmod = 0
+ cdscb = 0
+ cdscd = 0
+ cigbinv = 0.006
+ igbmod = 1
+ pvsat = -5e-11
+ wk2we = 0.0
+ pvth0 = 4.7221102e-16
+ drout = 0.56
+ pags = 2.5130854e-13
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ paigc = -1.411565e-17
+ ntox = -1.9260000000000002
+ pcit = 0
+ pclm = 1.2411167
+ pbswgd = 0.8
+ pbswgs = 0.8
+ voffl = 0
+ version = 4.5
+ igcmod = 1
+ phin = 0.15
+ tempmod = 0
+ weta0 = -2.4521569999999998e-8
+ wetab = 1.3741e-8
+ lkvth0we = 3e-12
+ lpclm = 0
+ pkt1 = -4.6411548e-15
+ pkt2 = -3.0623252e-15
+ aigbacc = 0.012071
+ cgidl = 1
+ acnqsmod = 0
+ rbdb = 50
+ pua1 = 3.4749829e-22
+ prwb = 0
+ pub1 = -1.3153018e-31
+ prwg = 0
+ puc1 = 2.216962e-23
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ paigsd = 1.9849821e-21
+ rbsb = 50
+ pvag = 2.1
+ pute = 5.6201301e-14
+ rdsw = 200
+ rbodymod = 0
+ pbswd = 0.9
+ pbsws = 0.9
+ aigbinv = 0.009974
+ permod = 1
+ pdits = 0
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ rshg = 14.1
+ voffcv = -0.125
+ wpemod = 1
+ wpdiblc2 = 4.9866096e-9
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ poxedge = 1
+ tnoia = 0
+ binunit = 2
+ peta0 = -1.5e-17
+ wketa = 6.9341182e-8
+ tnom = 25
+ tpbsw = 0.0025
+ toxe = 2.71e-9
+ toxm = 2.67e-9
+ cjswd = 5.457e-11
+ cjsws = 5.457e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ wkvth0we = 0.0
+ agidl = 3.2166e-9
+ tpbswg = 0.001
+ trnqsmod = 0
+ wags = -3.311005e-7
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ ptvoff = -4.0488554e-16
+ waigsd = 1.9105581e-12
+ voff = -0.13228318
+ acde = 0.5
+ scref = 1e-6
+ diomod = 1
+ vsat = 129757.01
+ pigcd = 2.572
+ rgatemod = 0
+ wint = 0
+ aigsd = 0.0063634264
+ vth0 = -0.41978391000000004
+ tnjtsswg = 1
+ wkt1 = 1.4275631e-8
+ wkt2 = 2.8375299e-9
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.9367000000000001e-10
+ pku0we = 0.0
+ wmax = 9.025999999999999e-7
+ wtvfbsdoff = 0
+ cjswgs = 1.9367000000000001e-10
+ aigc = 0.0067852248
+ lvoff = 5.3109112e-9
+ wmin = 5.426e-7
+ ags = 1.1875295
+ tvfbsdoff = 0.1
+ )

.model pch_ss_20 pmos (
+ level = 54
+ cjd = 0.00144022
+ cit = -0.00041212495
+ cjs = 0.00144022
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ lvsat = 0.00024
+ dlc = 1.38228675e-8
+ k3b = 2.1176
+ lvth0 = 5.9054743e-9
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ ltvfbsdoff = 0
+ wua1 = 2.4012676e-16
+ wub1 = -6.2487918e-26
+ delta = 0.018814
+ wuc1 = -3.9943707e-17
+ laigc = -2.2400472e-11
+ mjswgd = 0.95
+ mjswgs = 0.95
+ njtsswg = 6.489
+ bigc = 0.0012521
+ rnoia = 0
+ rnoib = 0
+ la0 = -7.2511148e-8
+ wwlc = 0
+ tcjswg = 0.00128
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0.001
+ kt1 = -0.20886849
+ kt2 = -0.049681978
+ lk2 = 1.6117426e-9
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ llc = -1.18e-13
+ lln = 0.7
+ lu0 = -4.7595715e-10
+ mjd = 0.335
+ mjs = 0.335
+ lua = -5.9775833e-17
+ lub = -8.2990392e-26
+ luc = -8.4878869e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = -2.0868237e-13
+ pketa = -1.8963071e-15
+ ckappad = 0.6
+ cdsc = 0
+ ckappas = 0.6
+ ngate = 1.7e+20
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ pk2 = -3.6576402e-16
+ pdiblc1 = 0
+ pdiblc2 = 0.01788848
+ cgbo = 0
+ cgdl = 2.799765e-11
+ cgdo = 2.4628259999999997e-11
+ xtid = 3
+ ngcon = 1
+ xtis = 3
+ pdiblcb = 0
+ pu0 = -2.2283222e-17
+ wpclm = -5.08417e-8
+ prt = 0
+ pua = -3.7414239e-23
+ pub = 6.4271496e-32
+ puc = -3.5764571e-25
+ pud = 0
+ cgsl = 2.799765e-11
+ cgso = 2.4628259999999997e-11
+ cigc = 0.15259
+ rsh = 15.2
+ wvfbsdoff = 0
+ tcj = 0.000832
+ ua1 = 1.3271195e-9
+ ub1 = -1.4620758e-18
+ uc1 = 1.6497662e-10
+ lvfbsdoff = 0
+ gbmin = 1e-12
+ tpb = 0.0016
+ wa0 = 8.4487289e-7
+ jswgd = 3.69e-13
+ ptvfbsdoff = 0
+ jswgs = 3.69e-13
+ ute = -1
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 1.4767164e-9
+ a0 = 1.2527531
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ wlc = 0
+ wln = 1
+ wu0 = 5.1646359e-10
+ at = 72000
+ cf = 7.598099999999999e-11
+ xgl = -8.2e-9
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.0030693202
+ xgw = 0
+ k3 = -2.5823
+ em = 20000000.0
+ wua = -8.6826164e-17
+ wub = 3.2435001e-26
+ wuc = -1.6113333e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ ll = -1.18e-13
+ lw = 0
+ u0 = 0.010416934000000001
+ w0 = 0
+ ua = 5.8580479e-11
+ ub = 1.4664474e-18
+ uc = 4.9122952e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 5.6700000000000005e-9
+ ww = 0
+ xw = 3.4e-9
+ bigbacc = 0.0054401
+ fprout = 200
+ xrcrg1 = 12
+ xrcrg2 = 1
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ kvth0we = -0.00022
+ lintnoi = -5e-9
+ wtvoff = -3.604609e-11
+ bigbinv = 0.00149
+ k2we = 5e-5
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ dsub = 0.5
+ dtox = 3.91e-10
+ ijthsfwd = 0.01
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ tvoff = 0.0020688013
+ capmod = 2
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ wku0we = 1.5e-11
+ eta0 = 0.191845
+ etab = -0.18516667
+ mobmod = 0
+ ijthsrev = 0.01
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = -5e-10
+ ppclm = 0
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ nfactor = 1
+ ppdiblc2 = 1.0915468e-15
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ nigbacc = 10
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ bigsd = 0.0003327
+ pkvth0we = 0.0
+ wvoff = -5.0330429e-9
+ nigbinv = 2.171
+ wvsat = -0.017628054
+ vfbsdoff = 0.01
+ wvth0 = 1.6926608000000005e-9
+ keta = -0.023696099
+ waigc = -1.2459534e-12
+ lags = 6.5053339e-7
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 2.2533498e-10
+ toxref = 3e-9
+ paramchk = 1
+ lketa = -1.4702559e-8
+ kt1l = 0
+ xpart = 1
+ fnoimod = 1
+ eigbinv = 1.1
+ lint = 9.7879675e-9
+ egidl = 0.001
+ lkt1 = -1.4875579e-8
+ lkt2 = -5.3979298e-9
+ lmax = 4.4741e-7
+ lmin = 2.1410000000000002e-7
+ lpe0 = 6.44e-8
+ lpeb = 0
+ ijthdfwd = 0.01
+ ltvoff = -2.3926284e-10
+ minv = -0.33
+ lua1 = 4.9692128e-17
+ lub1 = -7.8826099e-26
+ luc1 = -1.8826114e-17
+ pvfbsdoff = 0
+ ndep = 1e+18
+ lwlc = 0
+ moin = 5.5538
+ cigbacc = 0.245
+ ijthdrev = 0.01
+ nigc = 2.291
+ lku0we = 1.8e-11
+ epsrox = 3.9
+ tnoimod = 0
+ lpdiblc2 = -2.233586e-9
+ pvoff = 1.4096021e-16
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ rdsmod = 0
+ cdscb = 0
+ cdscd = 0
+ cigbinv = 0.006
+ igbmod = 1
+ pvsat = -5e-11
+ wk2we = 0.0
+ pvth0 = -1.8260727e-15
+ drout = 0.56
+ pags = 1.3163813e-13
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ paigc = -1.5565945e-18
+ ntox = -1.9260000000000002
+ pcit = -2.0500564e-17
+ pclm = 1.2411167
+ pbswgd = 0.8
+ pbswgs = 0.8
+ voffl = 0
+ version = 4.5
+ igcmod = 1
+ phin = 0.15
+ tempmod = 0
+ weta0 = -2.4521569999999998e-8
+ wetab = 1.3741e-8
+ lkvth0we = 3e-12
+ lpclm = 0
+ pkt1 = 1.1573276e-15
+ pkt2 = 6.9635068e-17
+ aigbacc = 0.012071
+ cgidl = 1
+ acnqsmod = 0
+ rbdb = 50
+ pua1 = -2.8450432e-23
+ prwb = 0
+ pub1 = -5.1585101e-32
+ prwg = 0
+ puc1 = 1.7937993e-23
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ rdsw = 200
+ rbodymod = 0
+ pbswd = 0.9
+ pbsws = 0.9
+ aigbinv = 0.009974
+ permod = 1
+ pdits = 0
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ rshg = 14.1
+ voffcv = -0.125
+ wpemod = 1
+ wpdiblc2 = -3.6871397e-9
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ poxedge = 1
+ tnoia = 0
+ binunit = 2
+ peta0 = -1.5e-17
+ wketa = 8.8109206e-9
+ tnom = 25
+ tpbsw = 0.0025
+ toxe = 2.71e-9
+ toxm = 2.67e-9
+ cjswd = 5.457e-11
+ cjsws = 5.457e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ wkvth0we = 0.0
+ agidl = 3.2166e-9
+ tpbswg = 0.001
+ trnqsmod = 0
+ wags = -5.9122303e-8
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ ptvoff = 4.9847489e-17
+ wcit = 4.6592191e-11
+ waigsd = 1.9150694e-12
+ voff = -0.10909205
+ acde = 0.5
+ scref = 1e-6
+ diomod = 1
+ vsat = 129757.01
+ pigcd = 2.572
+ rgatemod = 0
+ wint = 0
+ aigsd = 0.0063634182
+ vth0 = -0.43494766
+ tnjtsswg = 1
+ wkt1 = 1.0972613e-9
+ wkt2 = -4.2805615e-9
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.9367000000000001e-10
+ pku0we = 0.0
+ wmax = 9.025999999999999e-7
+ wtvfbsdoff = 0
+ cjswgs = 1.9367000000000001e-10
+ aigc = 0.0067947526
+ lvoff = -4.893186e-9
+ wmin = 5.426e-7
+ ags = -0.10644665
+ tvfbsdoff = 0.1
+ )

.model pch_ss_21 pmos (
+ level = 54
+ rbodymod = 0
+ version = 4.5
+ tempmod = 0
+ keta = -0.074839654
+ pvoff = 3.047289e-16
+ cdscb = 0
+ cdscd = 0
+ lags = 2.5597727e-7
+ pvsat = -5e-11
+ aigbacc = 0.012071
+ wk2we = 0.0
+ pvth0 = 3.5710493999999997e-16
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ drout = 0.56
+ fprout = 200
+ lcit = 1.4712816e-10
+ kt1l = 0
+ paigc = 3.3660127e-18
+ xrcrg1 = 12
+ xrcrg2 = 1
+ voffl = 0
+ wpdiblc2 = 2.1803424e-9
+ lint = 9.7879675e-9
+ weta0 = -2.4521569999999998e-8
+ wtvoff = -4.3702924e-10
+ aigbinv = 0.009974
+ wetab = 1.3741e-8
+ lkt1 = -7.1643470999999995e-9
+ lkt2 = -3.8990903e-9
+ lmax = 2.1410000000000002e-7
+ lpclm = 5.4900145e-8
+ lmin = 8.833e-8
+ lpe0 = 6.44e-8
+ lpeb = 0
+ cgidl = 1
+ minv = -0.33
+ capmod = 2
+ lua1 = -2.9544713e-16
+ lub1 = 3.7855773e-25
+ luc1 = 4.6029572e-17
+ wku0we = 1.5e-11
+ a0 = 0.98313605
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ ndep = 1e+18
+ at = 41320.114
+ cf = 7.598099999999999e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.016096302
+ k3 = -2.5823
+ em = 20000000.0
+ ll = -1.18e-13
+ lwlc = 0
+ lw = 0
+ u0 = 0.008966993000000001
+ mobmod = 0
+ w0 = 0
+ wkvth0we = 0.0
+ ua = 2.7312462e-10
+ ub = 6.1180894e-19
+ uc = 6.0007215e-11
+ ud = 0
+ moin = 5.5538
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 5.6700000000000005e-9
+ ww = 0
+ xw = 3.4e-9
+ pbswd = 0.9
+ pbsws = 0.9
+ nigc = 2.291
+ trnqsmod = 0
+ poxedge = 1
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ binunit = 2
+ pdits = 0
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ pags = -1.3976359e-13
+ ntox = -1.9260000000000002
+ pcit = -3.638512e-17
+ pclm = 0.98092641
+ rgatemod = 0
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ tnjtsswg = 1
+ phin = 0.15
+ pkt1 = 1.542035e-15
+ pkt2 = 2.2793112e-15
+ tnoia = 0
+ peta0 = -1.5e-17
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ wketa = -2.2984762e-8
+ tpbsw = 0.0025
+ rbdb = 50
+ pua1 = 7.9342593e-23
+ prwb = 0
+ pub1 = -9.194958e-32
+ prwg = 0
+ puc1 = -2.9723056e-23
+ cjswd = 5.457e-11
+ cjsws = 5.457e-11
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ mjswd = 0.01
+ rbsb = 50
+ pvag = 2.1
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ rdsw = 200
+ toxref = 3e-9
+ njtsswg = 6.489
+ ags = 1.7634876
+ scref = 1e-6
+ rshg = 14.1
+ cjd = 0.00144022
+ cit = -4.1476524e-5
+ cjs = 0.00144022
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ xtsswgd = 0.32
+ pigcd = 2.572
+ xtsswgs = 0.32
+ dlc = 1.38228675e-8
+ aigsd = 0.0063634182
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ tvfbsdoff = 0.1
+ ckappad = 0.6
+ ckappas = 0.6
+ lvoff = -2.4249846e-9
+ pdiblc1 = 0
+ pdiblc2 = 0.011594472
+ pdiblcb = 0
+ la0 = -1.5621959e-8
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0.007473456
+ lvsat = 0.00024
+ kt1 = -0.24541461
+ kt2 = -0.056785482
+ lk2 = 4.360422800000001e-9
+ llc = -1.18e-13
+ lvth0 = 3.3839767000000003e-9
+ lln = 0.7
+ ltvoff = -2.3342435e-10
+ lu0 = -1.7001950999999999e-10
+ mjd = 0.335
+ mjs = 0.335
+ lua = -1.0504465e-16
+ ijthsfwd = 0.01
+ lub = 9.7338322e-26
+ luc = -1.0784466e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ delta = 0.018814
+ pa0 = -2.5809676e-14
+ nsd = 1e+20
+ laigc = -2.5435198e-11
+ pbd = 0.75
+ pat = -8.1994638e-9
+ pbs = 0.75
+ pk2 = 1.2451684e-16
+ tnom = 25
+ pu0 = -7.9199366e-18
+ prt = 0
+ pua = 5.00917e-23
+ pub = -8.1076857e-32
+ puc = 8.6464743e-24
+ pud = 0
+ rnoia = 0
+ rnoib = 0
+ toxe = 2.71e-9
+ toxm = 2.67e-9
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 2.9628506e-9
+ ub1 = -3.6297717e-18
+ uc1 = -1.423963e-10
+ bigbacc = 0.0054401
+ tpb = 0.0016
+ wa0 = -2.1822352e-8
+ pketa = 4.8125819e-15
+ ute = -1
+ wat = 0.038860018
+ ngate = 1.7e+20
+ web = 6628.3
+ wec = -16935.0
+ lku0we = 1.8e-11
+ wk2 = -8.468563e-10
+ wlc = 0
+ wln = 1
+ ijthsrev = 0.01
+ wu0 = 4.4839114e-10
+ xgl = -8.2e-9
+ ngcon = 1
+ xgw = 0
+ epsrox = 3.9
+ wua = -5.0154626e-16
+ wub = 7.2128975e-25
+ wuc = -5.8786887e-17
+ wud = 0
+ wpclm = 1.8489068e-7
+ wwc = 0
+ kvth0we = -0.00022
+ wwl = 0
+ wwn = 1
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ gbmin = 1e-12
+ lintnoi = -5e-9
+ rdsmod = 0
+ jswgd = 3.69e-13
+ bigbinv = 0.00149
+ jswgs = 3.69e-13
+ wags = 1.2271418e-6
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ igbmod = 1
+ wcit = 1.2187445e-10
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ voff = -0.12078969
+ acde = 0.5
+ pbswgd = 0.8
+ pbswgs = 0.8
+ ppdiblc2 = -1.4649193e-16
+ vsat = 129757.01
+ wint = 0
+ vth0 = -0.42299743
+ igcmod = 1
+ wkt1 = -7.259963e-10
+ wkt2 = -1.475296e-8
+ wmax = 9.025999999999999e-7
+ aigc = 0.0068091352
+ wmin = 5.426e-7
+ wua1 = -2.7074066e-16
+ wub1 = 1.2881293e-25
+ wuc1 = 1.8593804e-16
+ tvoff = 0.0020411307
+ bigc = 0.0012521
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ wwlc = 0
+ pkvth0we = 0.0
+ nfactor = 1
+ cdsc = 0
+ cgbo = 0
+ cgdl = 2.799765e-11
+ cgdo = 2.4628259999999997e-11
+ xtid = 3
+ xtis = 3
+ permod = 1
+ ku0we = -0.0007
+ cgsl = 2.799765e-11
+ cgso = 2.4628259999999997e-11
+ cigc = 0.15259
+ beta0 = 13.32
+ vfbsdoff = 0.01
+ leta0 = -5e-10
+ ppclm = -4.9739531e-14
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ nigbacc = 10
+ paramchk = 1
+ voffcv = -0.125
+ wpemod = 1
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ nigbinv = 2.171
+ k2we = 5e-5
+ dsub = 0.5
+ ijthdfwd = 0.01
+ dtox = 3.91e-10
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ bigsd = 0.0003327
+ eta0 = 0.191845
+ tpbswg = 0.001
+ etab = -0.18516667
+ wvoff = -5.8091978e-9
+ fnoimod = 1
+ ijthdrev = 0.01
+ eigbinv = 1.1
+ wvsat = -0.017628054
+ wvth0 = -8.6541529e-9
+ lpdiblc2 = -9.0555048e-10
+ wtvfbsdoff = 0
+ ptvoff = 1.3445493e-16
+ waigc = -2.4575845e-11
+ waigsd = 1.9150694e-12
+ ltvfbsdoff = 0
+ lketa = -3.9112692e-9
+ diomod = 1
+ xpart = 1
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.9367000000000001e-10
+ pku0we = 0.0
+ cjswgs = 1.9367000000000001e-10
+ cigbacc = 0.245
+ egidl = 0.001
+ lkvth0we = 3e-12
+ tnoimod = 0
+ mjswgd = 0.95
+ mjswgs = 0.95
+ cigbinv = 0.006
+ tcjswg = 0.00128
+ pvfbsdoff = 0
+ ptvfbsdoff = 0
+ acnqsmod = 0
+ )

.model pch_ss_22 pmos (
+ level = 54
+ xrcrg1 = 12
+ xrcrg2 = 1
+ paramchk = 1
+ rshg = 14.1
+ nfactor = 1
+ wtvoff = 2.0697628e-9
+ ijthdfwd = 0.01
+ capmod = 2
+ tvoff = -0.0031746364
+ tnom = 25
+ wku0we = 1.5e-11
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ toxe = 2.71e-9
+ toxm = 2.67e-9
+ mobmod = 0
+ nigbacc = 10
+ ijthdrev = 0.01
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = -1.0551894999999999e-8
+ lpdiblc2 = 0
+ letab = 1.4778454e-8
+ nigbinv = 2.171
+ wags = -2.597049e-7
+ ppclm = 2.5985382e-14
+ wcit = 4.1443948999999997e-10
+ dlcig = 2.5e-9
+ laigsd = 2.2969081e-18
+ bgidl = 1834800000.0
+ voff = -0.11952627
+ acde = 0.5
+ vsat = 227676.61000000002
+ wint = 0
+ vth0 = -0.39483661000000003
+ a0 = 2.9368155
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ wkt1 = -1.289882e-8
+ wkt2 = 2.7006409e-8
+ at = 192293.99
+ cf = 7.598099999999999e-11
+ wmax = 9.025999999999999e-7
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.02088367
+ k3 = -2.5823
+ em = 20000000.0
+ fnoimod = 1
+ aigc = 0.0066428307
+ wmin = 5.426e-7
+ ll = 0
+ lw = 0
+ u0 = 0.008563541700000002
+ dmcgt = 0
+ w0 = 0
+ ua = -1.5734149e-9
+ ub = 3.4167628e-18
+ uc = -1.3540772e-10
+ ud = 0
+ tcjsw = 9.34e-5
+ wl = 0
+ lkvth0we = 3e-12
+ wr = 1
+ xj = 1.1e-7
+ eigbinv = 1.1
+ xl = 5.6700000000000005e-9
+ ww = 0
+ xw = 3.4e-9
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ wua1 = 6.2697239e-16
+ wub1 = -9.8389336e-25
+ wuc1 = -5.3295995e-16
+ bigc = 0.0012521
+ acnqsmod = 0
+ bigsd = 0.0003327
+ wwlc = 0
+ wvoff = -3.6240027e-9
+ cdsc = 0
+ rbodymod = 0
+ cgbo = 0
+ cgdl = 2.799765e-11
+ cgdo = 2.4628259999999997e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 2.799765e-11
+ cgso = 2.4628259999999997e-11
+ cigbacc = 0.245
+ wvsat = -0.079474309
+ cigc = 0.15259
+ wvth0 = -1.2111360000000054e-10
+ waigc = 3.8715701e-11
+ tnoimod = 0
+ toxref = 3e-9
+ lketa = 1.7736502e-8
+ cigbinv = 0.006
+ xpart = 1
+ wpdiblc2 = 6.2191766e-10
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ egidl = 0.001
+ version = 4.5
+ ltvoff = 2.5685776e-10
+ k2we = 5e-5
+ tempmod = 0
+ dsub = 0.5
+ dtox = 3.91e-10
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ pvfbsdoff = 0
+ aigbacc = 0.012071
+ eta0 = 0.29878005
+ etab = -0.34238426
+ wkvth0we = 0.0
+ lku0we = 1.8e-11
+ epsrox = 3.9
+ trnqsmod = 0
+ rdsmod = 0
+ aigbinv = 0.009974
+ pvoff = 9.9320558e-17
+ igbmod = 1
+ cdscb = 0
+ cdscd = 0
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ pvsat = 5.7635488000000005e-9
+ wk2we = 0.0
+ pvth0 = -4.450018500000001e-16
+ drout = 0.56
+ pbswgd = 0.8
+ pbswgs = 0.8
+ paigc = -2.5833927e-18
+ igcmod = 1
+ voffl = 0
+ rgatemod = 0
+ tnjtsswg = 1
+ weta0 = -7.0520749e-8
+ wetab = 2.4810139e-8
+ lpclm = -5.2812564e-8
+ poxedge = 1
+ cgidl = 1
+ binunit = 2
+ paigsd = -2.080997e-24
+ pbswd = 0.9
+ pbsws = 0.9
+ permod = 1
+ keta = -0.30513509
+ pdits = 0
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ jtsswgd = 1.75e-7
+ lcit = 2.6269861e-10
+ jtsswgs = 1.75e-7
+ voffcv = -0.125
+ wpemod = 1
+ kt1l = 0
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ lint = 0
+ lkt1 = -5.1189262e-9
+ lkt2 = 3.753071e-9
+ lmax = 8.833e-8
+ lmin = 5.233e-8
+ tnoia = 0
+ lpe0 = 6.44e-8
+ lpeb = 0
+ ijthsfwd = 0.01
+ peta0 = 4.3089229e-15
+ petab = -1.0404991e-15
+ wketa = 1.6222018e-7
+ minv = -0.33
+ wtvfbsdoff = 0
+ lua1 = 1.1693458e-16
+ lub1 = -2.0580342e-25
+ luc1 = -5.5456179e-17
+ tpbsw = 0.0025
+ tpbswg = 0.001
+ ndep = 1e+18
+ cjswd = 5.457e-11
+ njtsswg = 6.489
+ cjsws = 5.457e-11
+ mjswd = 0.01
+ lwlc = 0
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ moin = 5.5538
+ ltvfbsdoff = 0
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ ijthsrev = 0.01
+ nigc = 2.291
+ ckappad = 0.6
+ ckappas = 0.6
+ ags = 4.48665
+ pdiblc1 = 0
+ pdiblc2 = 0.0019609567
+ ptvoff = -1.0118352e-16
+ pdiblcb = 0
+ cjd = 0.00144022
+ cit = -0.0012709424099999998
+ waigsd = 1.9150916e-12
+ cjs = 0.00144022
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ noff = 2.2684
+ bvs = 8.2
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ dlc = 4.0349e-9
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ diomod = 1
+ scref = 1e-6
+ ntox = -1.9260000000000002
+ pcit = -6.38866987e-17
+ pclm = 2.1268063
+ la0 = -1.9926782e-7
+ pditsd = 0
+ pditsl = 0
+ ppdiblc2 = 0
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = -0.0067180887
+ cjswgd = 1.9367000000000001e-10
+ pku0we = 0.0
+ pigcd = 2.572
+ kt1 = -0.26717441
+ cjswgs = 1.9367000000000001e-10
+ kt2 = -0.13819145
+ lk2 = 4.8104354e-9
+ aigsd = 0.0063634181
+ bigbacc = 0.0054401
+ llc = 0
+ ptvfbsdoff = 0
+ lln = 1
+ lu0 = -1.3209508e-10
+ mjd = 0.335
+ mjs = 0.335
+ lua = 6.8530064e-17
+ lub = -1.6632734e-25
+ luc = 7.5845372e-18
+ lud = 0
+ tvfbsdoff = 0.1
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 2.4118768e-14
+ phin = 0.15
+ lvoff = -2.5437461e-9
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 2.0972465e-9
+ pbs = 0.75
+ pk2 = 2.0570947e-16
+ pu0 = 1.8416833e-16
+ kvth0we = -0.00022
+ prt = 0
+ pua = -1.7823119e-23
+ pub = 1.268951e-31
+ puc = -7.4643321e-24
+ pud = 0
+ pkt1 = 2.6862803e-15
+ pkt2 = -1.6460695e-15
+ lvsat = -0.0089644412
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = -1.4241889e-9
+ ub1 = 2.5868363e-18
+ mjswgd = 0.95
+ lvth0 = 7.3686409e-10
+ uc1 = 9.3723935e-10
+ mjswgs = 0.95
+ lintnoi = -5e-9
+ tpb = 0.0016
+ wa0 = -5.5297601e-7
+ delta = 0.018814
+ bigbinv = 0.00149
+ ute = -1
+ vtsswgd = 1.1
+ wat = -0.070679454
+ laigc = -9.8025804e-12
+ vtsswgs = 1.1
+ tcjswg = 0.00128
+ web = 6628.3
+ wec = -16935.0
+ wk2 = -1.7106076e-9
+ wlc = 0
+ wln = 1
+ wu0 = -1.5951011e-9
+ xgl = -8.2e-9
+ xgw = 0
+ wua = 2.2095182e-16
+ wub = -1.4911779e-24
+ wuc = 1.1260467e-16
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ rnoia = 0
+ rnoib = 0
+ rbdb = 50
+ pua1 = -5.0424332e-24
+ prwb = 0
+ pub1 = 1.2644812e-32
+ prwg = 0
+ puc1 = 3.7853356e-23
+ pkvth0we = 0.0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ pketa = -1.2596682e-14
+ ngate = 1.7e+20
+ rdsw = 200
+ ngcon = 1
+ wvfbsdoff = 0
+ wpclm = -6.2069351e-7
+ lvfbsdoff = 0
+ vfbsdoff = 0.01
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ fprout = 200
+ )

.model pch_ss_23 pmos (
+ level = 54
+ ijthsfwd = 0.01
+ dtox = 3.91e-10
+ cgidl = 1
+ wku0we = 1.5e-11
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ mobmod = 0
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ eta0 = 7.956713e-6
+ etab = -0.26192508
+ pbswd = 0.9
+ pbsws = 0.9
+ ijthsrev = 0.01
+ pdits = 0
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ ppdiblc2 = 0
+ njtsswg = 6.489
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ tnoia = 0
+ ckappad = 0.6
+ ckappas = 0.6
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ pdiblc1 = 0
+ pdiblc2 = 0.0019609567
+ pdiblcb = 0
+ peta0 = -2.8142439000000002e-15
+ petab = -1.6989745e-15
+ wketa = -4.2902456e-7
+ tpbsw = 0.0025
+ cjswd = 5.457e-11
+ cjsws = 5.457e-11
+ pkvth0we = 0.0
+ ags = 4.48665
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ cjd = 0.00144022
+ cit = -0.003819488
+ cjs = 0.00144022
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 4.0349e-9
+ bigbacc = 0.0054401
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ vfbsdoff = 0.01
+ a0 = 5.6551822
+ a1 = 0
+ a2 = 1
+ keta = 0.46798148
+ b0 = 0
+ b1 = 0
+ kvth0we = -0.00022
+ at = -40561.437
+ cf = 7.598099999999999e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.018874979
+ k3 = -2.5823
+ em = 20000000.0
+ la0 = -3.569331e-7
+ toxref = 3e-9
+ ll = 0
+ jsd = 1.5e-7
+ lw = 0
+ jss = 1.5e-7
+ lat = 0.0067875263
+ u0 = 0.0075684759
+ w0 = 0
+ kt1 = -0.46532049
+ kt2 = 0.0072316444
+ lk2 = 4.6939313e-9
+ ua = 5.3944309e-9
+ ub = -7.556367300000001e-18
+ uc = 1.0922891e-10
+ ud = 0
+ llc = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 5.6700000000000005e-9
+ ww = 0
+ lln = 1
+ xw = 3.4e-9
+ lu0 = -7.438127e-11
+ mjd = 0.335
+ lintnoi = -5e-9
+ mjs = 0.335
+ lua = -3.3560499e-16
+ lub = 4.7011424e-25
+ luc = -6.604387e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ bigbinv = 0.00149
+ njs = 1.02
+ pa0 = 1.517818e-13
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ nsd = 1e+20
+ lcit = 4.1051019e-10
+ pbd = 0.75
+ pat = -1.8496379e-9
+ pbs = 0.75
+ pk2 = 4.9657487e-16
+ paramchk = 1
+ pu0 = -8.1141216e-17
+ scref = 1e-6
+ kt1l = 0
+ prt = 0
+ pua = 1.7043409e-22
+ pub = -3.4495866000000004e-31
+ puc = 5.8491101e-24
+ pud = 0
+ pigcd = 2.572
+ rsh = 15.2
+ aigsd = 0.0063634182
+ tcj = 0.000832
+ ua1 = 9.464156e-9
+ tvfbsdoff = 0.1
+ ub1 = -1.352433e-17
+ uc1 = -1.5339544e-9
+ tpb = 0.0016
+ wa0 = -2.7540628e-6
+ lint = 0
+ ute = -1
+ wat = -0.002629722
+ lvoff = -5.520199e-9
+ web = 6628.3
+ wec = -16935.0
+ wk2 = -6.7255282e-9
+ wlc = 0
+ wln = 1
+ lkt1 = 6.3735466e-9
+ lkt2 = -4.6814687e-9
+ wu0 = 2.9792015e-9
+ xgl = -8.2e-9
+ xgw = 0
+ ltvoff = -2.6406105e-10
+ wua = -3.0248621e-15
+ wub = 6.6442312e-24
+ wuc = -1.1693744e-16
+ wud = 0
+ lmax = 5.233e-8
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ lmin = 4.333e-8
+ lvsat = 0.0064751142
+ lpe0 = 6.44e-8
+ lvth0 = -7.8098398e-9
+ lpeb = 0
+ ijthdfwd = 0.01
+ delta = 0.018814
+ laigc = -1.6050622e-11
+ minv = -0.33
+ lua1 = -5.1458943e-16
+ lub1 = 7.2864421e-25
+ luc1 = 8.7873061e-17
+ rnoia = 0
+ rnoib = 0
+ ndep = 1e+18
+ lku0we = 1.8e-11
+ lwlc = 0
+ epsrox = 3.9
+ moin = 5.5538
+ pketa = 2.1695512e-14
+ ngate = 1.7e+20
+ wvfbsdoff = 0
+ ijthdrev = 0.01
+ lvfbsdoff = 0
+ ngcon = 1
+ nigc = 2.291
+ wpclm = -1.0386396e-6
+ nfactor = 1
+ rdsmod = 0
+ igbmod = 1
+ lpdiblc2 = 0
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ noff = 2.2684
+ pscbe1 = 926400000.0
+ noia = 2.86e+42
+ pscbe2 = 1e-20
+ noib = 2.5e+24
+ noic = 31000000000.0
+ pbswgd = 0.8
+ pbswgs = 0.8
+ igcmod = 1
+ ntox = -1.9260000000000002
+ pcit = -2.400000000060939e-23
+ pclm = 4.4879115
+ nigbacc = 10
+ phin = 0.15
+ lkvth0we = 3e-12
+ pkt1 = -5.0612736e-15
+ pkt2 = 1.1767646e-15
+ nigbinv = 2.171
+ tvoff = 0.0058067224
+ acnqsmod = 0
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ rbdb = 50
+ pua1 = 2.7224008e-22
+ prwb = 0
+ pub1 = -3.6990718e-31
+ prwg = 0
+ puc1 = -5.7927018e-23
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ permod = 1
+ rbodymod = 0
+ rdsw = 200
+ ku0we = -0.0007
+ beta0 = 13.32
+ fnoimod = 1
+ leta0 = 6.7768865999999995e-9
+ letab = 1.0111821e-8
+ eigbinv = 1.1
+ ppclm = 5.0226256e-14
+ voffcv = -0.125
+ wpemod = 1
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ rshg = 14.1
+ wtvfbsdoff = 0
+ wpdiblc2 = 6.2191766e-10
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ ltvfbsdoff = 0
+ cigbacc = 0.245
+ tnoimod = 0
+ tnom = 25
+ tpbswg = 0.001
+ bigsd = 0.0003327
+ toxe = 2.71e-9
+ toxm = 2.67e-9
+ cigbinv = 0.006
+ wkvth0we = 0.0
+ wvoff = -2.1208799e-8
+ trnqsmod = 0
+ wvsat = 0.11762556
+ ptvoff = 1.2747838e-16
+ ptvfbsdoff = 0
+ wvth0 = -2.9965608e-8
+ waigsd = 1.9150557e-12
+ version = 4.5
+ waigc = -1.4751759e-11
+ wags = -2.597049e-7
+ tempmod = 0
+ wcit = -6.870588899999999e-10
+ diomod = 1
+ voff = -0.068208113
+ lketa = -2.7104259e-8
+ acde = 0.5
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.9367000000000001e-10
+ pku0we = 0.0
+ cjswgs = 1.9367000000000001e-10
+ aigbacc = 0.012071
+ xpart = 1
+ rgatemod = 0
+ vsat = -38522.667
+ wint = 0
+ vth0 = -0.24747999999999998
+ tnjtsswg = 1
+ wkt1 = 1.206797e-7
+ wkt2 = -2.1663145e-8
+ egidl = 0.001
+ wmax = 9.025999999999999e-7
+ aigc = 0.0067505556
+ wmin = 5.426e-7
+ mjswgd = 0.95
+ mjswgs = 0.95
+ aigbinv = 0.009974
+ tcjswg = 0.00128
+ pvfbsdoff = 0
+ wua1 = -4.1537606e-15
+ wub1 = 5.6118307e-24
+ wuc1 = 1.1184258e-15
+ bigc = 0.0012521
+ wwlc = 0
+ cdsc = 0
+ cgbo = 0
+ cgdl = 2.799765e-11
+ cgdo = 2.4628259999999997e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 2.799765e-11
+ cgso = 2.4628259999999997e-11
+ cigc = 0.15259
+ pvoff = 1.1192388e-15
+ poxedge = 1
+ cdscb = 0
+ cdscd = 0
+ fprout = 200
+ pvsat = -5.6682454999999995e-9
+ wk2we = 0.0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ pvth0 = 1.2859777e-15
+ drout = 0.56
+ binunit = 2
+ paigc = 5.1772001e-19
+ voffl = 0
+ dmcg = 3.1e-8
+ wtvoff = -1.8726837e-9
+ dmci = 3.1e-8
+ dmdg = 0
+ weta0 = 5.2292471e-8
+ wetab = 3.6163164e-8
+ lpclm = -1.8975667e-7
+ k2we = 5e-5
+ capmod = 2
+ dsub = 0.5
+ )

.model pch_ss_24 pmos (
+ level = 54
+ beta0 = 13.32
+ leta0 = -4.419176000000001e-11
+ letab = 2.8639817e-9
+ cigbacc = 0.245
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ ppclm = -6.983762e-15
+ laigsd = -1.7489044e-14
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ tnoimod = 0
+ ntox = -1.9260000000000002
+ pcit = -5.985074999999999e-17
+ pclm = 0.55996802
+ rgatemod = 0
+ cigbinv = 0.006
+ tnjtsswg = 1
+ phin = 0.15
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ pkt1 = 8.0439909e-15
+ pkt2 = -6.3201272e-16
+ version = 4.5
+ tempmod = 0
+ bigsd = 0.0003327
+ rbdb = 50
+ pua1 = -2.7866327e-22
+ prwb = 0
+ pub1 = 3.3701988e-31
+ prwg = 0
+ puc1 = 2.5974765e-23
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ aigbacc = 0.012071
+ wvoff = -2.6959456e-8
+ rdsw = 200
+ wvsat = 0.025612403
+ wvth0 = 5.670831900000001e-9
+ toxref = 3e-9
+ waigc = -9.7737582e-11
+ aigbinv = 0.009974
+ lketa = 1.4220453e-8
+ rshg = 14.1
+ xpart = 1
+ egidl = 0.001
+ ltvoff = -2.5344658e-10
+ pvfbsdoff = 0
+ ijthsfwd = 0.01
+ poxedge = 1
+ a0 = -2.5402778
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ tnom = 25
+ at = 223221.03
+ cf = 7.598099999999999e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.022656115
+ k3 = -2.5823
+ em = 20000000.0
+ lku0we = 1.8e-11
+ ll = 0
+ lw = 0
+ u0 = 0.0016778574000000002
+ w0 = 0
+ toxe = 2.71e-9
+ toxm = 2.67e-9
+ ua = -6.0379704e-9
+ ub = 7.7295729e-18
+ uc = -2.2784413e-10
+ ud = 0
+ binunit = 2
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 5.6700000000000005e-9
+ ww = 0
+ epsrox = 3.9
+ xw = 3.4e-9
+ ijthsrev = 0.01
+ rdsmod = 0
+ igbmod = 1
+ pvoff = 1.401021e-15
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ wags = -2.597049e-7
+ cdscb = 0
+ cdscd = 0
+ pbswgd = 0.8
+ pbswgs = 0.8
+ pvsat = -1.1596007e-9
+ wcit = 5.343688999999993e-10
+ wk2we = 0.0
+ pvth0 = -4.6020083e-16
+ drout = 0.56
+ igcmod = 1
+ voff = -0.080254273
+ paigc = 4.5840253e-18
+ acde = 0.5
+ ppdiblc2 = 0
+ voffl = 0
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ vsat = 108578.56
+ wint = 0
+ vth0 = -0.37982436
+ wkt1 = -1.4677468e-7
+ wkt2 = 1.5250678e-8
+ wmax = 9.025999999999999e-7
+ weta0 = -2.1433527999999997e-8
+ aigc = 0.0066531108
+ wetab = 8.325777e-9
+ wmin = 5.426e-7
+ lpclm = 2.7125638e-9
+ cgidl = 1
+ paigsd = 9.5490179e-21
+ wua1 = 7.089165e-15
+ wub1 = -8.8152527e-24
+ wuc1 = -5.9385548e-16
+ bigc = 0.0012521
+ wwlc = 0
+ pkvth0we = 0.0
+ permod = 1
+ cdsc = 0
+ pbswd = 0.9
+ pbsws = 0.9
+ njtsswg = 6.489
+ cgbo = 0
+ cgdl = 2.799765e-11
+ cgdo = 2.4628259999999997e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 2.799765e-11
+ cgso = 2.4628259999999997e-11
+ wtvfbsdoff = 0
+ cigc = 0.15259
+ vfbsdoff = 0.01
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ ckappad = 0.6
+ ckappas = 0.6
+ pdits = 0
+ voffcv = -0.125
+ wpemod = 1
+ pdiblc1 = 0
+ pdiblc2 = 0.0019609567
+ cigsd = 0.013281
+ ltvfbsdoff = 0
+ pdiblcb = 0
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ paramchk = 1
+ pk2we = 0.0
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ bigbacc = 0.0054401
+ tnoia = 0
+ k2we = 5e-5
+ ags = 4.48665
+ ijthdfwd = 0.01
+ dsub = 0.5
+ dtox = 3.91e-10
+ kvth0we = -0.00022
+ peta0 = 7.9833004e-16
+ ptvfbsdoff = 0
+ petab = -3.349425e-16
+ cjd = 0.00144022
+ cit = 0.0027658070000000003
+ cjs = 0.00144022
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dvt0 = 3.48
+ tpbswg = 0.001
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ wketa = 1.6324308e-7
+ dlc = 4.0349e-9
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ tpbsw = 0.0025
+ dwg = 0
+ lintnoi = -5e-9
+ dwj = 0
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ cjswd = 5.457e-11
+ cjsws = 5.457e-11
+ mjswd = 0.01
+ eta0 = 0.13921364
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ etab = -0.11400999
+ la0 = 4.4644444e-8
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = -0.0061378147
+ kt1 = 0.16833478
+ kt2 = -0.11193164
+ lk2 = 4.879207e-9
+ ijthdrev = 0.01
+ llc = 0
+ lln = 1
+ lu0 = 2.1425904e-10
+ mjd = 0.335
+ ptvoff = 8.5019581e-17
+ mjs = 0.335
+ lua = 2.2458267e-16
+ lub = -2.7889682000000003e-25
+ luc = 9.9121919e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = -8.9774533e-14
+ waigsd = 1.7201778e-12
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 7.328227899999999e-9
+ pbs = 0.75
+ lpdiblc2 = 0
+ pk2 = 1.0702031e-16
+ pu0 = -9.6657248e-17
+ prt = 0
+ pua = -9.0705467e-23
+ pub = 1.1140901e-31
+ puc = -1.0416838e-23
+ pud = 0
+ diomod = 1
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = -1.018181e-8
+ ub1 = 1.2730062e-17
+ uc1 = 9.111363e-10
+ tpb = 0.0016
+ wa0 = 2.1756583e-6
+ ute = -1
+ wat = -0.18993311000000002
+ pditsd = 0
+ web = 6628.3
+ wec = -16935.0
+ pditsl = 0
+ wk2 = 1.2245648e-9
+ cjswgd = 1.9367000000000001e-10
+ pku0we = 0.0
+ cjswgs = 1.9367000000000001e-10
+ wlc = 0
+ wln = 1
+ wu0 = 3.2958552e-9
+ xgl = -8.2e-9
+ xgw = 0
+ scref = 1e-6
+ wua = 2.3045166e-15
+ wub = -2.6693944999999998e-24
+ wuc = 2.150207e-16
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ tvfbsdoff = 0.1
+ pigcd = 2.572
+ aigsd = 0.0063637751
+ lvoff = -4.9299372e-9
+ mjswgd = 0.95
+ mjswgs = 0.95
+ lkvth0we = 3e-12
+ nfactor = 1
+ lvsat = -0.00073284372
+ tcjswg = 0.00128
+ lvth0 = -1.3249514899999999e-9
+ delta = 0.018814
+ laigc = -1.1275829e-11
+ acnqsmod = 0
+ rnoia = 0
+ rnoib = 0
+ wvfbsdoff = 0
+ pketa = -7.3256019e-15
+ ngate = 1.7e+20
+ lvfbsdoff = 0
+ rbodymod = 0
+ nigbacc = 10
+ ngcon = 1
+ wpclm = 1.2891178e-7
+ gbmin = 1e-12
+ keta = -0.37538
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ fprout = 200
+ xrcrg1 = 12
+ xrcrg2 = 1
+ nigbinv = 2.171
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 8.783704000000003e-11
+ kt1l = 0
+ wtvoff = -1.0061777e-9
+ wpdiblc2 = 6.2191766e-10
+ lint = 0
+ lkt1 = -2.4675560999999998e-8
+ lkt2 = 1.1575324e-9
+ lmax = 4.333e-8
+ lmin = 3.6e-8
+ capmod = 2
+ fnoimod = 1
+ lpe0 = 6.44e-8
+ lpeb = 0
+ wku0we = 1.5e-11
+ eigbinv = 1.1
+ tvoff = 0.0055901005
+ mobmod = 0
+ minv = -0.33
+ lua1 = 4.4806289e-16
+ lub1 = -5.5782098e-25
+ luc1 = -3.1936385e-17
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ ndep = 1e+18
+ wkvth0we = 0.0
+ lwlc = 0
+ moin = 5.5538
+ nigc = 2.291
+ trnqsmod = 0
+ ku0we = -0.0007
+ )

.model pch_ss_25 pmos (
+ level = 54
+ wint = 0
+ ags = 0.93810347
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ vth0 = -0.40498248000000003
+ wkt1 = -1.5318394e-9
+ wkt2 = 2.21858e-9
+ cjd = 0.00144022
+ cit = 5e-6
+ cjs = 0.00144022
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ wmax = 5.426e-7
+ bvs = 8.2
+ aigc = 0.0068215676
+ wmin = 2.726e-7
+ dlc = 1.0572421799999999e-8
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ k3b = 2.1176
+ lkvth0we = 3e-12
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ tnoia = 0
+ peta0 = -1.5e-17
+ la0 = 0
+ wua1 = 1.6452204e-16
+ wub1 = -6.9710259e-26
+ wuc1 = 2.1709154e-17
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0.001
+ wketa = 2.2687563e-8
+ kt1 = -0.17747938
+ lk2 = 4e-10
+ kt2 = -0.061438333
+ llc = 0
+ lln = 1
+ lu0 = 5e-12
+ tpbsw = 0.0025
+ acnqsmod = 0
+ mjd = 0.335
+ bigc = 0.0012521
+ mjs = 0.335
+ wute = 3.2371733e-8
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ wwlc = 0
+ pa0 = 0
+ cjswd = 5.457e-11
+ nsd = 1e+20
+ cjsws = 5.457e-11
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ pk2 = 0
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ pu0 = 0
+ prt = 0
+ pud = 0
+ rbodymod = 0
+ cdsc = 0
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 1.8507467e-10
+ ub1 = -1.7337534e-19
+ uc1 = -4.0886356e-11
+ cgbo = 0
+ cgdl = 2.799765e-11
+ cgdo = 2.4628259999999997e-11
+ xtid = 3
+ xtis = 3
+ tpb = 0.0016
+ wa0 = -1.5013787e-7
+ cgsl = 2.799765e-11
+ cgso = 2.4628259999999997e-11
+ cigc = 0.15259
+ ute = -1.2102889
+ toxref = 3e-9
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 4.440518e-10
+ wlc = 0
+ wln = 1
+ wu0 = 3.7953067e-11
+ xgl = -8.2e-9
+ xgw = 0
+ nfactor = 1
+ wua = -1.5196107e-16
+ wub = 9.0507286e-26
+ wuc = 5.3799588e-18
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ scref = 1e-6
+ tvfbsdoff = 0.1
+ pigcd = 2.572
+ aigsd = 0.0063632886
+ wpdiblc2 = -7.7579138e-11
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ ltvoff = 0
+ lvoff = 0
+ nigbacc = 10
+ lvsat = 0.00024
+ k2we = 5e-5
+ lvth0 = -6e-10
+ dsub = 0.5
+ dtox = 3.91e-10
+ delta = 0.018814
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ lku0we = 1.8e-11
+ rnoia = 0
+ rnoib = 0
+ epsrox = 3.9
+ nigbinv = 2.171
+ eta0 = 0.17962267
+ wvfbsdoff = 0
+ wkvth0we = 0.0
+ etab = -0.19577778
+ lvfbsdoff = 0
+ ngate = 1.7e+20
+ rdsmod = 0
+ ngcon = 1
+ igbmod = 1
+ wpclm = -1.1447315e-8
+ trnqsmod = 0
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ pbswgd = 0.8
+ pbswgs = 0.8
+ fnoimod = 1
+ eigbinv = 1.1
+ igcmod = 1
+ a0 = 3.3089778
+ a1 = 0
+ a2 = 1
+ rgatemod = 0
+ b0 = 0
+ b1 = 0
+ at = 72000
+ cf = 7.598099999999999e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.0028441163
+ k3 = -2.5823
+ em = 20000000.0
+ tnjtsswg = 1
+ ll = 0
+ lw = 0
+ u0 = 0.0099214889
+ w0 = 0
+ ua = 1.8228697e-10
+ ub = 9.7616315e-19
+ uc = -9.1826044e-12
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 5.6700000000000005e-9
+ ww = 0
+ xw = 3.4e-9
+ wtvfbsdoff = 0
+ cigbacc = 0.245
+ tvoff = 0.0026578776
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ permod = 1
+ ltvfbsdoff = 0
+ tnoimod = 0
+ cigbinv = 0.006
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = -5e-10
+ keta = -0.064397096
+ voffcv = -0.125
+ wpemod = 1
+ ppclm = 0
+ version = 4.5
+ dlcig = 2.5e-9
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ bgidl = 1834800000.0
+ lcit = 0
+ tempmod = 0
+ ptvfbsdoff = 0
+ kt1l = 0
+ aigbacc = 0.012071
+ lint = 6.5375218e-9
+ dmcgt = 0
+ lkt1 = -1e-9
+ tcjsw = 9.34e-5
+ lmax = 2.001e-5
+ lmin = 8.99743e-6
+ lpe0 = 6.44e-8
+ lpeb = 0
+ ijthsfwd = 0.01
+ tpbswg = 0.001
+ minv = -0.33
+ aigbinv = 0.009974
+ bigsd = 0.0003327
+ ndep = 1e+18
+ lwlc = 0
+ moin = 5.5538
+ wvoff = 2.5521431e-9
+ ptvoff = 0
+ ijthsrev = 0.01
+ nigc = 2.291
+ waigsd = 1.9763167e-12
+ wvsat = 0.0034765009
+ wvth0 = -4.6147147e-9
+ diomod = 1
+ waigc = 4.045116e-12
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.9367000000000001e-10
+ pku0we = 0.0
+ cjswgs = 1.9367000000000001e-10
+ poxedge = 1
+ lketa = 0
+ ntox = -1.9260000000000002
+ xpart = 1
+ pcit = 0
+ pclm = 1.1689658
+ ppdiblc2 = 0
+ binunit = 2
+ egidl = 0.001
+ mjswgd = 0.95
+ mjswgs = 0.95
+ phin = 0.15
+ tcjswg = 0.00128
+ pkt1 = 0
+ pvfbsdoff = 0
+ rbdb = 50
+ prwb = 0
+ prwg = 0
+ pkvth0we = 0.0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ jtsswgd = 1.75e-7
+ rdsw = 200
+ jtsswgs = 1.75e-7
+ vfbsdoff = 0.01
+ fprout = 200
+ pvoff = 2.5e-17
+ xrcrg1 = 12
+ xrcrg2 = 1
+ cdscb = 0
+ cdscd = 0
+ pvsat = -5e-11
+ wk2we = 0.0
+ pvth0 = -7e-17
+ drout = 0.56
+ paramchk = 1
+ wtvoff = -1.0551434e-10
+ rshg = 14.1
+ voffl = 0
+ weta0 = -1.7848176e-8
+ wetab = 1.9534667e-8
+ njtsswg = 6.489
+ capmod = 2
+ lpclm = 0
+ wku0we = 1.5e-11
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ ijthdfwd = 0.01
+ cgidl = 1
+ mobmod = 0
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.0030491463
+ tnom = 25
+ pdiblcb = 0
+ toxe = 2.71e-9
+ toxm = 2.67e-9
+ pbswd = 0.9
+ pbsws = 0.9
+ ijthdrev = 0.01
+ lpdiblc2 = 0
+ bigbacc = 0.0054401
+ wags = -6.1953916e-9
+ pdits = 0
+ cigsd = 0.013281
+ kvth0we = -0.00022
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ voff = -0.10784306
+ acde = 0.5
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ vsat = 91103.982
+ pk2we = 0.0
+ )

.model pch_ss_26 pmos (
+ level = 54
+ bigsd = 0.0003327
+ poxedge = 1
+ pkvth0we = 0.0
+ wvoff = 2.9007224e-9
+ binunit = 2
+ toxref = 3e-9
+ wvsat = 0.0034765009
+ wvth0 = -4.6762891999999995e-9
+ vfbsdoff = 0.01
+ keta = -0.06875265
+ waigc = 4.3476029e-12
+ lags = 1.0877241e-7
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 0
+ lketa = 3.9156432e-8
+ paramchk = 1
+ kt1l = 0
+ xpart = 1
+ ltvoff = -4.4286369e-10
+ egidl = 0.001
+ lint = 6.5375218e-9
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ lkt1 = -3.5853729e-8
+ lkt2 = -1.4641311e-8
+ lmax = 8.99743e-6
+ pvfbsdoff = 0
+ lmin = 8.974099999999999e-7
+ lpe0 = 6.44e-8
+ ijthdfwd = 0.01
+ lpeb = 0
+ lku0we = 1.8e-11
+ minv = -0.33
+ epsrox = 3.9
+ lua1 = 1.4818924e-15
+ lub1 = -2.0711788e-24
+ luc1 = 2.2491171e-16
+ ndep = 1e+18
+ lute = 1.330224e-7
+ rdsmod = 0
+ lwlc = 0
+ moin = 5.5538
+ igbmod = 1
+ ijthdrev = 0.01
+ nigc = 2.291
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ lpdiblc2 = 8.2033961e-9
+ njtsswg = 6.489
+ pbswgd = 0.8
+ pvoff = -3.1087282000000003e-15
+ pbswgs = 0.8
+ noff = 2.2684
+ cdscb = 0
+ cdscd = 0
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ igcmod = 1
+ pvsat = -5e-11
+ wk2we = 0.0
+ pvth0 = 4.835547400000001e-16
+ drout = 0.56
+ ckappad = 0.6
+ ckappas = 0.6
+ pags = 8.2314292e-14
+ wtvfbsdoff = 0
+ pdiblc1 = 0
+ pdiblc2 = 0.002136644
+ paigc = -2.7193569e-18
+ pdiblcb = 0
+ ntox = -1.9260000000000002
+ pcit = 0
+ pclm = 1.1689658
+ voffl = 0
+ ltvfbsdoff = 0
+ weta0 = -1.7848176e-8
+ phin = 0.15
+ wetab = 1.9534667e-8
+ lkvth0we = 3e-12
+ lpclm = 0
+ paigsd = -4.5957918e-20
+ pkt1 = 4.5592526e-15
+ pkt2 = 3.8774237e-15
+ bigbacc = 0.0054401
+ cgidl = 1
+ permod = 1
+ acnqsmod = 0
+ kvth0we = -0.00022
+ rbdb = 50
+ pua1 = -9.4343892e-23
+ prwb = 0
+ pub1 = 9.0084871e-32
+ prwg = 0
+ puc1 = -7.238167e-23
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ lintnoi = -5e-9
+ pute = -1.6539558e-14
+ bigbinv = 0.00149
+ rbodymod = 0
+ pbswd = 0.9
+ pbsws = 0.9
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ rdsw = 200
+ ptvfbsdoff = 0
+ a0 = 3.4253346
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 72000
+ cf = 7.598099999999999e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.0024652651
+ k3 = -2.5823
+ em = 20000000.0
+ ll = 0
+ voffcv = -0.125
+ lw = 0
+ wpemod = 1
+ u0 = 0.0098054275
+ w0 = 0
+ ua = 1.8429003e-10
+ ub = 9.3982253e-19
+ uc = -1.1498405e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 5.6700000000000005e-9
+ ww = 0
+ xw = 3.4e-9
+ pdits = 0
+ cigsd = 0.013281
+ ags = 0.9260042
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ cjd = 0.00144022
+ cit = 5e-6
+ cjs = 0.00144022
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 1.0572421799999999e-8
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ rshg = 14.1
+ wpdiblc2 = 3.818702e-12
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ la0 = -1.0460478e-6
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0.001
+ kt1 = -0.17360244
+ kt2 = -0.059809712
+ lk2 = -3.0058721000000003e-9
+ llc = 0
+ lln = 1
+ lu0 = 1.0483917e-9
+ mjd = 0.335
+ mjs = 0.335
+ lua = -1.8007487e-17
+ lub = 3.2670219e-25
+ luc = 2.0819042e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ tnoia = 0
+ njd = 1.02
+ njs = 1.02
+ pa0 = 1.483047e-13
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ tpbswg = 0.001
+ pk2 = 2.5596912e-15
+ pu0 = 1.7642195e-17
+ nfactor = 1
+ peta0 = -1.5e-17
+ prt = 0
+ pua = 1.2819791e-23
+ pub = -1.2787603e-32
+ puc = -1.6865938e-24
+ pud = 0
+ wketa = 2.5468383e-8
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 2.0236805e-11
+ ub1 = 5.7011626e-20
+ uc1 = -6.5904343e-11
+ tnom = 25
+ tpbsw = 0.0025
+ tpb = 0.0016
+ wa0 = -1.666345e-7
+ toxe = 2.71e-9
+ toxm = 2.67e-9
+ ute = -1.2250856
+ cjswd = 5.457e-11
+ cjsws = 5.457e-11
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 1.5932531e-10
+ mjswd = 0.01
+ wlc = 0
+ mjsws = 0.01
+ wln = 1
+ agidl = 3.2166e-9
+ wu0 = 3.5990642e-11
+ wkvth0we = 0.0
+ xgl = -8.2e-9
+ xgw = 0
+ wua = -1.5338707e-16
+ wub = 9.1929712e-26
+ wuc = 5.5675666e-18
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ ptvoff = -2.4168192e-17
+ waigsd = 1.9814288e-12
+ trnqsmod = 0
+ nigbacc = 10
+ diomod = 1
+ wags = -1.5351598e-8
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.9367000000000001e-10
+ pku0we = 0.0
+ cjswgs = 1.9367000000000001e-10
+ tvfbsdoff = 0.1
+ voff = -0.10676035
+ scref = 1e-6
+ acde = 0.5
+ nigbinv = 2.171
+ pigcd = 2.572
+ rgatemod = 0
+ aigsd = 0.0063632773
+ vsat = 91103.982
+ wint = 0
+ vth0 = -0.40356355000000005
+ tnjtsswg = 1
+ mjswgd = 0.95
+ mjswgs = 0.95
+ wkt1 = -2.0389865e-9
+ wkt2 = 1.7872759e-9
+ lvoff = -9.7335308e-9
+ wmax = 5.426e-7
+ aigc = 0.0068257672
+ wmin = 2.726e-7
+ tcjswg = 0.00128
+ lvsat = 0.00024
+ lvth0 = -1.3356137e-8
+ delta = 0.018814
+ laigc = -3.7754415e-11
+ wua1 = 1.7501635e-16
+ wub1 = -7.9730823e-26
+ wuc1 = 2.9760508e-17
+ fnoimod = 1
+ rnoia = 0
+ rnoib = 0
+ bigc = 0.0012521
+ eigbinv = 1.1
+ wute = 3.4211506e-8
+ wwlc = 0
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ pketa = -2.4999571e-14
+ ngate = 1.7e+20
+ cdsc = 0
+ ngcon = 1
+ cgbo = 0
+ wpclm = -1.1447315e-8
+ cgdl = 2.799765e-11
+ cgdo = 2.4628259999999997e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 2.799765e-11
+ cgso = 2.4628259999999997e-11
+ fprout = 200
+ cigc = 0.15259
+ gbmin = 1e-12
+ xrcrg1 = 12
+ xrcrg2 = 1
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ cigbacc = 0.245
+ wtvoff = -1.02826e-10
+ tnoimod = 0
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ capmod = 2
+ cigbinv = 0.006
+ wku0we = 1.5e-11
+ k2we = 5e-5
+ mobmod = 0
+ ijthsfwd = 0.01
+ dsub = 0.5
+ dtox = 3.91e-10
+ tvoff = 0.0027071394
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ xjbvd = 1
+ xjbvs = 1
+ version = 4.5
+ lk2we = 0.0
+ tempmod = 0
+ eta0 = 0.17962267
+ etab = -0.19577778
+ ijthsrev = 0.01
+ ku0we = -0.0007
+ aigbacc = 0.012071
+ beta0 = 13.32
+ leta0 = -5e-10
+ laigsd = 1.0132005e-13
+ ppclm = 0
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ aigbinv = 0.009974
+ ppdiblc2 = -7.3176658e-16
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ )

.model pch_ss_27 pmos (
+ level = 54
+ tvfbsdoff = 0.1
+ fnoimod = 1
+ scref = 1e-6
+ eigbinv = 1.1
+ rshg = 14.1
+ ltvoff = -3.7535707e-10
+ pigcd = 2.572
+ aigsd = 0.0063633912
+ lvoff = -1.1639377e-8
+ lvsat = 0.00024
+ lvth0 = 4.506701000000001e-10
+ ijthsfwd = 0.01
+ lku0we = 1.8e-11
+ delta = 0.018814
+ laigc = -5.5983746e-11
+ epsrox = 3.9
+ tnom = 25
+ rnoia = 0
+ rnoib = 0
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ cigbacc = 0.245
+ toxe = 2.71e-9
+ toxm = 2.67e-9
+ rdsmod = 0
+ igbmod = 1
+ pketa = 5.6398736e-15
+ ngate = 1.7e+20
+ wtvfbsdoff = 0
+ ijthsrev = 0.01
+ ngcon = 1
+ tnoimod = 0
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ wpclm = -1.1447315e-8
+ pbswgd = 0.8
+ pbswgs = 0.8
+ gbmin = 1e-12
+ cigbinv = 0.006
+ jswgd = 3.69e-13
+ ltvfbsdoff = 0
+ jswgs = 3.69e-13
+ igcmod = 1
+ wags = 3.4820603e-7
+ voff = -0.10461895
+ acde = 0.5
+ version = 4.5
+ ppdiblc2 = 9.4893758e-16
+ vsat = 91103.982
+ tempmod = 0
+ wint = 0
+ vth0 = -0.41907682
+ wkt1 = 1.4552168e-8
+ wkt2 = 6.9668931e-9
+ wmax = 5.426e-7
+ aigc = 0.0068462496
+ wmin = 2.726e-7
+ aigbacc = 0.012071
+ ptvfbsdoff = 0
+ tvoff = 0.0026312893
+ wua1 = 1.777316e-16
+ wub1 = 1.5048515e-26
+ wuc1 = -3.1929257e-17
+ permod = 1
+ xjbvd = 1
+ xjbvs = 1
+ bigc = 0.0012521
+ wute = 6.965504e-8
+ lk2we = 0.0
+ wwlc = 0
+ pkvth0we = 0.0
+ aigbinv = 0.009974
+ cdsc = 0
+ cgbo = 0
+ cgdl = 2.799765e-11
+ cgdo = 2.4628259999999997e-11
+ xtid = 3
+ xtis = 3
+ ku0we = -0.0007
+ beta0 = 13.32
+ cgsl = 2.799765e-11
+ cgso = 2.4628259999999997e-11
+ voffcv = -0.125
+ wpemod = 1
+ cigc = 0.15259
+ vfbsdoff = 0.01
+ leta0 = -5e-10
+ ppclm = 0
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ paramchk = 1
+ poxedge = 1
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ binunit = 2
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ tpbswg = 0.001
+ k2we = 5e-5
+ ijthdfwd = 0.01
+ dsub = 0.5
+ dtox = 3.91e-10
+ a0 = 2.4559917
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 72000
+ cf = 7.598099999999999e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.0065510297
+ k3 = -2.5823
+ em = 20000000.0
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ ll = 0
+ lw = 0
+ u0 = 0.011339968
+ w0 = 0
+ ua = 2.2475737e-10
+ ub = 1.3971204e-18
+ uc = 8.9671176e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 5.6700000000000005e-9
+ ww = 0
+ xw = 3.4e-9
+ bigsd = 0.0003327
+ ptvoff = 6.0034078e-17
+ eta0 = 0.17962267
+ etab = -0.19577778
+ waigsd = 1.9297907e-12
+ wvoff = -2.3606869e-9
+ ijthdrev = 0.01
+ wvsat = 0.0034765009
+ diomod = 1
+ wvth0 = -3.9167848e-9
+ lpdiblc2 = -1.0873556e-9
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ waigc = -6.0221967e-12
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.9367000000000001e-10
+ pku0we = 0.0
+ cjswgs = 1.9367000000000001e-10
+ lketa = -2.7133526e-8
+ xpart = 1
+ mjswgd = 0.95
+ mjswgs = 0.95
+ egidl = 0.001
+ tcjswg = 0.00128
+ pvfbsdoff = 0
+ lkvth0we = 3e-12
+ njtsswg = 6.489
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ acnqsmod = 0
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.012575691
+ pdiblcb = 0
+ rbodymod = 0
+ fprout = 200
+ xrcrg1 = 12
+ xrcrg2 = 1
+ pvoff = 1.5739261e-15
+ keta = 0.0057304489
+ cdscb = 0
+ cdscd = 0
+ pvsat = -5e-11
+ bigbacc = 0.0054401
+ lags = 9.833094e-7
+ wk2we = 0.0
+ pvth0 = -1.9240418e-16
+ wtvoff = -1.9743529e-10
+ drout = 0.56
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 8.2671111e-11
+ paigc = 6.5097646e-18
+ kt1l = 0
+ kvth0we = -0.00022
+ voffl = 0
+ wpdiblc2 = -1.8846129e-9
+ lintnoi = -5e-9
+ capmod = 2
+ lint = 6.5375218e-9
+ bigbinv = 0.00149
+ weta0 = -1.7848176e-8
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ wetab = 1.9534667e-8
+ wku0we = 1.5e-11
+ lkt1 = -5.3329349e-9
+ lkt2 = -2.567581e-9
+ lpclm = 0
+ lmax = 8.974099999999999e-7
+ lmin = 4.4741e-7
+ mobmod = 0
+ lpe0 = 6.44e-8
+ lpeb = 0
+ cgidl = 1
+ minv = -0.33
+ lua1 = 1.3348283e-16
+ lub1 = 2.1611253e-25
+ luc1 = 5.928335e-17
+ ndep = 1e+18
+ lute = 1.2896693e-7
+ wkvth0we = 0.0
+ lwlc = 0
+ moin = 5.5538
+ pbswd = 0.9
+ pbsws = 0.9
+ ags = -0.056621626
+ nigc = 2.291
+ trnqsmod = 0
+ cjd = 0.00144022
+ cit = -8.7888889e-5
+ cjs = 0.00144022
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 1.0572421799999999e-8
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ pdits = 0
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ cigsd = 0.013281
+ nfactor = 1
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ la0 = -1.8333262e-7
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0.001
+ pags = -2.41252e-13
+ kt1 = -0.20789546
+ kt2 = -0.0733757
+ lk2 = 6.3045842e-10
+ llc = 0
+ lln = 1
+ lu0 = -3.1734965000000004e-10
+ mjd = 0.335
+ mjs = 0.335
+ lua = -5.402342e-17
+ lub = -8.029291e-26
+ luc = -6.9221885e-17
+ lud = 0
+ ntox = -1.9260000000000002
+ lwc = 0
+ lwl = 0
+ pcit = 0
+ lwn = 1
+ pclm = 1.1689658
+ njd = 1.02
+ njs = 1.02
+ pa0 = -1.295362e-13
+ rgatemod = 0
+ nsd = 1e+20
+ pbd = 0.75
+ pk2we = 0.0
+ pat = 0
+ pbs = 0.75
+ pk2 = 6.34174e-16
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ tnjtsswg = 1
+ pu0 = -2.5304972e-16
+ prt = 0
+ pua = -1.1377853e-22
+ pub = 1.1787175e-31
+ puc = 2.8393052e-23
+ pud = 0
+ phin = 0.15
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 1.5353037e-9
+ ub1 = -2.5129786e-18
+ uc1 = 1.2019494e-10
+ tpb = 0.0016
+ tnoia = 0
+ wa0 = 1.4554629e-7
+ pkt1 = -1.0206874e-14
+ pkt2 = -7.3243565e-16
+ ute = -1.2205289
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 2.3228278e-9
+ nigbacc = 10
+ wlc = 0
+ wln = 1
+ wu0 = 3.4013886e-10
+ xgl = -8.2e-9
+ xgw = 0
+ peta0 = -1.5e-17
+ wua = -1.1141771e-17
+ wub = -5.4878553e-26
+ wuc = -2.8229789e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ wketa = -8.9579586e-9
+ tpbsw = 0.0025
+ cjswd = 5.457e-11
+ cjsws = 5.457e-11
+ rbdb = 50
+ pua1 = -9.6760461e-23
+ prwb = 0
+ pub1 = 5.7312604e-33
+ prwg = 0
+ puc1 = -1.747778e-23
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ nigbinv = 2.171
+ pute = -4.8084303e-14
+ rdsw = 200
+ toxref = 3e-9
+ )

.model pch_ss_28 pmos (
+ level = 54
+ wtvfbsdoff = 0
+ lku0we = 1.8e-11
+ k2we = 5e-5
+ epsrox = 3.9
+ dsub = 0.5
+ dtox = 3.91e-10
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ ltvfbsdoff = 0
+ bigbacc = 0.0054401
+ rdsmod = 0
+ igbmod = 1
+ wkvth0we = 0.0
+ eta0 = 0.17962267
+ etab = -0.19577778
+ kvth0we = -0.00022
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ trnqsmod = 0
+ pbswgd = 0.8
+ lintnoi = -5e-9
+ pbswgs = 0.8
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ pvoff = -2.0154208999999999e-16
+ igcmod = 1
+ cdscb = 0
+ cdscd = 0
+ pvsat = -5e-11
+ wk2we = 0.0
+ pvth0 = -7.6676914e-16
+ ptvfbsdoff = 0
+ drout = 0.56
+ paigc = -3.9499473e-18
+ voffl = 0
+ rgatemod = 0
+ tnjtsswg = 1
+ weta0 = -1.7848176e-8
+ wetab = 1.9534667e-8
+ lpclm = 0
+ cgidl = 1
+ permod = 1
+ ags = -1.2539967
+ nfactor = 1
+ cjd = 0.00144022
+ cit = -0.00036538451
+ cjs = 0.00144022
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 1.38228675e-8
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ pbswd = 0.9
+ pbsws = 0.9
+ voffcv = -0.125
+ wpemod = 1
+ la0 = -4.7253353e-7
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0.001
+ kt1 = -0.16257215
+ kt2 = -0.066291072
+ lk2 = 1.32447077e-9
+ llc = -1.18e-13
+ lln = 0.7
+ lu0 = -5.3790454e-10
+ keta = -0.0061234738
+ mjd = 0.335
+ mjs = 0.335
+ lua = -1.0290148e-16
+ lub = -5.3060964e-27
+ luc = -4.0794824e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pdits = 0
+ pa0 = 9.7298482e-15
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ cigsd = 0.013281
+ pk2 = -2.0891363e-16
+ nigbacc = 10
+ lags = 1.5101544e-6
+ pu0 = 1.1540053e-17
+ dvt0w = 0
+ dvt1w = 0
+ prt = 0
+ dvt2w = 0
+ pua = -1.3867635e-23
+ pub = 2.1855871e-32
+ puc = -2.7646346e-24
+ pud = 0
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 2.0476918e-10
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 1.7313241e-9
+ ub1 = -1.3316629e-18
+ uc1 = 2.2670111e-10
+ kt1l = 0
+ tpb = 0.0016
+ wa0 = -1.7096745e-7
+ ute = -0.86054925
+ web = 6628.3
+ wec = -16935.0
+ pk2we = 0.0
+ wk2 = 4.238936e-9
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ wlc = 0
+ wln = 1
+ wu0 = -2.6120153e-10
+ xgl = -8.2e-9
+ xgw = 0
+ wua = -2.3821198e-16
+ wub = 1.6333936e-25
+ wuc = 4.2583136e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ nigbinv = 2.171
+ lint = 9.7879675e-9
+ tpbswg = 0.001
+ lkt1 = -2.5275191999999998e-8
+ lkt2 = -5.6848171e-9
+ lmax = 4.4741e-7
+ tnoia = 0
+ lmin = 2.1410000000000002e-7
+ lpe0 = 6.44e-8
+ ijthsfwd = 0.01
+ lpeb = 0
+ peta0 = -1.5e-17
+ wketa = -7.8373297e-10
+ minv = -0.33
+ tpbsw = 0.0025
+ lua1 = 4.723388e-17
+ lub1 = -3.0366637e-25
+ luc1 = 1.2420632e-17
+ ptvoff = 5.0195791e-17
+ cjswd = 5.457e-11
+ cjsws = 5.457e-11
+ ndep = 1e+18
+ fnoimod = 1
+ mjswd = 0.01
+ lute = -2.9424109e-8
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ waigsd = 1.9297907e-12
+ lwlc = 0
+ eigbinv = 1.1
+ moin = 5.5538
+ ijthsrev = 0.01
+ nigc = 2.291
+ diomod = 1
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.9367000000000001e-10
+ pku0we = 0.0
+ cjswgs = 1.9367000000000001e-10
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ tvfbsdoff = 0.1
+ pags = -3.3771496e-13
+ scref = 1e-6
+ a0 = 3.1132665
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 72000
+ cf = 7.598099999999999e-11
+ ntox = -1.9260000000000002
+ mjswgd = 0.95
+ ef = 1.15
+ mjswgs = 0.95
+ k1 = 0.30425
+ k2 = -0.0081283305
+ k3 = -2.5823
+ pcit = -9.2716403e-18
+ em = 20000000.0
+ ppdiblc2 = -3.8737293e-16
+ pclm = 1.1689658
+ pigcd = 2.572
+ cigbacc = 0.245
+ ll = -1.18e-13
+ aigsd = 0.0063633912
+ lw = 0
+ u0 = 0.011841230000000001
+ w0 = 0
+ ua = 3.3584387e-10
+ ub = 1.2266958e-18
+ uc = -5.8379738e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 5.6700000000000005e-9
+ ww = 0
+ xw = 3.4e-9
+ tcjswg = 0.00128
+ lvoff = -4.2658924e-9
+ phin = 0.15
+ tnoimod = 0
+ lvsat = 0.00024
+ pkt1 = 6.8355166e-15
+ pkt2 = 2.2627554e-16
+ lvth0 = 3.965357899999999e-9
+ cigbinv = 0.006
+ delta = 0.018814
+ laigc = -1.8017042e-11
+ wvfbsdoff = 0
+ rnoia = 0
+ rnoib = 0
+ lvfbsdoff = 0
+ rbdb = 50
+ pua1 = -2.7108228e-23
+ pkvth0we = 0.0
+ prwb = 0
+ pub1 = 7.1177686e-32
+ prwg = 0
+ puc1 = 8.7727027e-25
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ pketa = 2.0432143e-15
+ version = 4.5
+ ngate = 1.7e+20
+ pute = 1.6065563e-14
+ fprout = 200
+ rdsw = 200
+ ngcon = 1
+ tempmod = 0
+ wpclm = -1.1447315e-8
+ xrcrg1 = 12
+ xrcrg2 = 1
+ vfbsdoff = 0.01
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ aigbacc = 0.012071
+ wtvoff = -1.7507555e-10
+ paramchk = 1
+ rshg = 14.1
+ capmod = 2
+ aigbinv = 0.009974
+ wku0we = 1.5e-11
+ mobmod = 0
+ ijthdfwd = 0.01
+ tvoff = 0.002323434
+ tnom = 25
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ toxe = 2.71e-9
+ toxm = 2.67e-9
+ poxedge = 1
+ ijthdrev = 0.01
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = -5e-10
+ lpdiblc2 = 4.7505822e-10
+ binunit = 2
+ ppclm = 0
+ wags = 5.6744004e-7
+ wcit = 2.107191e-11
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ voff = -0.12137687
+ acde = 0.5
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ vsat = 91103.982
+ wint = 0
+ vth0 = -0.42706475000000005
+ wkt1 = -2.4180539e-8
+ wkt2 = 4.7880041e-9
+ wmax = 5.426e-7
+ dmcgt = 0
+ aigc = 0.0067599617
+ wmin = 2.726e-7
+ tcjsw = 9.34e-5
+ lkvth0we = 3e-12
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ wua1 = 1.9431072e-17
+ wub1 = -1.3369336e-25
+ wuc1 = -7.3645279e-17
+ acnqsmod = 0
+ bigc = 0.0012521
+ bigsd = 0.0003327
+ wute = -7.6140111e-8
+ wwlc = 0
+ wvoff = 1.674468e-9
+ toxref = 3e-9
+ rbodymod = 0
+ cdsc = 0
+ cgbo = 0
+ cgdl = 2.799765e-11
+ cgdo = 2.4628259999999997e-11
+ xtid = 3
+ xtis = 3
+ wvsat = 0.0034765009
+ cgsl = 2.799765e-11
+ cgso = 2.4628259999999997e-11
+ wvth0 = -2.6114098999999997e-9
+ cigc = 0.15259
+ waigc = 1.7749876e-11
+ njtsswg = 6.489
+ lketa = -2.19178e-8
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ ltvoff = -2.3990075e-10
+ xpart = 1
+ ckappad = 0.6
+ wpdiblc2 = 1.1524564e-9
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.0090247504
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ pdiblcb = 0
+ egidl = 0.001
+ pvfbsdoff = 0
+ )

.model pch_ss_29 pmos (
+ level = 54
+ ijthdrev = 0.01
+ ngcon = 1
+ pbswgd = 0.8
+ pbswgs = 0.8
+ wpclm = -1.2079184e-7
+ aigbinv = 0.009974
+ nigc = 2.291
+ igcmod = 1
+ lpdiblc2 = -1.1954251e-9
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ ntox = -1.9260000000000002
+ pcit = -8.1298391e-18
+ pclm = 1.5407845
+ poxedge = 1
+ phin = 0.15
+ lkvth0we = 3e-12
+ pkt1 = -1.21482e-15
+ pkt2 = -1.4992738e-15
+ binunit = 2
+ permod = 1
+ tvoff = 0.00085372815
+ acnqsmod = 0
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ rbdb = 50
+ pua1 = 1.9617826e-23
+ prwb = 0
+ pub1 = -3.1346313e-32
+ prwg = 0
+ puc1 = 1.1713402e-23
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ rbodymod = 0
+ voffcv = -0.125
+ wpemod = 1
+ rdsw = 200
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = -5e-10
+ ppclm = 2.3071337e-14
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ rshg = 14.1
+ wpdiblc2 = -7.3926191e-10
+ tpbswg = 0.001
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ njtsswg = 6.489
+ ptvoff = -3.132788e-17
+ tnom = 25
+ bigsd = 0.0003327
+ waigsd = 1.9297907e-12
+ toxe = 2.71e-9
+ toxm = 2.67e-9
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ wkvth0we = 0.0
+ wvoff = 3.1859801e-10
+ diomod = 1
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.016941733
+ trnqsmod = 0
+ pdiblcb = 0
+ wvsat = 0.0032472346
+ pditsd = 0
+ wvth0 = -7.7669425e-9
+ pditsl = 0
+ cjswgd = 1.9367000000000001e-10
+ pku0we = 0.0
+ cjswgs = 1.9367000000000001e-10
+ waigc = -1.7260908e-11
+ wags = -1.0331048e-6
+ wcit = 1.566053e-11
+ lketa = 7.1935383e-9
+ voff = -0.13201276
+ mjswgd = 0.95
+ mjswgs = 0.95
+ bigbacc = 0.0054401
+ acde = 0.5
+ xpart = 1
+ rgatemod = 0
+ tcjswg = 0.00128
+ vsat = 91523.884
+ wint = 0
+ tnjtsswg = 1
+ vth0 = -0.42462236000000003
+ pvfbsdoff = 0
+ kvth0we = -0.00022
+ egidl = 0.001
+ wkt1 = 1.3972715e-8
+ wkt2 = 1.2965963e-8
+ wmax = 5.426e-7
+ aigc = 0.0067957378
+ wmin = 2.726e-7
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ wua1 = -2.0201942e-16
+ wub1 = 3.5220237e-25
+ wuc1 = -1.2500135e-16
+ bigc = 0.0012521
+ wwlc = 0
+ fprout = 200
+ cdsc = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ a0 = 1.1444157
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ cgbo = 0
+ cgdl = 2.799765e-11
+ cgdo = 2.4628259999999997e-11
+ at = 108550.2
+ xtid = 3
+ cf = 7.598099999999999e-11
+ xtis = 3
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.025395241
+ k3 = -2.5823
+ em = 20000000.0
+ ll = -1.18e-13
+ lw = 0
+ u0 = 0.0102017592
+ cgsl = 2.799765e-11
+ cgso = 2.4628259999999997e-11
+ w0 = 0
+ ua = -3.1599722e-11
+ ub = 1.4008434e-18
+ uc = -1.6299488e-10
+ ud = 0
+ cigc = 0.15259
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 5.6700000000000005e-9
+ ww = 0
+ xw = 3.4e-9
+ pvoff = 8.4546471e-17
+ wtvoff = 2.1129256e-10
+ cdscb = 0
+ cdscd = 0
+ pvsat = -1.6291000000000024e-12
+ wk2we = 0.0
+ pvth0 = 3.2104824e-16
+ drout = 0.56
+ paigc = 3.4373281e-18
+ nfactor = 1
+ capmod = 2
+ voffl = 0
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ wku0we = 1.5e-11
+ dmdg = 0
+ weta0 = -1.7848176e-8
+ wetab = 1.9534667e-8
+ mobmod = 0
+ ags = 5.9031333
+ lpclm = -7.8453093e-8
+ cjd = 0.00144022
+ cit = 0.00015305446
+ cjs = 0.00144022
+ clc = 1e-7
+ cle = 0.6
+ k2we = 5e-5
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 1.38228675e-8
+ ijthsfwd = 0.01
+ k3b = 2.1176
+ dsub = 0.5
+ cgidl = 1
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ dtox = 3.91e-10
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ nigbacc = 10
+ la0 = -5.7105222e-8
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = -0.0067120921
+ kt1 = -0.27233533
+ kt2 = -0.10755274
+ lk2 = 4.9677889e-9
+ eta0 = 0.17962267
+ llc = -1.18e-13
+ lln = 0.7
+ lu0 = -1.919763e-10
+ etab = -0.19577778
+ mjd = 0.335
+ mjs = 0.335
+ lua = -2.5370884e-17
+ lub = -4.2051244e-26
+ luc = 1.7994313e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ pbswd = 0.9
+ pbsws = 0.9
+ njd = 1.02
+ njs = 1.02
+ pa0 = -3.159814e-15
+ ijthsrev = 0.01
+ nsd = 1e+20
+ pbd = 0.75
+ pat = -4.5415452e-10
+ pbs = 0.75
+ pk2 = -2.0710507e-16
+ pu0 = 4.0684676e-18
+ prt = 0
+ pua = 6.5898257e-24
+ pub = -4.9701536e-33
+ puc = -7.066739e-24
+ pud = 0
+ nigbinv = 2.171
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 2.8369875e-9
+ ub1 = -4.0389099e-18
+ uc1 = 4.2708978e-10
+ tpb = 0.0016
+ wa0 = -1.0988104e-7
+ pdits = 0
+ ute = -1
+ wat = 0.0021523911
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 4.2303646e-9
+ cigsd = 0.013281
+ wlc = 0
+ wln = 1
+ wu0 = -2.2579117e-10
+ xgl = -8.2e-9
+ xgw = 0
+ wua = -3.3516677e-16
+ dvt0w = 0
+ wub = 2.9047692e-25
+ wuc = 6.2972257e-17
+ wud = 0
+ dvt1w = 0
+ dvt2w = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ ppdiblc2 = 1.1779633e-17
+ pk2we = 0.0
+ fnoimod = 1
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ eigbinv = 1.1
+ tnoia = 0
+ peta0 = -1.5e-17
+ wketa = 1.4826965e-8
+ tpbsw = 0.0025
+ cjswd = 5.457e-11
+ cjsws = 5.457e-11
+ pkvth0we = 0.0
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ toxref = 3e-9
+ cigbacc = 0.245
+ vfbsdoff = 0.01
+ tnoimod = 0
+ keta = -0.1440919
+ tvfbsdoff = 0.1
+ wtvfbsdoff = 0
+ cigbinv = 0.006
+ ltvoff = 7.0207177e-11
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 9.537856e-11
+ paramchk = 1
+ scref = 1e-6
+ kt1l = 0
+ pigcd = 2.572
+ aigsd = 0.0063633912
+ ltvfbsdoff = 0
+ version = 4.5
+ lvoff = -2.0217201e-9
+ lint = 9.7879675e-9
+ tempmod = 0
+ lkt1 = -2.1151622e-9
+ lkt2 = 3.021395e-9
+ lku0we = 1.8e-11
+ lmax = 2.1410000000000002e-7
+ lvsat = 0.0001514086
+ lmin = 8.833e-8
+ epsrox = 3.9
+ lvth0 = 3.4500146999999996e-9
+ lpe0 = 6.44e-8
+ ijthdfwd = 0.01
+ lpeb = 0
+ delta = 0.018814
+ laigc = -2.5565813e-11
+ aigbacc = 0.012071
+ wvfbsdoff = 0
+ rdsmod = 0
+ lvfbsdoff = 0
+ minv = -0.33
+ rnoia = 0
+ rnoib = 0
+ lua1 = -1.8606111e-16
+ lub1 = 2.6756274e-25
+ luc1 = -2.9861377e-17
+ igbmod = 1
+ ndep = 1e+18
+ ptvfbsdoff = 0
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ lwlc = 0
+ pketa = -1.250643e-15
+ ngate = 1.7e+20
+ moin = 5.5538
+ )

.model pch_ss_30 pmos (
+ level = 54
+ ijthdrev = 0.01
+ ngcon = 1
+ pbswgd = 0.8
+ pbswgs = 0.8
+ wpclm = 4.9341412e-7
+ aigbinv = 0.009974
+ nigc = 2.291
+ igcmod = 1
+ lpdiblc2 = 0
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ ntox = -1.9260000000000002
+ pcit = 1.0726434999999998e-17
+ pclm = 0.08631615
+ paigsd = 8.4526218e-25
+ poxedge = 1
+ phin = 0.15
+ lkvth0we = 3e-12
+ pkt1 = -1.7124191e-15
+ pkt2 = 2.1480498e-17
+ binunit = 2
+ permod = 1
+ tvoff = 0.0012365685
+ acnqsmod = 0
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ rbdb = 50
+ pua1 = 4.1792962e-25
+ prwb = 0
+ pub1 = 6.1746384e-33
+ prwg = 0
+ puc1 = 2.9246063e-24
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ rbodymod = 0
+ voffcv = -0.125
+ wpemod = 1
+ rdsw = 200
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = -9.065883199999999e-9
+ letab = 1.7579973e-8
+ ppclm = -3.4664022e-14
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ rshg = 14.1
+ wpdiblc2 = -6.1394667e-10
+ tpbswg = 0.001
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ njtsswg = 6.489
+ ptvoff = 2.0376593e-17
+ tnom = 25
+ bigsd = 0.0003327
+ waigsd = 1.9297817e-12
+ toxe = 2.71e-9
+ toxm = 2.67e-9
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ wkvth0we = 0.0
+ wvoff = -2.8254962e-9
+ diomod = 1
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.0042244444
+ trnqsmod = 0
+ pdiblcb = 0
+ wvsat = 0.023310745
+ pditsd = 0
+ wvth0 = 1.4897438999999999e-9
+ pditsl = 0
+ cjswgd = 1.9367000000000001e-10
+ pku0we = 0.0
+ cjswgs = 1.9367000000000001e-10
+ waigc = 7.1461687e-12
+ wags = -1.0331048e-6
+ wcit = -1.8493752e-10
+ lketa = -1.1878561e-8
+ voff = -0.12098873
+ mjswgd = 0.95
+ mjswgs = 0.95
+ bigbacc = 0.0054401
+ acde = 0.5
+ xpart = 1
+ rgatemod = 0
+ tcjswg = 0.00128
+ vsat = 39425.539000000004
+ wint = 0
+ tnjtsswg = 1
+ vth0 = -0.39778691000000005
+ pvfbsdoff = 0
+ kvth0we = -0.00022
+ egidl = 0.001
+ wkt1 = 1.9266322e-8
+ wkt2 = -3.2122744e-9
+ wmax = 5.426e-7
+ aigc = 0.0067006504
+ wmin = 2.726e-7
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ wua1 = 2.2347963e-18
+ wub1 = -4.6956688e-26
+ wuc1 = -3.1503526e-17
+ bigc = 0.0012521
+ wwlc = 0
+ fprout = 200
+ cdsc = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ a0 = 3.9744452
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ cgbo = 0
+ cgdl = 2.799765e-11
+ cgdo = 2.4628259999999997e-11
+ at = 69068.642
+ xtid = 3
+ cf = 7.598099999999999e-11
+ xtis = 3
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.022825095
+ k3 = -2.5823
+ em = 20000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.0043656963
+ cgsl = 2.799765e-11
+ cgso = 2.4628259999999997e-11
+ w0 = 0
+ ua = -9.2439852e-11
+ ub = -1.6232125e-18
+ uc = 5.3507127e-11
+ ud = 0
+ cigc = 0.15259
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 5.6700000000000005e-9
+ ww = 0
+ xw = 3.4e-9
+ pvoff = 3.8009132e-16
+ wtvoff = -3.3875503e-10
+ cdscb = 0
+ cdscd = 0
+ pvsat = -1.8875991e-9
+ wk2we = 0.0
+ pvth0 = -5.490808600000001e-16
+ drout = 0.56
+ paigc = 1.1430629e-18
+ nfactor = 1
+ capmod = 2
+ voffl = 0
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ wku0we = 1.5e-11
+ dmdg = 0
+ weta0 = -5.5215839e-8
+ wetab = 4.6876459e-8
+ mobmod = 0
+ ags = 5.9031333
+ lpclm = 5.8266931e-8
+ cjd = 0.00144022
+ cit = -0.00017317562
+ cjs = 0.00144022
+ clc = 1e-7
+ cle = 0.6
+ k2we = 5e-5
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 4.0349e-9
+ ijthsfwd = 0.01
+ k3b = 2.1176
+ dsub = 0.5
+ cgidl = 1
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ dtox = 3.91e-10
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ nigbacc = 10
+ la0 = -3.23128e-7
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = -0.0030008257
+ kt1 = -0.32608492
+ kt2 = -0.08284588
+ lk2 = 4.726195200000001e-9
+ eta0 = 0.27074908
+ llc = 0
+ lln = 1
+ lu0 = 3.5661361999999997e-10
+ etab = -0.38279877
+ mjd = 0.335
+ mjs = 0.335
+ lua = -1.9651912e-17
+ lub = 2.4221001e-25
+ luc = -2.356876e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ pbswd = 0.9
+ pbsws = 0.9
+ njd = 1.02
+ njs = 1.02
+ pa0 = 9.1746422e-14
+ laigsd = -3.0625433e-18
+ ijthsrev = 0.01
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 6.7620954e-11
+ pbs = 0.75
+ pk2 = 2.5170462e-16
+ pu0 = -8.2666616e-17
+ prt = 0
+ pua = 3.032424e-23
+ pub = -9.6166295e-32
+ puc = -2.0363205e-24
+ pud = 0
+ nigbinv = 2.171
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = -2.7998083e-10
+ ub1 = 8.7083504e-19
+ uc1 = 1.8820988e-11
+ tpb = 0.0016
+ wa0 = -1.1195219e-6
+ pdits = 0
+ ute = -1
+ wat = -0.0033984119
+ web = 6628.3
+ wec = -16935.0
+ wk2 = -6.5058945e-10
+ cigsd = 0.013281
+ wlc = 0
+ wln = 1
+ wu0 = 6.9692249e-10
+ xgl = -8.2e-9
+ xgw = 0
+ wua = -5.8766054e-16
+ dvt0w = 0
+ wub = 1.2606486e-24
+ wuc = 9.4571662e-18
+ wud = 0
+ dvt1w = 0
+ dvt2w = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ ppdiblc2 = 0
+ pk2we = 0.0
+ fnoimod = 1
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ eigbinv = 1.1
+ tnoia = 0
+ peta0 = 3.4975603e-15
+ petab = -2.5701285e-15
+ wketa = -3.6489897e-8
+ tpbsw = 0.0025
+ cjswd = 5.457e-11
+ cjsws = 5.457e-11
+ pkvth0we = 0.0
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ toxref = 3e-9
+ cigbacc = 0.245
+ vfbsdoff = 0.01
+ tnoimod = 0
+ keta = 0.058802768
+ tvfbsdoff = 0.1
+ wtvfbsdoff = 0
+ cigbinv = 0.006
+ ltvoff = 3.4220189e-11
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 1.26044219e-10
+ paramchk = 1
+ scref = 1e-6
+ kt1l = 0
+ pigcd = 2.572
+ aigsd = 0.0063633912
+ ltvfbsdoff = 0
+ version = 4.5
+ lvoff = -3.0579783e-9
+ lint = 0
+ tempmod = 0
+ lkt1 = 2.9372998999999997e-9
+ lkt2 = 6.989501e-10
+ lku0we = 1.8e-11
+ lmax = 8.833e-8
+ lvsat = 0.0050486503000000005
+ lmin = 5.233e-8
+ epsrox = 3.9
+ lvth0 = 9.274851999999998e-10
+ lpe0 = 6.44e-8
+ ijthdfwd = 0.01
+ lpeb = 0
+ delta = 0.018814
+ laigc = -1.6627591e-11
+ aigbacc = 0.012071
+ wvfbsdoff = 0
+ rdsmod = 0
+ lvfbsdoff = 0
+ minv = -0.33
+ rnoia = 0
+ rnoib = 0
+ lua1 = 1.0693391e-16
+ lub1 = -1.9395329e-25
+ luc1 = 8.5158894e-18
+ igbmod = 1
+ ndep = 1e+18
+ ptvfbsdoff = 0
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ lwlc = 0
+ pketa = 3.573142e-15
+ ngate = 1.7e+20
+ moin = 5.5538
+ )

.model pch_ss_31 pmos (
+ level = 54
+ paigc = -3.8652128e-18
+ voff = -0.11425646
+ nigbacc = 10
+ ags = 5.9031333
+ acde = 0.5
+ ppdiblc2 = 0
+ voffl = 0
+ cjd = 0.00144022
+ cit = -0.0111997498
+ cjs = 0.00144022
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ vsat = 280400.89
+ dlc = 4.0349e-9
+ wint = 0
+ k3b = 2.1176
+ vth0 = -0.28618022000000004
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ weta0 = 4.5369198e-8
+ wkt1 = -9.053012e-8
+ wkt2 = -4.5663135e-8
+ wetab = 2.1214781e-8
+ wmax = 5.426e-7
+ aigc = 0.0065523001
+ wmin = 2.726e-7
+ lpclm = -1.6067206e-7
+ permod = 1
+ nigbinv = 2.171
+ la0 = 2.2449695e-9
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 5.472133000000007e-5
+ kt1 = -0.078489325
+ kt2 = 0.051187672
+ lk2 = 5.823110100000001e-9
+ llc = 0
+ lln = 1
+ cgidl = 1
+ lu0 = -6.3649203e-10
+ mjd = 0.335
+ mjs = 0.335
+ lua = -5.2618623e-17
+ lub = -3.527729e-25
+ luc = -2.0280652e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ wua1 = 2.8402308e-15
+ njs = 1.02
+ wub1 = -3.9062366e-24
+ wuc1 = 2.0276364e-16
+ pa0 = -4.432942e-14
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 1.8264736e-9
+ pbs = 0.75
+ pk2 = -1.1995676e-16
+ pu0 = 2.2577126e-16
+ bigc = 0.0012521
+ prt = 0
+ pua = 1.5923531e-23
+ pub = 1.0433766599999999e-31
+ puc = 3.3504384e-24
+ pud = 0
+ wwlc = 0
+ pkvth0we = 0.0
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = -3.345352e-9
+ ub1 = 3.9080279e-18
+ uc1 = 1.4308247e-10
+ tpb = 0.0016
+ voffcv = -0.125
+ wpemod = 1
+ pbswd = 0.9
+ pbsws = 0.9
+ wa0 = 1.2266134e-6
+ cdsc = 0
+ ute = -1
+ wat = -0.033723458
+ web = 6628.3
+ wec = -16935.0
+ fnoimod = 1
+ wk2 = 5.7573654e-9
+ wlc = 0
+ cgbo = 0
+ wln = 1
+ cgdl = 2.799765e-11
+ cgdo = 2.4628259999999997e-11
+ wu0 = -4.6209719e-9
+ xtid = 3
+ xgl = -8.2e-9
+ xtis = 3
+ xgw = 0
+ wua = -3.3937245e-16
+ wub = -2.1963169e-24
+ wuc = -8.3417988e-17
+ wud = 0
+ eigbinv = 1.1
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ cgsl = 2.799765e-11
+ cgso = 2.4628259999999997e-11
+ vfbsdoff = 0.01
+ cigc = 0.15259
+ pdits = 0
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ paramchk = 1
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ tpbswg = 0.001
+ cigbacc = 0.245
+ tnoia = 0
+ k2we = 5e-5
+ tnoimod = 0
+ ijthdfwd = 0.01
+ peta0 = -2.3363718000000002e-15
+ dsub = 0.5
+ petab = -1.0817512e-15
+ dtox = 3.91e-10
+ wketa = 7.0696889e-8
+ ptvoff = -1.3332507e-17
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ tpbsw = 0.0025
+ waigsd = 1.9297962e-12
+ cigbinv = 0.006
+ cjswd = 5.457e-11
+ cjsws = 5.457e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ eta0 = 0.012687945
+ etab = -0.23454709
+ diomod = 1
+ ijthdrev = 0.01
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.9367000000000001e-10
+ pku0we = 0.0
+ version = 4.5
+ cjswgs = 1.9367000000000001e-10
+ lpdiblc2 = 0
+ tempmod = 0
+ tvfbsdoff = 0.1
+ aigbacc = 0.012071
+ mjswgd = 0.95
+ mjswgs = 0.95
+ scref = 1e-6
+ tcjswg = 0.00128
+ pigcd = 2.572
+ aigsd = 0.0063633912
+ lvoff = -3.4484499e-9
+ lkvth0we = 3e-12
+ aigbinv = 0.009974
+ lvsat = -0.0089279093
+ lvth0 = -5.5457143e-9
+ delta = 0.018814
+ wvfbsdoff = 0
+ laigc = -8.0232722e-12
+ lvfbsdoff = 0
+ rnoia = 0
+ rnoib = 0
+ acnqsmod = 0
+ fprout = 200
+ pketa = -2.6436916e-15
+ ngate = 1.7e+20
+ xrcrg1 = 12
+ xrcrg2 = 1
+ rbodymod = 0
+ ngcon = 1
+ wpclm = -6.9641486e-7
+ poxedge = 1
+ gbmin = 1e-12
+ wtvoff = 2.4243635e-10
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ keta = -0.44725926
+ binunit = 2
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 7.655849499999999e-10
+ capmod = 2
+ kt1l = 0
+ wku0we = 1.5e-11
+ wpdiblc2 = -6.1394667e-10
+ mobmod = 0
+ lint = 0
+ lkt1 = -1.1423245000000001e-8
+ lkt2 = -7.0749959e-9
+ lmax = 5.233e-8
+ lmin = 4.333e-8
+ a0 = -1.6354335
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 16386.797
+ cf = 7.598099999999999e-11
+ lpe0 = 6.44e-8
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.041737421
+ k3 = -2.5823
+ em = 20000000.0
+ lpeb = 0
+ ll = 0
+ lw = 0
+ u0 = 0.021488207
+ w0 = 0
+ tvoff = 0.0019328761
+ ua = 4.7595173e-10
+ ub = 8.6351132e-18
+ uc = 4.7837975e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 5.6700000000000005e-9
+ ww = 0
+ xw = 3.4e-9
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ minv = -0.33
+ xjbvd = 1
+ xjbvs = 1
+ lua1 = 2.8472544e-16
+ lub1 = -3.7011047e-25
+ lk2we = 0.0
+ luc1 = 1.3087235e-18
+ ndep = 1e+18
+ wkvth0we = 0.0
+ lwlc = 0
+ moin = 5.5538
+ ku0we = -0.0007
+ trnqsmod = 0
+ nigc = 2.291
+ beta0 = 13.32
+ leta0 = 5.9016629e-9
+ letab = 8.9813755e-9
+ ppclm = 3.4346058e-14
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ njtsswg = 6.489
+ ntox = -1.9260000000000002
+ pcit = -1.9387061000000002e-16
+ pclm = 3.8611263
+ rgatemod = 0
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ tnjtsswg = 1
+ dmcgt = 0
+ ckappad = 0.6
+ phin = 0.15
+ ckappas = 0.6
+ tcjsw = 9.34e-5
+ pdiblc1 = 0
+ pdiblc2 = 0.0042244444
+ pdiblcb = 0
+ pkt1 = 4.6557745e-15
+ pkt2 = 2.4836304e-15
+ bigsd = 0.0003327
+ toxref = 3e-9
+ rbdb = 50
+ pua1 = -1.6418584e-22
+ prwb = 0
+ pub1 = 2.3001287e-31
+ prwg = 0
+ puc1 = -1.0662889e-23
+ wtvfbsdoff = 0
+ bigbacc = 0.0054401
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ wvoff = 3.9335999e-9
+ rdsw = 200
+ wvsat = -0.056506619
+ kvth0we = -0.00022
+ ltvfbsdoff = 0
+ wvth0 = -8.835119e-9
+ waigc = 9.3495749e-11
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ ltvoff = -6.1656569e-12
+ lketa = 1.7473037e-8
+ xpart = 1
+ rshg = 14.1
+ pvfbsdoff = 0
+ egidl = 0.001
+ ptvfbsdoff = 0
+ lku0we = 1.8e-11
+ epsrox = 3.9
+ ijthsfwd = 0.01
+ rdsmod = 0
+ igbmod = 1
+ tnom = 25
+ toxe = 2.71e-9
+ toxm = 2.67e-9
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ nfactor = 1
+ pbswgd = 0.8
+ pbswgs = 0.8
+ ijthsrev = 0.01
+ igcmod = 1
+ pvoff = -1.1936247999999998e-17
+ cdscb = 0
+ cdscd = 0
+ wags = -1.0331048e-6
+ pvsat = 2.7418061e-9
+ wk2we = 0.0
+ pvth0 = 4.9761460000000076e-17
+ wcit = 3.34259593e-9
+ drout = 0.56
+ )

.model pch_ss_32 pmos (
+ level = 54
+ tvoff = 0.0050068134
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ voffcv = -0.125
+ wpemod = 1
+ njtsswg = 6.489
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = 4.4376338000000005e-9
+ ckappad = 0.6
+ letab = 1.8240871e-9
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.0042244444
+ pdiblcb = 0
+ keta = -0.10111506
+ ppclm = 1.7398739e-15
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = -4.892745e-10
+ kt1l = 0
+ tpbswg = 0.001
+ bigbacc = 0.0054401
+ lint = 0
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ lkt1 = -1.4409032e-8
+ lkt2 = 2.2261728e-10
+ lmax = 4.333e-8
+ kvth0we = -0.00022
+ lmin = 3.6e-8
+ lpe0 = 6.44e-8
+ ijthsfwd = 0.01
+ lpeb = 0
+ ptvoff = 3.2244316e-17
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ waigsd = 1.9257033e-12
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ minv = -0.33
+ bigsd = 0.0003327
+ lua1 = -1.7116539e-16
+ lub1 = 1.8575894699999999e-25
+ luc1 = 2.2025561e-17
+ ndep = 1e+18
+ diomod = 1
+ lwlc = 0
+ wvoff = 1.094003e-8
+ moin = 5.5538
+ ijthsrev = 0.01
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.9367000000000001e-10
+ pku0we = 0.0
+ cjswgs = 1.9367000000000001e-10
+ nigc = 2.291
+ wvsat = -0.013751414
+ wvth0 = -2.4112669999999983e-9
+ waigc = 1.753535e-10
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ mjswgd = 0.95
+ mjswgs = 0.95
+ lketa = 5.1197136e-10
+ tcjswg = 0.00128
+ xpart = 1
+ ntox = -1.9260000000000002
+ ppdiblc2 = 0
+ pcit = 2.5525304e-16
+ pclm = 0.85281474
+ pvfbsdoff = 0
+ nfactor = 1
+ egidl = 0.001
+ phin = 0.15
+ pkt1 = 2.438466e-15
+ pkt2 = -1.2154904e-16
+ fprout = 200
+ pkvth0we = 0.0
+ rbdb = 50
+ pua1 = 5.9435365e-23
+ prwb = 0
+ pub1 = -6.897475440000001e-32
+ prwg = 0
+ puc1 = -3.4884574e-24
+ xrcrg1 = 12
+ xrcrg2 = 1
+ nigbacc = 10
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ rdsw = 200
+ wtvoff = -6.8770288e-10
+ vfbsdoff = 0.01
+ pvoff = -3.5525133e-16
+ ags = 5.9031333
+ nigbinv = 2.171
+ cdscb = 0
+ cdscd = 0
+ cjd = 0.00144022
+ cit = 0.0144096321
+ cjs = 0.00144022
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ pvsat = 6.468032699999999e-10
+ dlc = 4.0349e-9
+ wk2we = 0.0
+ pvth0 = -2.650058000000001e-16
+ k3b = 2.1176
+ dwb = 0
+ drout = 0.56
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ capmod = 2
+ paramchk = 1
+ paigc = -7.8762427e-18
+ wku0we = 1.5e-11
+ rshg = 14.1
+ voffl = 0
+ la0 = -2.1218621e-7
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0.012168675999999998
+ mobmod = 0
+ kt1 = -0.017554887
+ kt2 = -0.09774321
+ lk2 = 4.457225800000001e-9
+ llc = 0
+ lln = 1
+ lu0 = -2.385917e-10
+ mjd = 0.335
+ mjs = 0.335
+ lua = 4.1444844e-17
+ lub = -1.0372545e-25
+ luc = -1.4956542e-17
+ lud = 0
+ lwc = 0
+ weta0 = 3.13360382e-8
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ wetab = -5.613608e-9
+ njs = 1.02
+ pa0 = 5.0455005e-14
+ fnoimod = 1
+ nsd = 1e+20
+ pbd = 0.75
+ pat = -2.6671169e-9
+ pbs = 0.75
+ pk2 = 3.3742201e-16
+ lpclm = -1.3264792e-8
+ pu0 = 1.5059926e-16
+ eigbinv = 1.1
+ prt = 0
+ pua = 9.2877876e-24
+ pub = 1.5765362e-32
+ puc = 3.1614905e-24
+ pud = 0
+ ijthdfwd = 0.01
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 5.9585425e-9
+ ub1 = -7.436245890000001e-18
+ uc1 = -2.7971012e-10
+ cgidl = 1
+ tpb = 0.0016
+ wa0 = -7.0776268e-7
+ ute = -1
+ wat = 0.057982464
+ web = 6628.3
+ wec = -16935.0
+ wk2 = -3.5768953e-9
+ wlc = 0
+ wln = 1
+ wu0 = -3.0868494e-9
+ tnom = 25
+ xgl = -8.2e-9
+ xgw = 0
+ wua = -2.0394912e-16
+ wub = -3.8871908000000002e-25
+ wuc = -7.9561907e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ toxe = 2.71e-9
+ toxm = 2.67e-9
+ laigsd = -3.6731852e-16
+ pbswd = 0.9
+ pbsws = 0.9
+ ijthdrev = 0.01
+ cigbacc = 0.245
+ lpdiblc2 = 0
+ pdits = 0
+ wags = -1.0331048e-6
+ cigsd = 0.013281
+ tnoimod = 0
+ dvt0w = 0
+ dvt1w = 0
+ wcit = -5.8231926000000004e-9
+ dvt2w = 0
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ a0 = 2.7407131
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = -230836.79
+ cf = 7.598099999999999e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.013862232
+ k3 = -2.5823
+ em = 20000000.0
+ voff = -0.14966725
+ ll = 0
+ lw = 0
+ u0 = 0.013367793000000001
+ w0 = 0
+ cigbinv = 0.006
+ acde = 0.5
+ ua = -1.4437109e-9
+ ub = 3.5525119e-18
+ uc = 3.1168444e-10
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 5.6700000000000005e-9
+ ww = 0
+ xw = 3.4e-9
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ vsat = 180673.32
+ wint = 0
+ vth0 = -0.36502203
+ wkt1 = -4.5278925e-8
+ wkt2 = 7.5037926e-9
+ wtvfbsdoff = 0
+ wmax = 5.426e-7
+ aigc = 0.006152944
+ wmin = 2.726e-7
+ lkvth0we = 3e-12
+ tnoia = 0
+ version = 4.5
+ tempmod = 0
+ peta0 = -1.64874789e-15
+ ltvfbsdoff = 0
+ petab = 2.3283989e-16
+ wketa = 1.3494424e-8
+ wua1 = -1.7234672e-15
+ wub1 = 2.19555176e-24
+ wuc1 = 5.6346661e-17
+ tpbsw = 0.0025
+ acnqsmod = 0
+ toxref = 3e-9
+ bigc = 0.0012521
+ aigbacc = 0.012071
+ cjswd = 5.457e-11
+ cjsws = 5.457e-11
+ wwlc = 0
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ rbodymod = 0
+ cdsc = 0
+ cgbo = 0
+ cgdl = 2.799765e-11
+ cgdo = 2.4628259999999997e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 2.799765e-11
+ cgso = 2.4628259999999997e-11
+ cigc = 0.15259
+ aigbinv = 0.009974
+ tvfbsdoff = 0.1
+ ptvfbsdoff = 0
+ ltvoff = -1.5678858e-10
+ scref = 1e-6
+ pigcd = 2.572
+ aigsd = 0.0063633987
+ wpdiblc2 = -6.1394667e-10
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ lku0we = 1.8e-11
+ lvoff = -1.7133213e-9
+ epsrox = 3.9
+ lvsat = -0.0040412681
+ poxedge = 1
+ lvth0 = -1.6824604e-9
+ k2we = 5e-5
+ wvfbsdoff = 0
+ rdsmod = 0
+ lvfbsdoff = 0
+ delta = 0.018814
+ dsub = 0.5
+ dtox = 3.91e-10
+ laigc = 1.1545174e-11
+ igbmod = 1
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ binunit = 2
+ rnoia = 0
+ rnoib = 0
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ pbswgd = 0.8
+ wkvth0we = 0.0
+ pbswgs = 0.8
+ eta0 = 0.04256602999999999
+ pketa = 1.5922924e-16
+ etab = -0.088479977
+ ngate = 1.7e+20
+ ngcon = 1
+ igcmod = 1
+ wpclm = -3.0982532e-8
+ trnqsmod = 0
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ paigsd = 2.0055591e-22
+ rgatemod = 0
+ tnjtsswg = 1
+ permod = 1
+ )

.model pch_ss_33 pmos (
+ level = 54
+ version = 4.5
+ pdits = 0
+ cigsd = 0.013281
+ tempmod = 0
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ tpbswg = 0.001
+ rshg = 14.1
+ aigbacc = 0.012071
+ wpdiblc2 = 3.3638075e-10
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ tnoia = 0
+ ptvoff = 0
+ aigbinv = 0.009974
+ peta0 = -1.5e-17
+ waigsd = 1.9846811e-12
+ wketa = -1.9384664e-9
+ tpbsw = 0.0025
+ tnom = 25
+ diomod = 1
+ cjswd = 5.457e-11
+ cjsws = 5.457e-11
+ toxe = 2.71e-9
+ toxm = 2.67e-9
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ wkvth0we = 0.0
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.9367000000000001e-10
+ pku0we = 0.0
+ cjswgs = 1.9367000000000001e-10
+ trnqsmod = 0
+ tvfbsdoff = 0.1
+ poxedge = 1
+ mjswgd = 0.95
+ wags = 5.1942014e-9
+ mjswgs = 0.95
+ tcjswg = 0.00128
+ binunit = 2
+ scref = 1e-6
+ voff = -0.10372023
+ acde = 0.5
+ pigcd = 2.572
+ aigsd = 0.0063632583
+ rgatemod = 0
+ vsat = 108525.44
+ tnjtsswg = 1
+ wint = 0
+ vth0 = -0.39987116
+ lvoff = 0
+ wkt1 = -3.0503659e-9
+ wkt2 = -7.2833333e-10
+ wmax = 2.726e-7
+ aigc = 0.0068302204
+ wmin = 1.08e-7
+ lvsat = 0.00024
+ lvth0 = -6e-10
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ delta = 0.018814
+ wua1 = -5.5326541e-17
+ wub1 = -1.0689498e-25
+ wuc1 = -1.2119467e-17
+ fprout = 200
+ rnoia = 0
+ rnoib = 0
+ bigc = 0.0012521
+ wute = -7.6523556e-8
+ xrcrg1 = 12
+ xrcrg2 = 1
+ wwlc = 0
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ ngate = 1.7e+20
+ ngcon = 1
+ cdsc = 0
+ wpclm = 7.1298978e-9
+ cgbo = 0
+ cgdl = 2.799765e-11
+ wtvoff = -7.3630015e-11
+ cgdo = 2.4628259999999997e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 2.799765e-11
+ cgso = 2.4628259999999997e-11
+ cigc = 0.15259
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ capmod = 2
+ wku0we = 1.5e-11
+ mobmod = 0
+ njtsswg = 6.489
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ k2we = 5e-5
+ ckappad = 0.6
+ ckappas = 0.6
+ ijthsfwd = 0.01
+ pdiblc1 = 0
+ pdiblc2 = 0.0015492917
+ dsub = 0.5
+ pdiblcb = 0
+ dtox = 3.91e-10
+ tvoff = 0.0025423547
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ eta0 = 0.10792519
+ etab = -0.13555556
+ ijthsrev = 0.01
+ ku0we = -0.0007
+ bigbacc = 0.0054401
+ beta0 = 13.32
+ leta0 = -5e-10
+ wtvfbsdoff = 0
+ kvth0we = -0.00022
+ ppclm = 0
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ dlcig = 2.5e-9
+ lintnoi = -5e-9
+ bgidl = 1834800000.0
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ ltvfbsdoff = 0
+ ppdiblc2 = 0
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ toxref = 3e-9
+ bigsd = 0.0003327
+ ptvfbsdoff = 0
+ pkvth0we = 0.0
+ wvoff = 1.4142431e-9
+ a0 = 2.5876667
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 72000
+ cf = 7.598099999999999e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.015389268
+ k3 = -2.5823
+ em = 20000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.0098471852
+ w0 = 0
+ ua = -1.9215717e-10
+ ub = 1.2747184e-18
+ uc = -1.7585185e-12
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 5.6700000000000005e-9
+ ww = 0
+ xw = 3.4e-9
+ wvsat = -0.0013318206
+ nfactor = 1
+ wvth0 = -6.0254372e-9
+ vfbsdoff = 0.01
+ waigc = 1.6569661e-12
+ keta = 0.02482765
+ ltvoff = 0
+ jswd = 3.69e-13
+ lketa = 0
+ jsws = 3.69e-13
+ paramchk = 1
+ lcit = 0
+ xpart = 1
+ pvfbsdoff = 0
+ kt1l = 0
+ lku0we = 1.8e-11
+ nigbacc = 10
+ egidl = 0.001
+ epsrox = 3.9
+ lint = 6.5375218e-9
+ lkt1 = -1e-9
+ lmax = 2.001e-5
+ lmin = 8.99743e-6
+ rdsmod = 0
+ ijthdfwd = 0.01
+ lpe0 = 6.44e-8
+ igbmod = 1
+ lpeb = 0
+ nigbinv = 2.171
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ minv = -0.33
+ pbswgd = 0.8
+ pbswgs = 0.8
+ ndep = 1e+18
+ ags = 0.89683683
+ lwlc = 0
+ igcmod = 1
+ moin = 5.5538
+ ijthdrev = 0.01
+ cjd = 0.00144022
+ cit = 5e-6
+ cjs = 0.00144022
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 1.0572421799999999e-8
+ nigc = 2.291
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ lpdiblc2 = 0
+ fnoimod = 1
+ pvoff = 2.5e-17
+ eigbinv = 1.1
+ cdscb = 0
+ cdscd = 0
+ la0 = 0
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ jsd = 1.5e-7
+ pvsat = -5e-11
+ jss = 1.5e-7
+ lat = 0.001
+ kt1 = -0.17197747
+ lk2 = 4e-10
+ kt2 = -0.050761111
+ wk2we = 0.0
+ pvth0 = -7e-17
+ llc = 0
+ lln = 1
+ lu0 = 5e-12
+ drout = 0.56
+ mjd = 0.335
+ mjs = 0.335
+ lub = 0
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 0
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ pk2 = 0
+ pu0 = 0
+ ntox = -1.9260000000000002
+ voffl = 0
+ prt = 0
+ pub = 0
+ pcit = 0
+ pud = 0
+ pclm = 1.101657
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 9.8162749e-10
+ ub1 = -3.8648101e-20
+ uc1 = 8.1681111e-11
+ tpb = 0.0016
+ weta0 = 1.9403288999999997e-9
+ permod = 1
+ wa0 = 4.8944e-8
+ wetab = 2.9133333e-9
+ ute = -0.81574074
+ phin = 0.15
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 3.9065138e-9
+ lkvth0we = 3e-12
+ lpclm = 0
+ wlc = 0
+ wln = 1
+ wu0 = 5.8460889e-11
+ xgl = -8.2e-9
+ xgw = 0
+ wua = -4.8614483e-17
+ wub = 8.106039e-27
+ wuc = 3.3309111e-18
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ cigbacc = 0.245
+ pkt1 = 0
+ cgidl = 1
+ tnoimod = 0
+ acnqsmod = 0
+ voffcv = -0.125
+ wpemod = 1
+ rbdb = 50
+ prwb = 0
+ prwg = 0
+ rbpb = 50
+ rbpd = 50
+ cigbinv = 0.006
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ pbswd = 0.9
+ rbodymod = 0
+ pbsws = 0.9
+ rdsw = 200
+ )

.model pch_ss_34 pmos (
+ level = 54
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ nfactor = 1
+ ptvoff = -5.393716e-17
+ k2we = 5e-5
+ waigsd = 1.9861139e-12
+ ijthdfwd = 0.01
+ dsub = 0.5
+ dtox = 3.91e-10
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ diomod = 1
+ bigsd = 0.0003327
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.9367000000000001e-10
+ pku0we = 0.0
+ cjswgs = 1.9367000000000001e-10
+ eta0 = 0.10792519
+ wvoff = 1.3100722e-9
+ etab = -0.13555556
+ ijthdrev = 0.01
+ nigbacc = 10
+ wvsat = -0.0013318206
+ wvth0 = -6.1211131e-9
+ lpdiblc2 = 6.2970633e-9
+ waigc = 1.4905459e-12
+ mjswgd = 0.95
+ mjswgs = 0.95
+ tcjswg = 0.00128
+ nigbinv = 2.171
+ lketa = -5.5366519e-8
+ pvfbsdoff = 0
+ xpart = 1
+ egidl = 0.001
+ lkvth0we = 3e-12
+ fnoimod = 1
+ ags = 0.84380759
+ eigbinv = 1.1
+ fprout = 200
+ cjd = 0.00144022
+ cit = 5e-6
+ cjs = 0.00144022
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ acnqsmod = 0
+ dlc = 1.0572421799999999e-8
+ xrcrg1 = 12
+ xrcrg2 = 1
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ rbodymod = 0
+ la0 = -3.9401851e-7
+ wtvoff = -6.7630331e-11
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0.001
+ kt1 = -0.17107141
+ kt2 = -0.050597496
+ lk2 = 5.931940300000001e-9
+ llc = 0
+ lln = 1
+ lu0 = 1.00178999e-9
+ mjd = 0.335
+ mjs = 0.335
+ lua = -7.2048384e-17
+ lub = 4.3514377e-25
+ luc = 1.4270275e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = -3.1655381e-14
+ pvoff = 9.6149624e-16
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ pk2 = 9.285497e-17
+ keta = 0.030986328
+ pu0 = 3.0504276e-17
+ prt = 0
+ cdscb = 0
+ cdscd = 0
+ pua = 2.7735079e-23
+ pub = -4.2717478e-32
+ puc = 1.20866e-25
+ pud = 0
+ cigbacc = 0.245
+ capmod = 2
+ pvsat = -5e-11
+ rsh = 15.2
+ wk2we = 0.0
+ tcj = 0.000832
+ ua1 = 8.0734953e-10
+ pvth0 = 7.901263899999999e-16
+ ub1 = 2.6826436e-19
+ uc1 = 8.9789043e-11
+ drout = 0.56
+ lags = 4.7673289e-7
+ wku0we = 1.5e-11
+ tpb = 0.0016
+ wa0 = 5.2465177e-8
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ ute = -0.817454
+ paigc = 1.4961177e-18
+ lcit = 0
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 3.8961851e-9
+ tnoimod = 0
+ mobmod = 0
+ wlc = 0
+ wln = 1
+ wu0 = 5.5067755e-11
+ xgl = -8.2e-9
+ xgw = 0
+ kt1l = 0
+ wua = -5.1699586e-17
+ wub = 1.2857705e-26
+ wuc = 3.3174666e-18
+ wud = 0
+ voffl = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ wpdiblc2 = 3.5925269e-10
+ cigbinv = 0.006
+ weta0 = 1.9403288999999997e-9
+ wetab = 2.9133333e-9
+ lint = 6.5375218e-9
+ lpclm = 0
+ lkt1 = -9.1454893e-9
+ lkt2 = -1.4709041e-9
+ lmax = 8.99743e-6
+ lmin = 8.974099999999999e-7
+ lpe0 = 6.44e-8
+ cgidl = 1
+ lpeb = 0
+ version = 4.5
+ tempmod = 0
+ minv = -0.33
+ wtvfbsdoff = 0
+ laigsd = -1.8524358e-14
+ lua1 = 1.5667589e-15
+ lub1 = -2.759143e-24
+ luc1 = -7.2890309e-17
+ ndep = 1e+18
+ wkvth0we = 0.0
+ lute = 1.5402209e-8
+ lwlc = 0
+ pbswd = 0.9
+ pbsws = 0.9
+ moin = 5.5538
+ aigbacc = 0.012071
+ ltvfbsdoff = 0
+ trnqsmod = 0
+ nigc = 2.291
+ pdits = 0
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ noff = 2.2684
+ cigsd = 0.013281
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ aigbinv = 0.009974
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ pags = -1.92428e-14
+ ntox = -1.9260000000000002
+ pcit = 0
+ rgatemod = 0
+ pclm = 1.101657
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ ptvfbsdoff = 0
+ tnjtsswg = 1
+ phin = 0.15
+ tnoia = 0
+ pkt1 = -2.8122214e-15
+ pkt2 = 2.4239149e-16
+ peta0 = -1.5e-17
+ toxref = 3e-9
+ wketa = -2.0595747e-9
+ poxedge = 1
+ tpbsw = 0.0025
+ cjswd = 5.457e-11
+ cjsws = 5.457e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ rbdb = 50
+ pua1 = -1.1776704e-22
+ binunit = 2
+ prwb = 0
+ pub1 = 2.7996299e-31
+ prwg = 0
+ puc1 = 9.811687e-24
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ pute = 1.5923616e-14
+ rdsw = 200
+ tvfbsdoff = 0.1
+ ltvoff = -3.3500511e-10
+ scref = 1e-6
+ pigcd = 2.572
+ rshg = 14.1
+ aigsd = 0.0063632604
+ lku0we = 1.8e-11
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ epsrox = 3.9
+ lvoff = -2.4480721e-8
+ a0 = 2.6314952
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ rdsmod = 0
+ wvfbsdoff = 0
+ at = 72000
+ cf = 7.598099999999999e-11
+ lvsat = 0.00024
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.016004612
+ k3 = -2.5823
+ em = 20000000.0
+ lvfbsdoff = 0
+ lvth0 = -1.4466904e-8
+ igbmod = 1
+ ll = 0
+ lw = 0
+ u0 = 0.009736307500000001
+ w0 = 0
+ ua = -1.8414289e-10
+ ub = 1.2263153e-18
+ uc = -3.3458683e-12
+ ud = 0
+ ijthsfwd = 0.01
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 5.6700000000000005e-9
+ ww = 0
+ xw = 3.4e-9
+ delta = 0.018814
+ laigc = -5.3027874e-11
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ rnoia = 0
+ rnoib = 0
+ pbswgd = 0.8
+ pbswgs = 0.8
+ tnom = 25
+ toxe = 2.71e-9
+ toxm = 2.67e-9
+ igcmod = 1
+ pketa = 1.0887638e-15
+ ngate = 1.7e+20
+ ngcon = 1
+ ijthsrev = 0.01
+ wpclm = 7.1298978e-9
+ njtsswg = 6.489
+ gbmin = 1e-12
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ wags = 7.3346686e-9
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.00084883969
+ pdiblcb = 0
+ paigsd = -1.2880862e-20
+ voff = -0.10099712
+ acde = 0.5
+ ppdiblc2 = -2.0561872e-16
+ vsat = 108525.44
+ wint = 0
+ permod = 1
+ vth0 = -0.39832868000000005
+ wkt1 = -2.7375492e-9
+ wkt2 = -7.5529568e-10
+ wmax = 2.726e-7
+ aigc = 0.0068361189
+ wmin = 1.08e-7
+ bigbacc = 0.0054401
+ tvoff = 0.0025796189
+ kvth0we = -0.00022
+ wua1 = -4.222676e-17
+ wub1 = -1.3803658e-25
+ wuc1 = -1.3210867e-17
+ xjbvd = 1
+ xjbvs = 1
+ voffcv = -0.125
+ wpemod = 1
+ lk2we = 0.0
+ lintnoi = -5e-9
+ bigc = 0.0012521
+ wute = -7.8294814e-8
+ bigbinv = 0.00149
+ pkvth0we = 0.0
+ wwlc = 0
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ cdsc = 0
+ ku0we = -0.0007
+ cgbo = 0
+ cgdl = 2.799765e-11
+ cgdo = 2.4628259999999997e-11
+ xtid = 3
+ xtis = 3
+ beta0 = 13.32
+ leta0 = -5e-10
+ vfbsdoff = 0.01
+ cgsl = 2.799765e-11
+ cgso = 2.4628259999999997e-11
+ cigc = 0.15259
+ ppclm = 0
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ paramchk = 1
+ tpbswg = 0.001
+ )

.model pch_ss_35 pmos (
+ level = 54
+ cjsws = 5.457e-11
+ cjswgd = 1.9367000000000001e-10
+ pku0we = 0.0
+ cjswgs = 1.9367000000000001e-10
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ ndep = 1e+18
+ lute = -1.0958354e-8
+ lwlc = 0
+ moin = 5.5538
+ ijthsrev = 0.01
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ tvfbsdoff = 0.1
+ nigc = 2.291
+ mjswgd = 0.95
+ mjswgs = 0.95
+ tcjswg = 0.00128
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ scref = 1e-6
+ pags = 1.1742809e-13
+ ppdiblc2 = -6.1367245e-16
+ pigcd = 2.572
+ ntox = -1.9260000000000002
+ aigsd = 0.0063632396
+ pcit = 0
+ pclm = 1.101657
+ lvoff = -2.4340257e-9
+ phin = 0.15
+ wvfbsdoff = 0
+ njtsswg = 6.489
+ lvfbsdoff = 0
+ lvsat = 0.00024
+ lvth0 = -6.2799405e-10
+ pkt1 = 5.7473332e-15
+ pkt2 = -5.7270183e-16
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ delta = 0.018814
+ fprout = 200
+ laigc = -3.3884553e-11
+ xrcrg1 = 12
+ xrcrg2 = 1
+ ckappad = 0.6
+ ckappas = 0.6
+ rnoia = 0
+ rnoib = 0
+ pdiblc1 = 0
+ pdiblc2 = 0.0027845581
+ pdiblcb = 0
+ pkvth0we = 0.0
+ rbdb = 50
+ pua1 = -9.8048843e-24
+ prwb = 0
+ pub1 = -2.3189739e-32
+ prwg = 0
+ puc1 = -4.5795492e-24
+ pketa = -3.0075994e-15
+ rbpb = 50
+ rbpd = 50
+ ngate = 1.7e+20
+ rbps = 50
+ rbsb = 50
+ wtvoff = -2.2790108e-10
+ pvag = 2.1
+ pute = -9.4649237e-15
+ ngcon = 1
+ wpclm = 7.1298978e-9
+ rdsw = 200
+ vfbsdoff = 0.01
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ bigbacc = 0.0054401
+ capmod = 2
+ wku0we = 1.5e-11
+ kvth0we = -0.00022
+ mobmod = 0
+ paramchk = 1
+ lintnoi = -5e-9
+ rshg = 14.1
+ bigbinv = 0.00149
+ wtvfbsdoff = 0
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ ltvfbsdoff = 0
+ ijthdfwd = 0.01
+ tvoff = 0.0027416725
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ tnom = 25
+ toxe = 2.71e-9
+ toxm = 2.67e-9
+ ijthdrev = 0.01
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = -5e-10
+ lpdiblc2 = 4.574275e-9
+ ptvfbsdoff = 0
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ nfactor = 1
+ ppclm = 0
+ wags = -1.4622812e-7
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ voff = -0.12576869
+ acde = 0.5
+ vsat = 108525.44
+ wint = 0
+ vth0 = -0.41387802
+ wkt1 = -1.2355026e-8
+ wkt2 = 1.605395e-10
+ dmcgt = 0
+ wmax = 2.726e-7
+ tcjsw = 9.34e-5
+ lkvth0we = 3e-12
+ aigc = 0.0068146096
+ wmin = 1.08e-7
+ nigbacc = 10
+ toxref = 3e-9
+ wua1 = -1.6353255e-16
+ wub1 = 2.0258446e-25
+ wuc1 = 2.9590615e-18
+ acnqsmod = 0
+ bigsd = 0.0003327
+ bigc = 0.0012521
+ wute = -4.9768365e-8
+ nigbinv = 2.171
+ wwlc = 0
+ wvoff = 3.4766421e-9
+ rbodymod = 0
+ cdsc = 0
+ cgbo = 0
+ cgdl = 2.799765e-11
+ cgdo = 2.4628259999999997e-11
+ wvsat = -0.0013318206
+ xtid = 3
+ xtis = 3
+ wvth0 = -5.3516532e-9
+ ltvoff = -4.7923289e-10
+ cgsl = 2.799765e-11
+ cgso = 2.4628259999999997e-11
+ cigc = 0.15259
+ waigc = 2.7104678e-12
+ fnoimod = 1
+ eigbinv = 1.1
+ pvfbsdoff = 0
+ lketa = 4.197898e-9
+ xpart = 1
+ lku0we = 1.8e-11
+ epsrox = 3.9
+ wpdiblc2 = 8.1773971e-10
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ ags = 1.7348065
+ dmdg = 0
+ egidl = 0.001
+ cjd = 0.00144022
+ rdsmod = 0
+ cit = -8.7888889e-5
+ cjs = 0.00144022
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 1.0572421799999999e-8
+ igbmod = 1
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ k2we = 5e-5
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ dsub = 0.5
+ dtox = 3.91e-10
+ pbswgd = 0.8
+ la0 = -1.044589e-6
+ cigbacc = 0.245
+ pbswgs = 0.8
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0.001
+ kt1 = -0.11040563
+ kt2 = -0.048714998
+ lk2 = 3.4890726e-9
+ llc = 0
+ lln = 1
+ lu0 = -1.8122817999999998e-9
+ mjd = 0.335
+ mjs = 0.335
+ lua = -6.2776752e-16
+ lub = 4.4518935e-25
+ luc = 5.1177769e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ igcmod = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 1.0817056e-13
+ wkvth0we = 0.0
+ nsd = 1e+20
+ pbd = 0.75
+ tnoimod = 0
+ pat = 0
+ pbs = 0.75
+ pk2 = -1.5480351e-16
+ eta0 = 0.10792519
+ etab = -0.13555556
+ pu0 = 1.5955157e-16
+ prt = 0
+ pua = 4.4574845e-23
+ pub = -2.7161351e-32
+ puc = -4.8372521e-24
+ pud = 0
+ rsh = 15.2
+ trnqsmod = 0
+ tcj = 0.000832
+ ua1 = 2.771768e-9
+ ub1 = -3.1924567e-18
+ uc1 = -6.2120134e-12
+ cigbinv = 0.006
+ tpb = 0.0016
+ wa0 = -1.0464262e-7
+ ute = -0.78783539
+ pvoff = -9.6675093e-16
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 4.174453e-9
+ wlc = 0
+ wln = 1
+ wu0 = -8.9929205e-11
+ xgl = -8.2e-9
+ xgw = 0
+ wua = -7.0620672e-17
+ wub = -4.621089e-27
+ wuc = 8.8883858e-18
+ wud = 0
+ cdscb = 0
+ cdscd = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ pvsat = -5e-11
+ a0 = 3.3624733
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ wk2we = 0.0
+ pvth0 = 1.0530712e-16
+ at = 72000
+ cf = 7.598099999999999e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.013259817
+ k3 = -2.5823
+ em = 20000000.0
+ drout = 0.56
+ version = 4.5
+ ll = 0
+ lw = 0
+ u0 = 0.012898186
+ w0 = 0
+ ua = 4.4026063e-10
+ ub = 1.2150282e-18
+ uc = -4.4814963e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 5.6700000000000005e-9
+ ww = 0
+ paigc = 4.1038726e-19
+ xw = 3.4e-9
+ tempmod = 0
+ voffl = 0
+ rgatemod = 0
+ permod = 1
+ tnjtsswg = 1
+ weta0 = 1.9403288999999997e-9
+ wetab = 2.9133333e-9
+ aigbacc = 0.012071
+ lpclm = 0
+ cgidl = 1
+ voffcv = -0.125
+ wpemod = 1
+ aigbinv = 0.009974
+ pbswd = 0.9
+ pbsws = 0.9
+ keta = -0.035939983
+ pdits = 0
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ lags = -3.1625612e-7
+ tpbswg = 0.001
+ poxedge = 1
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 8.2671111e-11
+ kt1l = 0
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ binunit = 2
+ lint = 6.5375218e-9
+ ptvoff = 8.8703803e-17
+ lkt1 = -6.3138035e-8
+ lkt2 = -3.1463267e-9
+ tnoia = 0
+ lmax = 8.974099999999999e-7
+ waigsd = 1.9716411e-12
+ lmin = 4.4741e-7
+ ijthsfwd = 0.01
+ peta0 = -1.5e-17
+ lpe0 = 6.44e-8
+ lpeb = 0
+ wketa = 2.5430806e-9
+ diomod = 1
+ tpbsw = 0.0025
+ minv = -0.33
+ lua1 = -1.8157361e-16
+ lub1 = 3.2089876e-25
+ luc1 = 1.2550631e-17
+ pditsd = 0
+ cjswd = 5.457e-11
+ pditsl = 0
+ )

.model pch_ss_36 pmos (
+ level = 54
+ ags = 0.79842724
+ pvfbsdoff = 0
+ wcit = 5.8162887e-11
+ lketa = -1.0850486e-8
+ cigbacc = 0.245
+ cjd = 0.00144022
+ cit = -0.00049977211
+ cjs = 0.00144022
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ voff = -0.11894985
+ xpart = 1
+ dlc = 1.38228675e-8
+ k3b = 2.1176
+ acde = 0.5
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ rgatemod = 0
+ tnjtsswg = 1
+ vsat = 108525.44
+ tnoimod = 0
+ wint = 0
+ vth0 = -0.42050626
+ egidl = 0.001
+ wkt1 = 8.365112e-10
+ wkt2 = -1.4765978e-9
+ la0 = -3.2362015e-7
+ wmax = 2.726e-7
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0.001
+ aigc = 0.0068096243
+ wmin = 1.08e-7
+ kt1 = -0.25321364
+ kt2 = -0.04359324
+ lk2 = 5.726910000000002e-11
+ llc = -1.18e-13
+ lln = 0.7
+ cigbinv = 0.006
+ lu0 = -4.4559608e-10
+ mjd = 0.335
+ mjs = 0.335
+ lua = -1.7021816e-16
+ lub = 1.0550853e-25
+ luc = -1.2975077e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ fprout = 200
+ njs = 1.02
+ pa0 = -3.1370244e-14
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ pk2 = 1.4083403e-16
+ xrcrg1 = 12
+ xrcrg2 = 1
+ pu0 = -1.3937081e-17
+ prt = 0
+ pua = 4.7117679e-24
+ pub = -8.7289665e-33
+ puc = -3.0945045e-25
+ pud = 0
+ wua1 = -2.3000717e-16
+ wub1 = 1.2114667e-25
+ wuc1 = -1.9684753e-17
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 2.6350858e-9
+ ub1 = -2.2549964e-18
+ uc1 = 3.1191962e-11
+ bigc = 0.0012521
+ wute = -1.1762912e-7
+ version = 4.5
+ tpb = 0.0016
+ wa0 = 2.1249557e-7
+ wwlc = 0
+ ute = -0.71022675
+ wtvoff = -1.1036076e-10
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 3.5025496e-9
+ tempmod = 0
+ wlc = 0
+ wln = 1
+ wu0 = 3.0436319e-10
+ xgl = -8.2e-9
+ xgw = 0
+ wua = 1.9977231e-17
+ wub = -4.6512873e-26
+ wuc = -1.4020724e-18
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ cdsc = 0
+ cgbo = 0
+ cgdl = 2.799765e-11
+ cgdo = 2.4628259999999997e-11
+ xtid = 3
+ xtis = 3
+ wtvfbsdoff = 0
+ aigbacc = 0.012071
+ cgsl = 2.799765e-11
+ cgso = 2.4628259999999997e-11
+ cigc = 0.15259
+ pvoff = 1.20942711e-16
+ capmod = 2
+ cdscb = 0
+ cdscd = 0
+ wku0we = 1.5e-11
+ pvsat = -5e-11
+ wk2we = 0.0
+ pvth0 = -3.0393785e-16
+ ltvfbsdoff = 0
+ drout = 0.56
+ mobmod = 0
+ paigc = -1.759214e-19
+ aigbinv = 0.009974
+ voffl = 0
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ weta0 = 1.9403288999999997e-9
+ wetab = 2.9133333e-9
+ lpclm = 0
+ k2we = 5e-5
+ ijthsfwd = 0.01
+ cgidl = 1
+ dsub = 0.5
+ ptvfbsdoff = 0
+ dtox = 3.91e-10
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ poxedge = 1
+ eta0 = 0.10792519
+ pbswd = 0.9
+ etab = -0.13555556
+ pbsws = 0.9
+ ijthsrev = 0.01
+ binunit = 2
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ pdits = 0
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ ppdiblc2 = 9.2177422e-17
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ tnoia = 0
+ toxref = 3e-9
+ peta0 = -1.5e-17
+ wketa = -1.9938172e-9
+ tpbsw = 0.0025
+ cjswd = 5.457e-11
+ cjsws = 5.457e-11
+ pkvth0we = 0.0
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ tvfbsdoff = 0.1
+ ltvoff = -1.9203223e-10
+ vfbsdoff = 0.01
+ njtsswg = 6.489
+ keta = -0.0017391106
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ lags = 9.5750741e-8
+ lku0we = 1.8e-11
+ paramchk = 1
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ scref = 1e-6
+ ckappad = 0.6
+ ckappas = 0.6
+ lcit = 2.6389973e-10
+ pdiblc1 = 0
+ pdiblc2 = 0.016049816
+ epsrox = 3.9
+ pdiblcb = 0
+ pigcd = 2.572
+ kt1l = 0
+ aigsd = 0.0063632396
+ rdsmod = 0
+ lvoff = -5.4343156e-9
+ wvfbsdoff = 0
+ lint = 9.7879675e-9
+ igbmod = 1
+ lvfbsdoff = 0
+ lkt1 = -3.021340000000001e-10
+ lkt2 = -5.3999005e-9
+ lvsat = 0.00024
+ lmax = 4.4741e-7
+ lvth0 = 2.2884329e-9
+ lmin = 2.1410000000000002e-7
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ ijthdfwd = 0.01
+ lpe0 = 6.44e-8
+ delta = 0.018814
+ bigbacc = 0.0054401
+ lpeb = 0
+ pbswgd = 0.8
+ laigc = -3.1691048e-11
+ pbswgs = 0.8
+ rnoia = 0
+ rnoib = 0
+ minv = -0.33
+ igcmod = 1
+ lua1 = -1.2143343e-16
+ lub1 = -9.158653e-26
+ luc1 = -3.907118e-18
+ kvth0we = -0.00022
+ ndep = 1e+18
+ lute = -4.5106156e-8
+ pketa = -1.0113644e-15
+ ngate = 1.7e+20
+ lwlc = 0
+ lintnoi = -5e-9
+ moin = 5.5538
+ ijthdrev = 0.01
+ ngcon = 1
+ bigbinv = 0.00149
+ wpclm = 7.1298978e-9
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ nigc = 2.291
+ lpdiblc2 = -1.262443e-9
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ pags = 5.2660461e-14
+ permod = 1
+ ntox = -1.9260000000000002
+ pcit = -2.559167e-17
+ pclm = 1.101657
+ phin = 0.15
+ lkvth0we = 3e-12
+ pkt1 = -5.70475e-17
+ pkt2 = 1.4763857e-16
+ voffcv = -0.125
+ wpemod = 1
+ tvoff = 0.0020889601
+ nfactor = 1
+ xjbvd = 1
+ acnqsmod = 0
+ xjbvs = 1
+ lk2we = 0.0
+ a0 = 1.7239078
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ rbdb = 50
+ pua1 = 1.9443948e-23
+ prwb = 0
+ pub1 = 1.2643651e-32
+ prwg = 0
+ at = 72000
+ puc1 = 5.3837292e-24
+ cf = 7.598099999999999e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.0054602636
+ k3 = -2.5823
+ em = 20000000.0
+ rbpb = 50
+ rbpd = 50
+ ll = -1.18e-13
+ lw = 0
+ rbps = 50
+ u0 = 0.009792082
+ rbsb = 50
+ pvag = 2.1
+ w0 = 0
+ rbodymod = 0
+ ua = -5.9962427e-10
+ ub = 1.98703e-18
+ uc = 1.0098696e-10
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 5.6700000000000005e-9
+ ww = 0
+ pute = 2.0393808e-14
+ xw = 3.4e-9
+ rdsw = 200
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = -5e-10
+ nigbacc = 10
+ ppclm = 0
+ tpbswg = 0.001
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ rshg = 14.1
+ nigbinv = 2.171
+ wpdiblc2 = -7.8646151e-10
+ ptvoff = 3.6984079e-17
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ waigsd = 1.9716411e-12
+ diomod = 1
+ fnoimod = 1
+ pditsd = 0
+ pditsl = 0
+ bigsd = 0.0003327
+ cjswgd = 1.9367000000000001e-10
+ pku0we = 0.0
+ tnom = 25
+ cjswgs = 1.9367000000000001e-10
+ eigbinv = 1.1
+ toxe = 2.71e-9
+ toxm = 2.67e-9
+ wkvth0we = 0.0
+ wvoff = 1.0046111e-9
+ trnqsmod = 0
+ wvsat = -0.0013318206
+ mjswgd = 0.95
+ wvth0 = -4.421551e-9
+ mjswgs = 0.95
+ tcjswg = 0.00128
+ waigc = 4.0429874e-12
+ wags = 9.7102189e-10
+ )

.model pch_ss_37 pmos (
+ level = 54
+ fprout = 200
+ lvth0 = 4.927490499999999e-9
+ xrcrg1 = 12
+ xrcrg2 = 1
+ delta = 0.018814
+ wtvfbsdoff = 0
+ laigc = -4.357169e-12
+ rnoia = 0
+ rnoib = 0
+ acnqsmod = 0
+ wtvoff = 1.2048366e-10
+ ltvfbsdoff = 0
+ pketa = 4.1278959e-16
+ ngate = 1.7e+20
+ rbodymod = 0
+ ngcon = 1
+ wpclm = 6.8691006e-8
+ capmod = 2
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ wku0we = 1.5e-11
+ keta = -0.058692164
+ mobmod = 0
+ nfactor = 1
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 2.5291477e-11
+ ptvfbsdoff = 0
+ kt1l = 0
+ wpdiblc2 = -7.28246e-10
+ lint = 9.7879675e-9
+ lkt1 = -5.6770694e-9
+ lkt2 = -3.7791597e-9
+ lmax = 2.1410000000000002e-7
+ lmin = 8.833e-8
+ lpe0 = 6.44e-8
+ nigbacc = 10
+ lpeb = 0
+ tvoff = 0.0011827459
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ minv = -0.33
+ lua1 = -2.1218464e-16
+ lub1 = 2.7818737e-25
+ luc1 = 2.2554944e-17
+ ndep = 1e+18
+ wkvth0we = 0.0
+ lute = 1.5508066e-9
+ lwlc = 0
+ moin = 5.5538
+ nigbinv = 2.171
+ ku0we = -0.0007
+ trnqsmod = 0
+ beta0 = 13.32
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ nigc = 2.291
+ leta0 = -5e-10
+ ppclm = -1.2989269e-14
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ fnoimod = 1
+ eigbinv = 1.1
+ ntox = -1.9260000000000002
+ rgatemod = 0
+ pcit = 1.1214196e-17
+ pclm = 0.85425247
+ tnjtsswg = 1
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ phin = 0.15
+ toxref = 3e-9
+ pkt1 = -2.317336e-16
+ pkt2 = 3.7767926e-16
+ bigsd = 0.0003327
+ cigbacc = 0.245
+ rbdb = 50
+ pua1 = 2.6827919e-23
+ prwb = 0
+ pub1 = -3.4278711e-32
+ prwg = 0
+ puc1 = -2.7535024e-24
+ wvoff = 8.5374562e-10
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ pute = -4.2802262e-16
+ ltvoff = -8.1627e-13
+ rdsw = 200
+ tnoimod = 0
+ wvsat = -0.00089129698
+ ags = 1.2522222
+ wvth0 = -5.450948e-9
+ cjd = 0.00144022
+ cit = 0.00063107268
+ cjs = 0.00144022
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 1.38228675e-8
+ waigc = 1.4660694e-11
+ k3b = 2.1176
+ cigbinv = 0.006
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ pvfbsdoff = 0
+ lku0we = 1.8e-11
+ lketa = 1.1666086e-9
+ epsrox = 3.9
+ la0 = 6.219346e-9
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = -0.0065443287
+ xpart = 1
+ kt1 = -0.22773883
+ kt2 = -0.051274476
+ lk2 = 4.0711471e-9
+ llc = -1.18e-13
+ lln = 0.7
+ lu0 = -1.5814862e-10
+ mjd = 0.335
+ version = 4.5
+ mjs = 0.335
+ lua = 1.3101868e-17
+ lub = -8.7271368e-26
+ luc = -1.2812174e-17
+ lud = 0
+ rshg = 14.1
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = -2.0637395e-14
+ rdsmod = 0
+ nsd = 1e+20
+ pbd = 0.75
+ tempmod = 0
+ pat = -5.0045721e-10
+ pbs = 0.75
+ pk2 = 4.0368065e-17
+ egidl = 0.001
+ igbmod = 1
+ pu0 = -5.2679707e-18
+ prt = 0
+ pua = -4.0286539e-24
+ pub = 7.5106005e-33
+ puc = 1.4358513e-24
+ pud = 0
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 3.0651863e-9
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ ub1 = -4.0074881e-18
+ uc1 = -9.4220652e-11
+ tpb = 0.0016
+ aigbacc = 0.012071
+ wa0 = 1.6162969e-7
+ pbswgd = 0.8
+ pbswgs = 0.8
+ ute = -0.93134979
+ ijthsfwd = 0.01
+ wat = 0.0023718351
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 3.9786916e-9
+ wlc = 0
+ wln = 1
+ wu0 = 2.6327735e-10
+ xgl = -8.2e-9
+ xgw = 0
+ wua = 6.1401032e-17
+ wub = -1.2347765e-25
+ wuc = -9.6736445e-18
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ igcmod = 1
+ tnom = 25
+ toxe = 2.71e-9
+ toxm = 2.67e-9
+ aigbinv = 0.009974
+ ijthsrev = 0.01
+ pvoff = 1.5277532e-16
+ cdscb = 0
+ cdscd = 0
+ pvsat = -1.42948987e-10
+ wags = 2.5054667e-7
+ wk2we = 0.0
+ pvth0 = -8.6735092e-17
+ drout = 0.56
+ wcit = -1.162725e-10
+ paigc = -2.4162575e-18
+ permod = 1
+ voff = -0.1339517
+ acde = 0.5
+ ppdiblc2 = 7.9894307e-17
+ voffl = 0
+ poxedge = 1
+ vsat = 106518.57
+ wint = 0
+ vth0 = -0.43301365
+ weta0 = 1.9403288999999997e-9
+ wetab = 2.9133333e-9
+ wkt1 = 1.664079e-9
+ wkt2 = -2.566838e-9
+ wmax = 2.726e-7
+ lpclm = 5.2201277e-8
+ binunit = 2
+ aigc = 0.0066800799
+ wmin = 1.08e-7
+ voffcv = -0.125
+ wpemod = 1
+ cgidl = 1
+ wua1 = -2.6500229e-16
+ wub1 = 3.4352994e-25
+ wuc1 = 1.8880326e-17
+ bigc = 0.0012521
+ wute = -1.8947457e-8
+ pkvth0we = 0.0
+ wwlc = 0
+ pbswd = 0.9
+ pbsws = 0.9
+ cdsc = 0
+ cgbo = 0
+ cgdl = 2.799765e-11
+ cgdo = 2.4628259999999997e-11
+ xtid = 3
+ xtis = 3
+ vfbsdoff = 0.01
+ cgsl = 2.799765e-11
+ cgso = 2.4628259999999997e-11
+ cigc = 0.15259
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ pdits = 0
+ tpbswg = 0.001
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ paramchk = 1
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ ptvoff = -1.1725409e-17
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ a0 = 0.16068118
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ waigsd = 1.9716411e-12
+ at = 107755.11
+ cf = 7.598099999999999e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.024483382
+ k3 = -2.5823
+ em = 20000000.0
+ ll = -1.18e-13
+ lw = 0
+ u0 = 0.008429771800000001
+ tnoia = 0
+ w0 = 0
+ ua = -1.4684396e-9
+ ub = 2.9006788e-18
+ uc = 1.0021491e-10
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 5.6700000000000005e-9
+ ww = 0
+ xw = 3.4e-9
+ diomod = 1
+ k2we = 5e-5
+ ijthdfwd = 0.01
+ peta0 = -1.5e-17
+ njtsswg = 6.489
+ dsub = 0.5
+ dtox = 3.91e-10
+ wketa = -8.743362e-9
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.9367000000000001e-10
+ pku0we = 0.0
+ cjswgs = 1.9367000000000001e-10
+ tpbsw = 0.0025
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ cjswd = 5.457e-11
+ cjsws = 5.457e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.01690182
+ eta0 = 0.10792519
+ pdiblcb = 0
+ etab = -0.13555556
+ tvfbsdoff = 0.1
+ ijthdrev = 0.01
+ mjswgd = 0.95
+ mjswgs = 0.95
+ lpdiblc2 = -1.4422174e-9
+ tcjswg = 0.00128
+ bigbacc = 0.0054401
+ scref = 1e-6
+ pigcd = 2.572
+ aigsd = 0.0063632396
+ kvth0we = -0.00022
+ wvfbsdoff = 0
+ lvoff = -2.268926e-9
+ lintnoi = -5e-9
+ lvfbsdoff = 0
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ lkvth0we = 3e-12
+ lvsat = 0.00066343719
+ )

.model pch_ss_38 pmos (
+ level = 54
+ poxedge = 1
+ ptvfbsdoff = 0
+ rdsw = 200
+ capmod = 2
+ vfbsdoff = 0.01
+ wku0we = 1.5e-11
+ pvoff = -1.1873467e-16
+ binunit = 2
+ cdscb = 0
+ cdscd = 0
+ mobmod = 0
+ pvsat = 1.2296039999999998e-10
+ wk2we = 0.0
+ pvth0 = 2.8090213400000003e-16
+ drout = 0.56
+ paramchk = 1
+ paigc = -1.1563004e-18
+ voffl = 0
+ rshg = 14.1
+ weta0 = 1.2757501e-8
+ wetab = 4.1458967e-9
+ lpclm = -1.0127779e-7
+ ijthdfwd = 0.01
+ jtsswgd = 1.75e-7
+ cgidl = 1
+ jtsswgs = 1.75e-7
+ tnom = 25
+ toxe = 2.71e-9
+ toxm = 2.67e-9
+ pbswd = 0.9
+ pbsws = 0.9
+ ijthdrev = 0.01
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ lpdiblc2 = -1.4113545e-11
+ pdits = 0
+ cigsd = 0.013281
+ wags = 2.5054667e-7
+ dvt0w = 0
+ dvt1w = 0
+ njtsswg = 6.489
+ dvt2w = 0
+ wcit = -1.17261256e-10
+ xtsswgd = 0.32
+ voff = -0.14478455
+ xtsswgs = 0.32
+ acde = 0.5
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ ckappad = 0.6
+ ckappas = 0.6
+ vsat = 137363.5
+ wint = 0
+ pdiblc1 = 0
+ pdiblc2 = 0.0017092259
+ vth0 = -0.35846913
+ pdiblcb = 0
+ wkt1 = -1.350742e-8
+ wkt2 = 1.8825744e-9
+ toxref = 3e-9
+ wmax = 2.726e-7
+ lkvth0we = 3e-12
+ aigc = 0.0067219883
+ wmin = 1.08e-7
+ tnoia = 0
+ peta0 = -1.0318142000000001e-15
+ petab = -1.1586096e-16
+ wketa = -6.6698086e-9
+ wua1 = 1.6631395e-16
+ wub1 = -2.121384e-25
+ wuc1 = 2.5860689e-17
+ tpbsw = 0.0025
+ acnqsmod = 0
+ bigbacc = 0.0054401
+ cjswd = 5.457e-11
+ bigc = 0.0012521
+ cjsws = 5.457e-11
+ wute = -6.1363432e-8
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ wwlc = 0
+ tvfbsdoff = 0.1
+ ltvoff = 3.7319947e-11
+ rbodymod = 0
+ kvth0we = -0.00022
+ cdsc = 0
+ cgbo = 0
+ cgdl = 2.799765e-11
+ cgdo = 2.4628259999999997e-11
+ xtid = 3
+ xtis = 3
+ lintnoi = -5e-9
+ cgsl = 2.799765e-11
+ cgso = 2.4628259999999997e-11
+ bigbinv = 0.00149
+ cigc = 0.15259
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ lku0we = 1.8e-11
+ epsrox = 3.9
+ scref = 1e-6
+ pigcd = 2.572
+ aigsd = 0.0063632396
+ rdsmod = 0
+ wpdiblc2 = 8.0253658e-11
+ igbmod = 1
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ lvoff = -1.2506377e-9
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ lvsat = -0.0022359865
+ pbswgd = 0.8
+ pbswgs = 0.8
+ lvth0 = -2.0796987e-9
+ k2we = 5e-5
+ delta = 0.018814
+ laigc = -8.2965642e-12
+ dsub = 0.5
+ igcmod = 1
+ dtox = 3.91e-10
+ rnoia = 0
+ rnoib = 0
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ nfactor = 1
+ wkvth0we = 0.0
+ pketa = 2.1787556e-16
+ ngate = 1.7e+20
+ eta0 = 0.024468866
+ etab = -0.22797789
+ ngcon = 1
+ wpclm = -1.6917696e-7
+ trnqsmod = 0
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ nigbacc = 10
+ permod = 1
+ rgatemod = 0
+ tnjtsswg = 1
+ nigbinv = 2.171
+ voffcv = -0.125
+ wpemod = 1
+ tvoff = 0.00077704148
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ fnoimod = 1
+ eigbinv = 1.1
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = 7.344893999999999e-9
+ letab = 8.6876992e-9
+ tpbswg = 0.001
+ ppclm = 9.3703198e-15
+ keta = -0.049241031
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 1.2394067e-10
+ kt1l = 0
+ ptvoff = 1.952106e-17
+ cigbacc = 0.245
+ waigsd = 1.9716411e-12
+ dmcgt = 0
+ lint = 0
+ tcjsw = 9.34e-5
+ tnoimod = 0
+ lkt1 = -7.5946074e-9
+ lkt2 = 9.2375447e-10
+ diomod = 1
+ lmax = 8.833e-8
+ lmin = 5.233e-8
+ ijthsfwd = 0.01
+ lpe0 = 6.44e-8
+ pditsd = 0
+ pditsl = 0
+ lpeb = 0
+ cigbinv = 0.006
+ cjswgd = 1.9367000000000001e-10
+ pku0we = 0.0
+ cjswgs = 1.9367000000000001e-10
+ bigsd = 0.0003327
+ minv = -0.33
+ ags = 1.2522222
+ lua1 = 1.5814311e-16
+ lub1 = -2.3663254e-25
+ luc1 = 3.1466117e-17
+ cjd = 0.00144022
+ cit = -0.00041837991
+ cjs = 0.00144022
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ ndep = 1e+18
+ bvs = 8.2
+ lute = -1.2895214e-8
+ dlc = 4.0349e-9
+ wvoff = 3.7421498e-9
+ k3b = 2.1176
+ lwlc = 0
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ version = 4.5
+ moin = 5.5538
+ mjswgd = 0.95
+ mjswgs = 0.95
+ ijthsrev = 0.01
+ tempmod = 0
+ wvsat = -0.0037201203
+ nigc = 2.291
+ tcjswg = 0.00128
+ wvth0 = -9.361984e-9
+ la0 = 3.4503642e-8
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = -0.0070528058999999995
+ kt1 = -0.20733948
+ kt2 = -0.10130548
+ lk2 = 5.947863e-9
+ waigc = 1.256895e-12
+ llc = 0
+ lln = 1
+ a0 = -0.1402156
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ lu0 = 5.0809140000000005e-11
+ mjd = 0.335
+ mjs = 0.335
+ lua = 1.1003971e-16
+ lub = -1.3258131e-25
+ luc = -1.072064e-17
+ at = 113164.44
+ lud = 0
+ cf = 7.598099999999999e-11
+ lwc = 0
+ pvfbsdoff = 0
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.044448444
+ k3 = -2.5823
+ lwl = 0
+ lwn = 1
+ em = 20000000.0
+ aigbacc = 0.012071
+ njd = 1.02
+ njs = 1.02
+ ll = 0
+ noff = 2.2684
+ pa0 = -6.959911e-15
+ lw = 0
+ u0 = 0.0062068169
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ w0 = 0
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 1.1859675e-9
+ ua = -2.4996932e-9
+ ub = 3.3826995e-18
+ uc = 7.7964547e-11
+ ud = 0
+ pbs = 0.75
+ pk2 = -8.547569e-17
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 5.6700000000000005e-9
+ ww = 0
+ xw = 3.4e-9
+ pu0 = 1.7354187e-18
+ prt = 0
+ lketa = 2.7820203e-10
+ pua = -5.4706466e-24
+ pub = 7.2761107e-33
+ puc = 2.7207836e-25
+ pud = 0
+ wtvfbsdoff = 0
+ xpart = 1
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = -8.7447052e-10
+ ub1 = 1.4693195e-18
+ uc1 = -1.8902037e-10
+ ppdiblc2 = 3.8953385e-18
+ ntox = -1.9260000000000002
+ tpb = 0.0016
+ pcit = 1.1307033299999999e-17
+ pclm = 2.4870084
+ wa0 = 1.612455e-8
+ ute = -0.77766872
+ wat = -0.015568853
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 5.3174549e-9
+ aigbinv = 0.009974
+ wlc = 0
+ egidl = 0.001
+ wln = 1
+ wu0 = 1.8877321e-10
+ xgl = -8.2e-9
+ xgw = 0
+ wua = 7.6741379e-17
+ wub = -1.2098307e-25
+ wuc = 2.7069183e-18
+ wud = 0
+ wwc = 0
+ ltvfbsdoff = 0
+ wwl = 0
+ wwn = 1
+ phin = 0.15
+ fprout = 200
+ xrcrg1 = 12
+ xrcrg2 = 1
+ pkt1 = 1.1943873e-15
+ pkt2 = -4.056551e-17
+ wtvoff = -2.1192558e-10
+ pkvth0we = 0.0
+ rbdb = 50
+ pua1 = -1.3715808e-23
+ prwb = 0
+ pub1 = 1.7954113e-32
+ prwg = 0
+ puc1 = -3.4096566e-24
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ pute = 3.5590791e-15
+ )

.model pch_ss_39 pmos (
+ level = 54
+ fnoimod = 1
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ eigbinv = 1.1
+ k2we = 5e-5
+ ijthsfwd = 0.01
+ tvoff = 0.00092289205
+ dsub = 0.5
+ dtox = 3.91e-10
+ xjbvd = 1
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ xjbvs = 1
+ lk2we = 0.0
+ eta0 = 0.19463541
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ etab = -0.16706384
+ ijthsrev = 0.01
+ cigbacc = 0.245
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = -2.5247657e-9
+ letab = 5.1546845e-9
+ tnoimod = 0
+ ppclm = 7.8094068e-15
+ dlcig = 2.5e-9
+ cigbinv = 0.006
+ bgidl = 1834800000.0
+ ppdiblc2 = 0
+ toxref = 3e-9
+ version = 4.5
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ tempmod = 0
+ ags = 1.2522222
+ cjd = 0.00144022
+ cit = -0.0001366287
+ cjs = 0.00144022
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 4.0349e-9
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ aigbacc = 0.012071
+ bigsd = 0.0003327
+ pkvth0we = 0.0
+ la0 = -1.4904033e-7
+ ltvoff = 2.8860613e-11
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0.010372508999999999
+ kt1 = -0.53950997
+ kt2 = -0.12590838
+ lk2 = 4.6165993000000006e-9
+ wvoff = 1.4341134e-10
+ llc = 0
+ lln = 1
+ lu0 = 4.2151088999999996e-10
+ mjd = 0.335
+ mjs = 0.335
+ lua = 7.9060667e-17
+ lub = -2.7964918e-26
+ luc = 5.5424848e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = -2.574678e-15
+ nsd = 1e+20
+ pbd = 0.75
+ pat = -1.0212358e-9
+ wvsat = -0.0016609281000000001
+ pbs = 0.75
+ pk2 = 2.1304022e-16
+ aigbinv = 0.009974
+ wvth0 = 1.32392e-10
+ pu0 = -6.6237547e-17
+ vfbsdoff = 0.01
+ prt = 0
+ pua = -2.0419953e-23
+ pub = 1.469069e-32
+ puc = 1.2609666e-24
+ pud = 0
+ waigc = 6.0357037e-12
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 8.3453493e-9
+ ub1 = -1.1410668e-17
+ pvfbsdoff = 0
+ uc1 = 1.6197295e-9
+ keta = -0.31465021
+ lku0we = 1.8e-11
+ tpb = 0.0016
+ wa0 = -5.9482929e-8
+ epsrox = 3.9
+ ute = -1
+ wat = 0.022486376
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 1.7062889e-10
+ wlc = 0
+ wln = 1
+ wu0 = 1.3607209e-9
+ xgl = -8.2e-9
+ xgw = 0
+ wua = 3.3448805e-16
+ wub = -2.4882066e-25
+ wuc = -1.434288e-17
+ wud = 0
+ lketa = 1.5671934e-8
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ paramchk = 1
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 1.0759785999999998e-10
+ xpart = 1
+ rdsmod = 0
+ kt1l = 0
+ igbmod = 1
+ egidl = 0.001
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ lint = 0
+ poxedge = 1
+ pbswgd = 0.8
+ pbswgs = 0.8
+ lkt1 = 1.1671281e-8
+ lkt2 = 2.350723e-9
+ lmax = 5.233e-8
+ lmin = 4.333e-8
+ ijthdfwd = 0.01
+ igcmod = 1
+ binunit = 2
+ lpe0 = 6.44e-8
+ lpeb = 0
+ minv = -0.33
+ lua1 = -3.7660644e-16
+ lub1 = 5.1040674e-25
+ luc1 = -7.3441373e-17
+ ndep = 1e+18
+ lwlc = 0
+ ijthdrev = 0.01
+ moin = 5.5538
+ nigc = 2.291
+ lpdiblc2 = 0
+ pvoff = 8.9992158e-17
+ cdscb = 0
+ cdscd = 0
+ pvsat = 3.527869999999998e-12
+ noff = 2.2684
+ wk2we = 0.0
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ pvth0 = -2.69772397e-16
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ permod = 1
+ drout = 0.56
+ paigc = -1.4334713e-18
+ voffl = 0
+ ntox = -1.9260000000000002
+ pcit = -1.2266278e-17
+ pclm = 1.8533357
+ weta0 = -4.8483037e-9
+ wetab = 2.5894049e-9
+ lpclm = -6.4524768e-8
+ lkvth0we = 3e-12
+ phin = 0.15
+ voffcv = -0.125
+ wpemod = 1
+ pkt1 = -1.7183146e-15
+ pkt2 = -1.1786798e-16
+ cgidl = 1
+ acnqsmod = 0
+ njtsswg = 6.489
+ rbdb = 50
+ pua1 = 1.8341764e-23
+ prwb = 0
+ pub1 = -1.3009877e-32
+ prwg = 0
+ puc1 = 9.9681375e-24
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ pbswd = 0.9
+ rbpb = 50
+ rbpd = 50
+ pbsws = 0.9
+ rbps = 50
+ rbodymod = 0
+ rbsb = 50
+ pvag = 2.1
+ ckappad = 0.6
+ ckappas = 0.6
+ rdsw = 200
+ pdiblc1 = 0
+ pdiblc2 = 0.0014658889
+ pdiblcb = 0
+ tpbswg = 0.001
+ pdits = 0
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ bigbacc = 0.0054401
+ ptvoff = -2.2999757e-17
+ pk2we = 0.0
+ wpdiblc2 = 1.4741467e-10
+ rshg = 14.1
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ waigsd = 1.9716411e-12
+ kvth0we = -0.00022
+ diomod = 1
+ tnoia = 0
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ pditsd = 0
+ pditsl = 0
+ vtsswgd = 1.1
+ peta0 = -1.06775094e-17
+ vtsswgs = 1.1
+ cjswgd = 1.9367000000000001e-10
+ pku0we = 0.0
+ cjswgs = 1.9367000000000001e-10
+ petab = -2.558443e-17
+ wketa = 3.409679e-8
+ tpbsw = 0.0025
+ tnom = 25
+ cjswd = 5.457e-11
+ cjsws = 5.457e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ tvfbsdoff = 0.1
+ toxe = 2.71e-9
+ toxm = 2.67e-9
+ wkvth0we = 0.0
+ mjswgd = 0.95
+ mjswgs = 0.95
+ wtvfbsdoff = 0
+ tcjswg = 0.00128
+ trnqsmod = 0
+ ltvfbsdoff = 0
+ wags = 2.5054667e-7
+ wcit = 2.8917948e-10
+ scref = 1e-6
+ voff = -0.1005239
+ pigcd = 2.572
+ acde = 0.5
+ aigsd = 0.0063632396
+ nfactor = 1
+ rgatemod = 0
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ tnjtsswg = 1
+ vsat = 81684.56
+ wint = 0
+ lvoff = -3.8177557e-9
+ vth0 = -0.31867124
+ fprout = 200
+ wkt1 = 3.6711578e-8
+ wkt2 = 3.2153756e-9
+ wmax = 2.726e-7
+ xrcrg1 = 12
+ xrcrg2 = 1
+ aigc = 0.0068691843
+ wmin = 1.08e-7
+ lvsat = 0.00099339504
+ lvth0 = -4.3879777000000005e-9
+ ptvfbsdoff = 0
+ delta = 0.018814
+ laigc = -1.683393e-11
+ wtvoff = 5.2119196e-10
+ wua1 = -3.864028e-16
+ wub1 = 3.2172349e-25
+ wuc1 = -2.0479093e-16
+ rnoia = 0
+ rnoib = 0
+ a0 = 3.0243356
+ a1 = 0
+ a2 = 1
+ nigbacc = 10
+ b0 = 0
+ b1 = 0
+ at = -187272.02
+ cf = 7.598099999999999e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.021495622
+ k3 = -2.5823
+ em = 20000000.0
+ bigc = 0.0012521
+ ll = 0
+ lw = 0
+ u0 = -0.00018459259
+ w0 = 0
+ wwlc = 0
+ ua = -1.9655718e-9
+ ub = 1.5789686e-18
+ uc = -2.0243416e-10
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 5.6700000000000005e-9
+ ww = 0
+ xw = 3.4e-9
+ pketa = -2.1465872e-15
+ ngate = 1.7e+20
+ ngcon = 1
+ capmod = 2
+ wpclm = -1.4226467e-7
+ cdsc = 0
+ cgbo = 0
+ cgdl = 2.799765e-11
+ cgdo = 2.4628259999999997e-11
+ wku0we = 1.5e-11
+ xtid = 3
+ xtis = 3
+ gbmin = 1e-12
+ nigbinv = 2.171
+ cgsl = 2.799765e-11
+ cgso = 2.4628259999999997e-11
+ cigc = 0.15259
+ jswgd = 3.69e-13
+ mobmod = 0
+ jswgs = 3.69e-13
+ )

.model pch_ss_40 pmos (
+ level = 54
+ fnoimod = 1
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ eigbinv = 1.1
+ laigsd = 6.1219753e-16
+ k2we = 5e-5
+ ijthsfwd = 0.01
+ tvoff = -0.00058332606
+ dsub = 0.5
+ dtox = 3.91e-10
+ xjbvd = 1
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ xjbvs = 1
+ lk2we = 0.0
+ eta0 = 0.19272491
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ etab = -0.15063456
+ ijthsrev = 0.01
+ cigbacc = 0.245
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = -2.4311511e-9
+ letab = 4.3496496e-9
+ tnoimod = 0
+ ppclm = -3.5647768e-15
+ dlcig = 2.5e-9
+ cigbinv = 0.006
+ bgidl = 1834800000.0
+ ppdiblc2 = 0
+ toxref = 3e-9
+ version = 4.5
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ tempmod = 0
+ ags = 1.2522222
+ cjd = 0.00144022
+ cit = -0.0098195899
+ cjs = 0.00144022
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 4.0349e-9
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ aigbacc = 0.012071
+ bigsd = 0.0003327
+ pkvth0we = 0.0
+ la0 = -3.4726683e-8
+ ltvoff = 1.026653e-10
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0.0027111306999999998
+ kt1 = -0.31430817
+ kt2 = -0.12562663
+ lk2 = 6.6841473e-9
+ wvoff = 3.3909703e-9
+ llc = 0
+ lln = 1
+ lu0 = 5.3141728e-10
+ mjd = 0.335
+ mjs = 0.335
+ lua = 9.0470184e-17
+ lub = -2.7144874e-26
+ luc = 2.7216576e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 1.4761752e-15
+ nsd = 1e+20
+ pbd = 0.75
+ pat = -5.6834015e-11
+ wvsat = -0.011345602
+ pbs = 0.75
+ pk2 = -2.7720832e-16
+ aigbinv = 0.009974
+ wvth0 = 1.2795535899999999e-9
+ pu0 = -6.1923224e-17
+ vfbsdoff = 0.01
+ prt = 0
+ pua = -4.2432063e-24
+ pub = -5.3708285e-33
+ puc = -1.7176927e-24
+ pud = 0
+ waigc = -4.0606639e-11
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 2.1566906e-9
+ ub1 = -3.7269546e-18
+ pvfbsdoff = 0
+ uc1 = -1.7258848e-10
+ keta = 0.15497942
+ lku0we = 1.8e-11
+ tpb = 0.0016
+ wa0 = -1.421534e-7
+ epsrox = 3.9
+ ute = -1
+ wat = 0.002804707
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 1.0175701e-8
+ wlc = 0
+ wln = 1
+ wu0 = 1.2726735e-9
+ xgl = -8.2e-9
+ xgw = 0
+ wua = 4.3503521e-18
+ wub = 1.6059812e-25
+ wuc = 4.6446086e-17
+ wud = 0
+ lketa = -7.3399177e-9
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ paramchk = 1
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 5.8206353e-10
+ xpart = 1
+ rdsmod = 0
+ kt1l = 0
+ igbmod = 1
+ egidl = 0.001
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ lint = 0
+ poxedge = 1
+ pbswgd = 0.8
+ pbswgs = 0.8
+ lkt1 = 6.363929e-10
+ lkt2 = 2.3369169e-9
+ lmax = 4.333e-8
+ lmin = 3.6e-8
+ ijthdfwd = 0.01
+ igcmod = 1
+ binunit = 2
+ lpe0 = 6.44e-8
+ lpeb = 0
+ minv = -0.33
+ lua1 = -7.3362164e-17
+ lub1 = 1.3390478e-25
+ luc1 = 1.4382206e-17
+ ndep = 1e+18
+ lwlc = 0
+ ijthdrev = 0.01
+ moin = 5.5538
+ nigc = 2.291
+ paigsd = -6.9790518e-23
+ lpdiblc2 = 0
+ pvoff = -6.9138231e-17
+ cdscb = 0
+ cdscd = 0
+ pvsat = 4.7807606e-10
+ noff = 2.2684
+ wk2we = 0.0
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ pvth0 = -3.2598297e-16
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ permod = 1
+ drout = 0.56
+ paigc = 8.520035e-19
+ voffl = 0
+ ntox = -1.9260000000000002
+ pcit = -4.0436162e-17
+ pclm = 0.41497396
+ weta0 = -1.0107776999999999e-8
+ wetab = 1.1541057e-8
+ lpclm = 5.9549575e-9
+ lkvth0we = 3e-12
+ phin = 0.15
+ voffcv = -0.125
+ wpemod = 1
+ pkt1 = -1.7140714e-15
+ pkt2 = -7.0509572e-16
+ cgidl = 1
+ acnqsmod = 0
+ njtsswg = 6.489
+ rbdb = 50
+ pua1 = 3.2441676e-23
+ prwb = 0
+ pub1 = -5.4663004e-32
+ prwg = 0
+ puc1 = -1.3788915e-24
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ pbswd = 0.9
+ rbpb = 50
+ rbpd = 50
+ pbsws = 0.9
+ rbps = 50
+ rbodymod = 0
+ rbsb = 50
+ pvag = 2.1
+ ckappad = 0.6
+ ckappas = 0.6
+ rdsw = 200
+ pdiblc1 = 0
+ pdiblc2 = 0.0014658889
+ pdiblcb = 0
+ tpbswg = 0.001
+ pdits = 0
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ bigbacc = 0.0054401
+ ptvoff = -3.9364956e-17
+ pk2we = 0.0
+ wpdiblc2 = 1.4741467e-10
+ rshg = 14.1
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ waigsd = 1.9730654e-12
+ kvth0we = -0.00022
+ diomod = 1
+ tnoia = 0
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ pditsd = 0
+ pditsl = 0
+ vtsswgd = 1.1
+ peta0 = 2.4703678e-16
+ vtsswgs = 1.1
+ cjswgd = 1.9367000000000001e-10
+ pku0we = 0.0
+ cjswgs = 1.9367000000000001e-10
+ petab = -4.6421536e-16
+ wketa = -5.7187654e-8
+ tpbsw = 0.0025
+ tnom = 25
+ cjswd = 5.457e-11
+ cjsws = 5.457e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ tvfbsdoff = 0.1
+ toxe = 2.71e-9
+ toxm = 2.67e-9
+ wkvth0we = 0.0
+ mjswgd = 0.95
+ mjswgs = 0.95
+ wtvfbsdoff = 0
+ tcjswg = 0.00128
+ trnqsmod = 0
+ ltvfbsdoff = 0
+ wags = 2.5054667e-7
+ wcit = 8.6407259e-10
+ scref = 1e-6
+ voff = -0.12231559
+ pigcd = 2.572
+ acde = 0.5
+ aigsd = 0.0063632271
+ nfactor = 1
+ rgatemod = 0
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ tnjtsswg = 1
+ vsat = 171956.58000000002
+ wint = 0
+ lvoff = -2.7499629e-9
+ vth0 = -0.37839467000000004
+ fprout = 200
+ wkt1 = 3.6624982e-8
+ wkt2 = 1.5199615e-8
+ wmax = 2.726e-7
+ xrcrg1 = 12
+ xrcrg2 = 1
+ aigc = 0.0069354083
+ wmin = 1.08e-7
+ lvsat = -0.0034299414
+ lvth0 = -1.4615239000000001e-9
+ ptvfbsdoff = 0
+ delta = 0.018814
+ laigc = -2.0078906e-11
+ wtvoff = 8.5517561e-10
+ wua1 = -6.7415611e-16
+ wub1 = 1.1717873e-24
+ wuc1 = 2.6781086e-17
+ rnoia = 0
+ rnoib = 0
+ a0 = 0.69140412
+ a1 = 0
+ a2 = 1
+ nigbacc = 10
+ b0 = 0
+ b1 = 0
+ at = -30917.36
+ cf = 7.598099999999999e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.06369048
+ k3 = -2.5823
+ em = 20000000.0
+ bigc = 0.0012521
+ ll = 0
+ lw = 0
+ u0 = -0.0024275803
+ w0 = 0
+ wwlc = 0
+ ua = -2.1984191e-9
+ ub = 1.5622339e-18
+ uc = -1.4486626e-10
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 5.6700000000000005e-9
+ ww = 0
+ xw = 3.4e-9
+ pketa = 2.3263506e-15
+ ngate = 1.7e+20
+ ngcon = 1
+ capmod = 2
+ wpclm = 8.9861524e-8
+ cdsc = 0
+ cgbo = 0
+ cgdl = 2.799765e-11
+ cgdo = 2.4628259999999997e-11
+ wku0we = 1.5e-11
+ xtid = 3
+ xtis = 3
+ gbmin = 1e-12
+ nigbinv = 2.171
+ cgsl = 2.799765e-11
+ cgso = 2.4628259999999997e-11
+ cigc = 0.15259
+ jswgd = 3.69e-13
+ mobmod = 0
+ jswgs = 3.69e-13
+ )

.model pch_tt_1 pmos (
+ level = 54
+ ppclm = 0
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ bigbacc = 0.0054401
+ wpdiblc2 = 0
+ tnom = 25
+ kvth0we = -0.00022
+ tvfbsdoff = 0.1
+ dmcgt = 0
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ tcjsw = 9.34e-5
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ toxref = 3e-9
+ bigsd = 0.0003327
+ wkvth0we = 0.0
+ wvoff = 0
+ trnqsmod = 0
+ voff = -0.11110337
+ acde = 0.5
+ wvsat = 0
+ wvfbsdoff = 0
+ wvth0 = 0.0
+ lvfbsdoff = 0
+ vsat = 120000
+ wint = 0
+ vth0 = -0.38513527
+ ltvoff = 0
+ wmax = 0.00090001
+ aigc = 0.0068307507
+ wmin = 9e-6
+ a0 = 2.531
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 72000
+ cf = 8.17e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.00077592763
+ k3 = -2.5823
+ em = 20000000.0
+ lketa = 0
+ ll = 0
+ lw = 0
+ u0 = 0.009795
+ w0 = 0
+ rgatemod = 0
+ ua = 1.297e-10
+ ub = 1.182572e-18
+ uc = 2.014e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xpart = 1
+ xw = 6e-9
+ nfactor = 1
+ tnjtsswg = 1
+ lku0we = 1.8e-11
+ bigc = 0.0012521
+ egidl = 0.001
+ wwlc = 0
+ epsrox = 3.9
+ cdsc = 0
+ rdsmod = 0
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ igbmod = 1
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigc = 0.15259
+ nigbacc = 10
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ pbswgd = 0.8
+ pbswgs = 0.8
+ igcmod = 1
+ nigbinv = 2.171
+ pvoff = 0
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ cdscb = 0
+ cdscd = 0
+ pvsat = 0
+ wk2we = 0.0
+ pvth0 = 0.0
+ drout = 0.56
+ k2we = 5e-5
+ dsub = 0.5
+ dtox = 3.91e-10
+ voffl = 0
+ fnoimod = 1
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ eigbinv = 1.1
+ weta0 = 0
+ permod = 1
+ lpclm = 0
+ eta0 = 0.1672
+ etab = -0.23
+ ijthsfwd = 0.01
+ cgidl = 1
+ voffcv = -0.125
+ wpemod = 1
+ ijthsrev = 0.01
+ pbswd = 0.9
+ pbsws = 0.9
+ cigbacc = 0.245
+ tnoimod = 0
+ pdits = 0
+ cigsd = 0.013281
+ cigbinv = 0.006
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ ppdiblc2 = 0
+ tpbswg = 0.001
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ version = 4.5
+ tempmod = 0
+ tnoia = 0
+ peta0 = 0
+ ptvoff = 0
+ aigbacc = 0.012071
+ tpbsw = 0.0025
+ pkvth0we = 0.0
+ pvfbsdoff = 0
+ keta = -0.042350111
+ cjswd = 5.1e-11
+ cjsws = 5.1e-11
+ diomod = 1
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ pditsd = 0
+ pditsl = 0
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ cjswgd = 1.81e-10
+ pku0we = 0.0
+ cjswgs = 1.81e-10
+ lcit = 0
+ aigbinv = 0.009974
+ vfbsdoff = 0.01
+ wtvfbsdoff = 0
+ kt1l = 0
+ lint = 6.5375218e-9
+ ltvfbsdoff = 0
+ mjswgd = 0.95
+ mjswgs = 0.95
+ lkt1 = 0
+ paramchk = 1
+ lmax = 2.001e-5
+ lmin = 8.9991e-6
+ tcjswg = 0.00128
+ scref = 1e-6
+ lpe0 = 6.44e-8
+ lpeb = 0
+ pigcd = 2.572
+ aigsd = 0.0063636
+ minv = -0.33
+ lvoff = 0
+ poxedge = 1
+ ndep = 1e+18
+ lwlc = 0
+ ijthdfwd = 0.01
+ lvsat = 0
+ moin = 5.5538
+ lvth0 = 0.0
+ binunit = 2
+ ptvfbsdoff = 0
+ nigc = 2.291
+ delta = 0.018814
+ rnoia = 0
+ rnoib = 0
+ fprout = 200
+ noff = 2.2684
+ ags = 0.8379228
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ ijthdrev = 0.01
+ ngate = 1.7e+20
+ cjd = 0.001346
+ cit = 5e-6
+ cjs = 0.001346
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 1.0572421799999999e-8
+ ngcon = 1
+ k3b = 2.1176
+ wpclm = 0
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ lpdiblc2 = 0
+ ntox = 1
+ wtvoff = 0
+ pcit = 0
+ pclm = 1.484
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ la0 = 0
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0
+ kt1 = -0.17107633
+ lk2 = 0
+ kt2 = -0.04747
+ jtsswgd = 1.75e-7
+ phin = 0.15
+ llc = 0
+ jtsswgs = 1.75e-7
+ lln = 1
+ lu0 = 0
+ mjd = 0.335
+ mjs = 0.335
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 0
+ capmod = 2
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ pk2 = 0
+ pkt1 = 0
+ pu0 = 0
+ prt = 0
+ wku0we = 1.5e-11
+ pud = 0
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 1.1969344e-9
+ ub1 = -1.3666143e-18
+ uc1 = 6.873e-11
+ mobmod = 0
+ tpb = 0.0016
+ wa0 = 0
+ lkvth0we = 3e-12
+ ute = -1
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 0
+ wlc = 0
+ wln = 1
+ rbdb = 50
+ prwb = 0
+ wu0 = 0
+ prwg = 0
+ xgl = -8.2e-9
+ xgw = 0
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ rdsw = 200
+ tvoff = 0.0026155642
+ acnqsmod = 0
+ njtsswg = 6.489
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ xtsswgd = 0.32
+ rbodymod = 0
+ xtsswgs = 0.32
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.0026729629
+ ku0we = -0.0007
+ pdiblcb = 0
+ beta0 = 13.32
+ rshg = 14.1
+ leta0 = 0
+ )

.model pch_tt_2 pmos (
+ level = 54
+ aigbinv = 0.009974
+ eta0 = 0.1672
+ tnoia = 0
+ etab = -0.23
+ ijthdfwd = 0.01
+ peta0 = 0
+ toxref = 3e-9
+ pvfbsdoff = 0
+ tpbsw = 0.0025
+ cjswd = 5.1e-11
+ cjsws = 5.1e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ ijthdrev = 0.01
+ lpdiblc2 = 7.1311563e-9
+ poxedge = 1
+ ltvoff = -4.7585658e-10
+ binunit = 2
+ scref = 1e-6
+ pigcd = 2.572
+ aigsd = 0.0063636
+ lku0we = 1.8e-11
+ epsrox = 3.9
+ lkvth0we = 3e-12
+ lvoff = -8.0044387e-9
+ lvsat = 0
+ rdsmod = 0
+ lvth0 = -5.1267661e-9
+ ags = 0.80385259
+ igbmod = 1
+ delta = 0.018814
+ laigc = -4.8397409e-11
+ cjd = 0.001346
+ cit = 5e-6
+ cjs = 0.001346
+ clc = 1e-7
+ cle = 0.6
+ acnqsmod = 0
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 1.0572421799999999e-8
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ k3b = 2.1176
+ rnoia = 0
+ rnoib = 0
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ keta = -0.040853613
+ pbswgd = 0.8
+ pbswgs = 0.8
+ rbodymod = 0
+ a0 = 2.5747309
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 72000
+ lags = 3.062912e-7
+ ngate = 1.7e+20
+ cf = 8.17e-11
+ igcmod = 1
+ la0 = -3.9314047e-7
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.0012551498
+ k3 = -2.5823
+ em = 20000000.0
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0
+ ll = 0
+ lw = 0
+ kt1 = -0.16652617
+ kt2 = -0.046491549
+ lk2 = 4.3082075e-9
+ u0 = 0.0097948901
+ ngcon = 1
+ w0 = 0
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ ua = 1.4083134e-10
+ ub = 1.1675774e-18
+ uc = 1.8373185e-11
+ ud = 0
+ llc = 0
+ wpclm = 0
+ lln = 1
+ lcit = 0
+ wl = 0
+ wr = 1
+ lu0 = 9.8779012e-13
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 6e-9
+ mjd = 0.335
+ mjs = 0.335
+ lua = -1.0007073e-16
+ lub = 1.3480174e-25
+ luc = 1.5883665e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ kt1l = 0
+ njs = 1.02
+ pa0 = 0
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ pk2 = 0
+ gbmin = 1e-12
+ pu0 = 0
+ jswgd = 3.69e-13
+ prt = 0
+ jswgs = 3.69e-13
+ pud = 0
+ lint = 6.5375218e-9
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 1.1817684e-9
+ ub1 = -1.3634053e-18
+ uc1 = 6.7786161e-11
+ tpb = 0.0016
+ lkt1 = -4.0906013e-8
+ lkt2 = -8.7962711e-9
+ wa0 = 0
+ lmax = 8.9991e-6
+ ute = -1
+ lmin = 8.9908e-7
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 0
+ wlc = 0
+ wln = 1
+ wu0 = 0
+ xgl = -8.2e-9
+ xgw = 0
+ njtsswg = 6.489
+ lpe0 = 6.44e-8
+ wud = 0
+ wpdiblc2 = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ lpeb = 0
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ minv = -0.33
+ lua1 = 1.3634229e-16
+ lub1 = -2.8849398e-26
+ luc1 = 8.4851172e-18
+ permod = 1
+ ckappad = 0.6
+ ckappas = 0.6
+ ndep = 1e+18
+ pdiblc1 = 0
+ pdiblc2 = 0.0018797309
+ pdiblcb = 0
+ lwlc = 0
+ moin = 5.5538
+ nigc = 2.291
+ tvoff = 0.002668496
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ wkvth0we = 0.0
+ voffcv = -0.125
+ wpemod = 1
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ bigbacc = 0.0054401
+ trnqsmod = 0
+ ku0we = -0.0007
+ beta0 = 13.32
+ kvth0we = -0.00022
+ ntox = 1
+ pcit = 0
+ pclm = 1.484
+ leta0 = 0
+ lintnoi = -5e-9
+ ppclm = 0
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ phin = 0.15
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ pkt1 = 0
+ rgatemod = 0
+ tpbswg = 0.001
+ tnjtsswg = 1
+ tvfbsdoff = 0.1
+ dmcgt = 0
+ rbdb = 50
+ tcjsw = 9.34e-5
+ prwb = 0
+ prwg = 0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ ptvoff = 0
+ wtvfbsdoff = 0
+ rdsw = 200
+ bigsd = 0.0003327
+ diomod = 1
+ ltvfbsdoff = 0
+ pditsd = 0
+ pditsl = 0
+ nfactor = 1
+ wvoff = 0
+ cjswgd = 1.81e-10
+ pku0we = 0.0
+ cjswgs = 1.81e-10
+ wvfbsdoff = 0
+ wvsat = 0
+ lvfbsdoff = 0
+ wvth0 = 0.0
+ rshg = 14.1
+ mjswgd = 0.95
+ mjswgs = 0.95
+ tcjswg = 0.00128
+ lketa = -1.3453518e-8
+ ptvfbsdoff = 0
+ nigbacc = 10
+ xpart = 1
+ tnom = 25
+ egidl = 0.001
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ ijthsfwd = 0.01
+ nigbinv = 2.171
+ fprout = 200
+ xrcrg1 = 12
+ xrcrg2 = 1
+ ijthsrev = 0.01
+ fnoimod = 1
+ voff = -0.110213
+ wtvoff = 0
+ acde = 0.5
+ eigbinv = 1.1
+ pvoff = 0
+ vsat = 120000
+ wint = 0
+ vth0 = -0.384565
+ cdscb = 0
+ cdscd = 0
+ wmax = 0.00090001
+ pvsat = 0
+ aigc = 0.0068361342
+ wmin = 9e-6
+ wk2we = 0.0
+ capmod = 2
+ pvth0 = 0.0
+ drout = 0.56
+ wku0we = 1.5e-11
+ ppdiblc2 = 0
+ mobmod = 0
+ voffl = 0
+ bigc = 0.0012521
+ weta0 = 0
+ cigbacc = 0.245
+ wwlc = 0
+ lpclm = 0
+ cdsc = 0
+ tnoimod = 0
+ cgbo = 0
+ cgidl = 1
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigc = 0.15259
+ pkvth0we = 0.0
+ cigbinv = 0.006
+ pbswd = 0.9
+ pbsws = 0.9
+ vfbsdoff = 0.01
+ version = 4.5
+ tempmod = 0
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ pdits = 0
+ cigsd = 0.013281
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ dvt0w = 0
+ paramchk = 1
+ dvt1w = 0
+ dvt2w = 0
+ aigbacc = 0.012071
+ k2we = 5e-5
+ dsub = 0.5
+ dtox = 3.91e-10
+ pk2we = 0.0
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ )

.model pch_tt_3 pmos (
+ level = 54
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ nigbacc = 10
+ ijthsrev = 0.01
+ wvoff = 0
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ wvsat = 0
+ ntox = 1
+ wvth0 = 0.0
+ pcit = 0
+ pclm = 1.484
+ ltvoff = -2.3123852e-10
+ nigbinv = 2.171
+ phin = 0.15
+ lketa = -1.5940244e-8
+ pkt1 = 0
+ ppdiblc2 = 0
+ xpart = 1
+ lku0we = 1.8e-11
+ epsrox = 3.9
+ egidl = 0.001
+ rbdb = 50
+ fnoimod = 1
+ prwb = 0
+ prwg = 0
+ rdsmod = 0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ eigbinv = 1.1
+ igbmod = 1
+ rdsw = 200
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ pbswgd = 0.8
+ pbswgs = 0.8
+ pkvth0we = 0.0
+ igcmod = 1
+ vfbsdoff = 0.01
+ rshg = 14.1
+ cigbacc = 0.245
+ pvoff = 0
+ cdscb = 0
+ cdscd = 0
+ pvsat = 0
+ tnoimod = 0
+ wk2we = 0.0
+ pvth0 = 0.0
+ paramchk = 1
+ drout = 0.56
+ cigbinv = 0.006
+ voffl = 0
+ permod = 1
+ tnom = 25
+ weta0 = 0
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ a0 = 2.8917556
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ lpclm = 0
+ at = 72000
+ cf = 8.17e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = 0.0040664684
+ k3 = -2.5823
+ em = 20000000.0
+ ijthdfwd = 0.01
+ version = 4.5
+ ll = 0
+ lw = 0
+ u0 = 0.010026756
+ w0 = 0
+ ua = 1.1413788e-10
+ ub = 1.1978347e-18
+ uc = 4.3035111e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 6e-9
+ tempmod = 0
+ cgidl = 1
+ voffcv = -0.125
+ wpemod = 1
+ aigbacc = 0.012071
+ ijthdrev = 0.01
+ pbswd = 0.9
+ pbsws = 0.9
+ voff = -0.10886793
+ lpdiblc2 = 1.7469722e-9
+ acde = 0.5
+ vsat = 120000
+ aigbinv = 0.009974
+ wint = 0
+ vth0 = -0.38718963
+ pdits = 0
+ cigsd = 0.013281
+ wmax = 0.00090001
+ aigc = 0.00683106
+ wmin = 9e-6
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ wtvfbsdoff = 0
+ tpbswg = 0.001
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ ltvfbsdoff = 0
+ lkvth0we = 3e-12
+ bigc = 0.0012521
+ wwlc = 0
+ tnoia = 0
+ ptvoff = 0
+ poxedge = 1
+ cdsc = 0
+ peta0 = 0
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ acnqsmod = 0
+ pvfbsdoff = 0
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigc = 0.15259
+ binunit = 2
+ diomod = 1
+ tpbsw = 0.0025
+ cjswd = 5.1e-11
+ cjsws = 5.1e-11
+ mjswd = 0.01
+ pditsd = 0
+ mjsws = 0.01
+ pditsl = 0
+ rbodymod = 0
+ agidl = 3.2166e-9
+ cjswgd = 1.81e-10
+ pku0we = 0.0
+ cjswgs = 1.81e-10
+ ptvfbsdoff = 0
+ dmcg = 3.1e-8
+ mjswgd = 0.95
+ dmci = 3.1e-8
+ dmdg = 0
+ mjswgs = 0.95
+ tcjswg = 0.00128
+ k2we = 5e-5
+ jtsswgd = 1.75e-7
+ scref = 1e-6
+ jtsswgs = 1.75e-7
+ wpdiblc2 = 0
+ dsub = 0.5
+ pigcd = 2.572
+ dtox = 3.91e-10
+ aigsd = 0.0063635603
+ ags = 0.82774541
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ lvoff = -9.201547e-9
+ cjd = 0.001346
+ cit = -8.7888889e-5
+ cjs = 0.001346
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 1.0572421799999999e-8
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ eta0 = 0.1672
+ etab = -0.23
+ lvsat = 0
+ lvth0 = -2.7908401e-9
+ delta = 0.018814
+ laigc = -4.3881382e-11
+ la0 = -6.7529244e-7
+ fprout = 200
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0
+ kt1 = -0.19559142
+ kt2 = -0.048919444
+ lk2 = -4.2803272e-10
+ llc = 0
+ lln = 1
+ lu0 = -2.0537244e-10
+ rnoia = 0
+ rnoib = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ mjd = 0.335
+ mjs = 0.335
+ lua = -7.6313554e-17
+ lub = 1.0787275e-25
+ luc = -6.0654489e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ wkvth0we = 0.0
+ njs = 1.02
+ pa0 = 0
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ pk2 = 0
+ njtsswg = 6.489
+ pu0 = 0
+ prt = 0
+ pud = 0
+ ngate = 1.7e+20
+ trnqsmod = 0
+ wtvoff = 0
+ ngcon = 1
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 1.2804108e-9
+ ub1 = -1.1625424e-18
+ uc1 = 4.6637333e-11
+ wpclm = 0
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ tpb = 0.0016
+ wa0 = 0
+ ute = -1
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 0
+ ckappad = 0.6
+ ckappas = 0.6
+ gbmin = 1e-12
+ wlc = 0
+ wln = 1
+ wu0 = 0
+ xgl = -8.2e-9
+ xgw = 0
+ pdiblc1 = 0
+ pdiblc2 = 0.0079293759
+ wud = 0
+ jswgd = 3.69e-13
+ wwc = 0
+ jswgs = 3.69e-13
+ wwl = 0
+ wwn = 1
+ pdiblcb = 0
+ capmod = 2
+ wku0we = 1.5e-11
+ rgatemod = 0
+ mobmod = 0
+ tnjtsswg = 1
+ bigbacc = 0.0054401
+ kvth0we = -0.00022
+ lintnoi = -5e-9
+ tvoff = 0.0023936443
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ laigsd = 3.5374533e-14
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ keta = -0.03805954
+ lags = 2.8502658e-7
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 8.2671111e-11
+ ku0we = -0.0007
+ beta0 = 13.32
+ kt1l = 0
+ leta0 = 0
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ ppclm = 0
+ lint = 6.5375218e-9
+ lkt1 = -1.5037939e-8
+ lkt2 = -6.6354444e-9
+ dlcig = 2.5e-9
+ lmax = 8.9908e-7
+ bgidl = 1834800000.0
+ lmin = 4.4908e-7
+ lpe0 = 6.44e-8
+ lpeb = 0
+ tvfbsdoff = 0.1
+ minv = -0.33
+ lua1 = 4.8550568e-17
+ nfactor = 1
+ lub1 = -2.0761736e-25
+ luc1 = 2.7307573e-17
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ ndep = 1e+18
+ lwlc = 0
+ ijthsfwd = 0.01
+ moin = 5.5538
+ nigc = 2.291
+ toxref = 3e-9
+ bigsd = 0.0003327
+ )

.model pch_tt_4 pmos (
+ level = 54
+ aigc = 0.0067884199
+ wmin = 9e-6
+ cjd = 0.001346
+ cit = -0.00054497817
+ cjs = 0.001346
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 1.38228675e-8
+ scref = 1e-6
+ k3b = 2.1176
+ rgatemod = 0
+ lku0we = 1.8e-11
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ pigcd = 2.572
+ tnjtsswg = 1
+ epsrox = 3.9
+ aigsd = 0.0063636407
+ njtsswg = 6.489
+ lvoff = -3.8830249e-9
+ bigc = 0.0012521
+ la0 = -4.3379389e-8
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0
+ rdsmod = 0
+ kt1 = -0.2000222
+ kt2 = -0.054670852
+ lk2 = 1.3630221e-9
+ wwlc = 0
+ llc = -1.18e-13
+ xtsswgd = 0.32
+ lln = 0.7
+ xtsswgs = 0.32
+ lu0 = -4.832545e-10
+ igbmod = 1
+ mjd = 0.335
+ mjs = 0.335
+ lua = -1.5477844e-16
+ lub = 5.0676856e-26
+ luc = -5.2541764e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ lvsat = 0
+ njd = 1.02
+ njs = 1.02
+ pa0 = 0
+ lvth0 = 4.3404654e-9
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ ckappad = 0.6
+ pk2 = 0
+ ckappas = 0.6
+ cdsc = 0
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ pu0 = 0
+ pdiblc1 = 0
+ pdiblc2 = 0.013802718
+ delta = 0.018814
+ cgbo = 0
+ prt = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ pud = 0
+ pdiblcb = 0
+ xtid = 3
+ xtis = 3
+ laigc = -2.5119727e-11
+ pbswgd = 0.8
+ pbswgs = 0.8
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ rsh = 15.2
+ tcj = 0.000832
+ cigc = 0.15259
+ ua1 = 1.2553592e-9
+ ub1 = -1.2671808e-18
+ uc1 = 1.0455371e-10
+ rnoia = 0
+ rnoib = 0
+ tpb = 0.0016
+ wa0 = 0
+ igcmod = 1
+ ute = -1
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 0
+ wlc = 0
+ wln = 1
+ wu0 = 0
+ xgl = -8.2e-9
+ xgw = 0
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ ngate = 1.7e+20
+ ngcon = 1
+ wpclm = 0
+ bigbacc = 0.0054401
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ kvth0we = -0.00022
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ k2we = 5e-5
+ vtsswgs = 1.1
+ dsub = 0.5
+ dtox = 3.91e-10
+ permod = 1
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ eta0 = 0.1672
+ ijthsfwd = 0.01
+ etab = -0.23
+ tvoff = 0.002134918
+ voffcv = -0.125
+ wpemod = 1
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ ijthsrev = 0.01
+ wtvfbsdoff = 0
+ ku0we = -0.0007
+ beta0 = 13.32
+ nfactor = 1
+ leta0 = 0
+ ltvfbsdoff = 0
+ ppclm = 0
+ a0 = 1.4555895
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 72000
+ cf = 8.17e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -4.1106394e-6
+ k3 = -2.5823
+ em = 20000000.0
+ ll = -1.18e-13
+ dlcig = 2.5e-9
+ lw = 0
+ u0 = 0.010658306
+ w0 = 0
+ tpbswg = 0.001
+ ua = 2.9246716e-10
+ ub = 1.3278253e-18
+ uc = 4.119131e-11
+ ud = 0
+ bgidl = 1834800000.0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 6e-9
+ ppdiblc2 = 0
+ tvfbsdoff = 0.1
+ nigbacc = 10
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ ptvoff = 0
+ ptvfbsdoff = 0
+ diomod = 1
+ nigbinv = 2.171
+ pkvth0we = 0.0
+ bigsd = 0.0003327
+ keta = -0.029364427
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.81e-10
+ pku0we = 0.0
+ cjswgs = 1.81e-10
+ wvoff = 0
+ lags = 5.4107004e-7
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 2.8379039e-10
+ vfbsdoff = 0.01
+ wvsat = 0
+ kt1l = 0
+ wvth0 = 0.0
+ mjswgd = 0.95
+ mjswgs = 0.95
+ fnoimod = 1
+ eigbinv = 1.1
+ tcjswg = 0.00128
+ lint = 9.7879675e-9
+ lkt1 = -1.3088393e-8
+ lkt2 = -4.1048253e-9
+ paramchk = 1
+ lmax = 4.4908e-7
+ lmin = 2.1577e-7
+ lketa = -1.9766093e-8
+ lpe0 = 6.44e-8
+ xpart = 1
+ lpeb = 0
+ minv = -0.33
+ lua1 = 5.9573279e-17
+ lub1 = -1.6157647e-25
+ egidl = 0.001
+ luc1 = 1.8243668e-18
+ ndep = 1e+18
+ lwlc = 0
+ ijthdfwd = 0.01
+ moin = 5.5538
+ cigbacc = 0.245
+ fprout = 200
+ nigc = 2.291
+ xrcrg1 = 12
+ xrcrg2 = 1
+ tnoimod = 0
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ ijthdrev = 0.01
+ cigbinv = 0.006
+ wtvoff = 0
+ lpdiblc2 = -8.3729822e-10
+ ntox = 1
+ pcit = 0
+ pclm = 1.484
+ pvoff = 0
+ capmod = 2
+ version = 4.5
+ cdscb = 0
+ cdscd = 0
+ pvsat = 0
+ phin = 0.15
+ wku0we = 1.5e-11
+ tempmod = 0
+ wk2we = 0.0
+ pvth0 = 0.0
+ drout = 0.56
+ mobmod = 0
+ pkt1 = 0
+ voffl = 0
+ aigbacc = 0.012071
+ lkvth0we = 3e-12
+ weta0 = 0
+ rbdb = 50
+ prwb = 0
+ prwg = 0
+ lpclm = 0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ rdsw = 200
+ aigbinv = 0.009974
+ cgidl = 1
+ acnqsmod = 0
+ rbodymod = 0
+ pbswd = 0.9
+ pbsws = 0.9
+ rshg = 14.1
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ pdits = 0
+ poxedge = 1
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ binunit = 2
+ wpdiblc2 = 0
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ tnom = 25
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ tnoia = 0
+ toxref = 3e-9
+ peta0 = 0
+ pvfbsdoff = 0
+ tpbsw = 0.0025
+ wkvth0we = 0.0
+ cjswd = 5.1e-11
+ cjsws = 5.1e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ trnqsmod = 0
+ voff = -0.12095548
+ acde = 0.5
+ ltvoff = -1.1739897e-10
+ vsat = 120000
+ wint = 0
+ vth0 = -0.40339715
+ wmax = 0.00090001
+ ags = 0.24582847
+ )

.model pch_tt_5 pmos (
+ level = 54
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ pbswgd = 0.8
+ pbswgs = 0.8
+ acnqsmod = 0
+ version = 4.5
+ tempmod = 0
+ igcmod = 1
+ keta = -0.12863898
+ rbodymod = 0
+ lags = 3.2185083e-8
+ aigbacc = 0.012071
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 7.5945573e-11
+ kt1l = 0
+ pvoff = 0
+ cdscb = 0
+ cdscd = 0
+ lint = 9.7879675e-9
+ pvsat = 0.0
+ wk2we = 0.0
+ pvth0 = 0.0
+ aigbinv = 0.009974
+ lkt1 = -4.7409966e-9
+ lkt2 = -5.2805906e-10
+ drout = 0.56
+ lmax = 2.1577e-7
+ lmin = 9e-8
+ wpdiblc2 = 0
+ lpe0 = 6.44e-8
+ permod = 1
+ lpeb = 0
+ voffl = 0
+ minv = -0.33
+ lua1 = -1.5051887e-16
+ lub1 = 1.742578e-25
+ luc1 = 7.2216103e-18
+ weta0 = 0
+ ndep = 1e+18
+ lpclm = -1.4239795e-8
+ wtvfbsdoff = 0
+ lwlc = 0
+ moin = 5.5538
+ cgidl = 1
+ voffcv = -0.125
+ wpemod = 1
+ nigc = 2.291
+ ltvfbsdoff = 0
+ poxedge = 1
+ wkvth0we = 0.0
+ noff = 2.2684
+ binunit = 2
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ pbswd = 0.9
+ pbsws = 0.9
+ trnqsmod = 0
+ ntox = 1
+ pcit = 0.0
+ pclm = 1.5514872
+ pdits = 0
+ cigsd = 0.013281
+ phin = 0.15
+ tpbswg = 0.001
+ ptvfbsdoff = 0
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ pkt1 = 0
+ rgatemod = 0
+ tnjtsswg = 1
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ ptvoff = 0
+ rbdb = 50
+ prwb = 0
+ prwg = 0
+ tnoia = 0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ pvfbsdoff = 0
+ rdsw = 200
+ peta0 = 0
+ diomod = 1
+ tpbsw = 0.0025
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.81e-10
+ pku0we = 0.0
+ cjswgs = 1.81e-10
+ cjswd = 5.1e-11
+ a0 = 1.4508547
+ a1 = 0
+ a2 = 1
+ cjsws = 5.1e-11
+ b0 = 0
+ b1 = 0
+ mjswd = 0.01
+ at = 72000
+ cf = 8.17e-11
+ mjsws = 0.01
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.013949949
+ k3 = -2.5823
+ agidl = 3.2166e-9
+ em = 20000000.0
+ ll = -1.18e-13
+ lw = 0
+ u0 = 0.0092421197
+ w0 = 0
+ ua = -3.1871506e-10
+ ub = 1.6925299e-18
+ uc = 2.1642376e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 6e-9
+ ags = 2.6576055
+ njtsswg = 6.489
+ mjswgd = 0.95
+ mjswgs = 0.95
+ cjd = 0.001346
+ cit = 0.00044006838
+ cjs = 0.001346
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ rshg = 14.1
+ bvs = 8.2
+ dlc = 1.38228675e-8
+ xtsswgd = 0.32
+ k3b = 2.1176
+ xtsswgs = 0.32
+ tcjswg = 0.00128
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.016932267
+ pdiblcb = 0
+ la0 = -4.2380342e-8
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0
+ kt1 = -0.23958332
+ kt2 = -0.07162235
+ lk2 = 4.3055939e-9
+ scref = 1e-6
+ llc = -1.18e-13
+ lln = 0.7
+ lu0 = -1.8443925e-10
+ mjd = 0.335
+ mjs = 0.335
+ lua = -2.581899e-17
+ lub = -2.6275812e-26
+ luc = -1.1293514e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ pigcd = 2.572
+ njd = 1.02
+ njs = 1.02
+ aigsd = 0.0063636407
+ pa0 = 0
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ pk2 = 0
+ pu0 = 0
+ prt = 0
+ pud = 0
+ tnom = 25
+ lvoff = -1.3382853e-9
+ rsh = 15.2
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ tcj = 0.000832
+ ua1 = 2.2510566e-9
+ ub1 = -2.8588123e-18
+ uc1 = 7.8974359e-11
+ bigbacc = 0.0054401
+ tpb = 0.0016
+ lvsat = 0.00084760684
+ ijthsfwd = 0.01
+ wa0 = 0
+ ute = -1
+ lvth0 = 5.1777832e-9
+ web = 6628.3
+ wec = -16935.0
+ fprout = 200
+ wk2 = 0
+ wlc = 0
+ wln = 1
+ wu0 = 0
+ xgl = -8.2e-9
+ xgw = 0
+ delta = 0.018814
+ wud = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ laigc = -2.0986759e-11
+ kvth0we = -0.00022
+ rnoia = 0
+ rnoib = 0
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ wtvoff = 0
+ vtsswgs = 1.1
+ ijthsrev = 0.01
+ ngate = 1.7e+20
+ wcit = 0.0
+ ngcon = 1
+ wpclm = 0
+ voff = -0.13301586
+ acde = 0.5
+ gbmin = 1e-12
+ capmod = 2
+ vsat = 115982.91
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ wint = 0
+ vth0 = -0.40736548
+ wku0we = 1.5e-11
+ wmax = 0.00090001
+ aigc = 0.0067688324
+ wmin = 9e-6
+ mobmod = 0
+ ppdiblc2 = 0
+ bigc = 0.0012521
+ wwlc = 0
+ nfactor = 1
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ tvoff = 0.0018930751
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigc = 0.15259
+ xjbvd = 1
+ xjbvs = 1
+ pkvth0we = 0.0
+ lk2we = 0.0
+ vfbsdoff = 0.01
+ ku0we = -0.0007
+ nigbacc = 10
+ beta0 = 13.32
+ leta0 = 0
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ ppclm = 0
+ paramchk = 1
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ nigbinv = 2.171
+ k2we = 5e-5
+ tvfbsdoff = 0.1
+ dsub = 0.5
+ dtox = 3.91e-10
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ eta0 = 0.1672
+ ijthdfwd = 0.01
+ etab = -0.23
+ toxref = 3e-9
+ fnoimod = 1
+ eigbinv = 1.1
+ bigsd = 0.0003327
+ ijthdrev = 0.01
+ wvfbsdoff = 0
+ wvoff = 0
+ lvfbsdoff = 0
+ ltvoff = -6.6370123e-11
+ lpdiblc2 = -1.4976331e-9
+ wvsat = 0.0
+ wvth0 = 0.0
+ cigbacc = 0.245
+ lku0we = 1.8e-11
+ lketa = 1.1808374e-9
+ tnoimod = 0
+ epsrox = 3.9
+ xpart = 1
+ rdsmod = 0
+ cigbinv = 0.006
+ egidl = 0.001
+ lkvth0we = 3e-12
+ igbmod = 1
+ )

.model pch_tt_6 pmos (
+ level = 54
+ wpclm = 0
+ vfbsdoff = 0.01
+ rshg = 14.1
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ nfactor = 1
+ wtvfbsdoff = 0
+ paramchk = 1
+ permod = 1
+ ltvfbsdoff = 0
+ tnom = 25
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ nigbacc = 10
+ ijthdfwd = 0.01
+ voffcv = -0.125
+ wpemod = 1
+ tvoff = 0.00091084129
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ nigbinv = 2.171
+ ptvfbsdoff = 0
+ ijthdrev = 0.01
+ wcit = 0.0
+ ku0we = -0.0007
+ lpdiblc2 = 0
+ voff = -0.11896044
+ beta0 = 13.32
+ acde = 0.5
+ leta0 = -1.1141465e-9
+ letab = 2.0255694e-8
+ vsat = 185878.73
+ wint = 0
+ vth0 = -0.33730292
+ ppclm = 0
+ tpbswg = 0.001
+ wmax = 0.00090001
+ fnoimod = 1
+ aigc = 0.0067067782
+ wmin = 9e-6
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ eigbinv = 1.1
+ tvfbsdoff = 0.1
+ ptvoff = 0
+ lkvth0we = 3e-12
+ bigc = 0.0012521
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ wwlc = 0
+ diomod = 1
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ acnqsmod = 0
+ pditsd = 0
+ pditsl = 0
+ cgsl = 3.0105e-11
+ cjswgd = 1.81e-10
+ pku0we = 0.0
+ cgso = 2.6482e-11
+ cigbacc = 0.245
+ cjswgs = 1.81e-10
+ cigc = 0.15259
+ bigsd = 0.0003327
+ rbodymod = 0
+ wvfbsdoff = 0
+ tnoimod = 0
+ lvfbsdoff = 0
+ wvoff = 0
+ mjswgd = 0.95
+ mjswgs = 0.95
+ wvsat = 0.0
+ cigbinv = 0.006
+ wvth0 = 0.0
+ tcjswg = 0.00128
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ version = 4.5
+ lketa = 8.4925319e-9
+ k2we = 5e-5
+ tempmod = 0
+ wpdiblc2 = 0
+ xpart = 1
+ dsub = 0.5
+ dtox = 3.91e-10
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ egidl = 0.001
+ a0 = 3.4166667
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 140456.11
+ cf = 8.17e-11
+ aigbacc = 0.012071
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.010241786
+ k3 = -2.5823
+ em = 20000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.0052338889
+ w0 = 0
+ ua = -1.1682959e-9
+ ub = 1.3034444e-18
+ uc = -8.7638e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 6e-9
+ fprout = 200
+ eta0 = 0.17905262
+ etab = -0.44548611
+ xrcrg1 = 12
+ xrcrg2 = 1
+ aigbinv = 0.009974
+ wkvth0we = 0.0
+ wtvoff = 0
+ trnqsmod = 0
+ capmod = 2
+ pvoff = 0
+ wku0we = 1.5e-11
+ cdscb = 0
+ cdscd = 0
+ mobmod = 0
+ pvsat = 0.0
+ wk2we = 0.0
+ pvth0 = 0.0
+ drout = 0.56
+ poxedge = 1
+ rgatemod = 0
+ voffl = 0
+ tnjtsswg = 1
+ binunit = 2
+ weta0 = 0
+ lpclm = -9.8438889e-8
+ cgidl = 1
+ keta = -0.20642296
+ pbswd = 0.9
+ pbsws = 0.9
+ lags = -2.8753242e-8
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ lcit = 1.8551944e-10
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ kt1l = 0
+ pdits = 0
+ cigsd = 0.013281
+ lint = 0
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ lkt1 = -1.23119e-9
+ lkt2 = 1.5220167e-10
+ lmax = 9e-8
+ lmin = 5.4e-8
+ lpe0 = 6.44e-8
+ lpeb = 0
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ minv = -0.33
+ lua1 = -7.3062676e-18
+ lub1 = 1.0038041e-26
+ luc1 = 7.6176556e-18
+ ndep = 1e+18
+ toxref = 3e-9
+ njtsswg = 6.489
+ tnoia = 0
+ ijthsfwd = 0.01
+ lwlc = 0
+ pvfbsdoff = 0
+ moin = 5.5538
+ xtsswgd = 0.32
+ peta0 = 0
+ xtsswgs = 0.32
+ nigc = 2.291
+ ckappad = 0.6
+ ckappas = 0.6
+ tpbsw = 0.0025
+ ags = 3.3058856
+ pdiblc1 = 0
+ pdiblc2 = 0.001
+ pdiblcb = 0
+ cjswd = 5.1e-11
+ cjd = 0.001346
+ cjsws = 5.1e-11
+ cit = -0.00072561111
+ cjs = 0.001346
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ dlc = 4.0349e-9
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ k3b = 2.1176
+ ijthsrev = 0.01
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ ltvoff = 2.5959859e-11
+ la0 = -2.2716667e-7
+ ntox = 1
+ pcit = 0.0
+ jsd = 1.5e-7
+ pclm = 2.4472222
+ jss = 1.5e-7
+ lat = -0.0064348744
+ kt1 = -0.27692169
+ kt2 = -0.078859167
+ lk2 = 3.9570266e-9
+ llc = 0
+ lln = 1
+ lu0 = 1.9233444e-10
+ mjd = 0.335
+ bigbacc = 0.0054401
+ mjs = 0.335
+ lua = 5.4041604e-17
+ lub = 1.0298222e-26
+ luc = 9.143004e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 0
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ pk2 = 0
+ phin = 0.15
+ pu0 = 0
+ lku0we = 1.8e-11
+ prt = 0
+ pub = 0.0
+ pud = 0
+ kvth0we = -0.00022
+ epsrox = 3.9
+ ppdiblc2 = 0
+ rsh = 15.2
+ scref = 1e-6
+ pkt1 = 0
+ tcj = 0.000832
+ ua1 = 7.2751825e-10
+ ub1 = -1.1117937e-18
+ uc1 = 7.4761111e-11
+ tpb = 0.0016
+ pigcd = 2.572
+ lintnoi = -5e-9
+ wa0 = 0
+ aigsd = 0.0063636407
+ ute = -1
+ web = 6628.3
+ wec = -16935.0
+ bigbinv = 0.00149
+ wk2 = 0
+ rdsmod = 0
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ wlc = 0
+ wln = 1
+ wu0 = 0
+ xgl = -8.2e-9
+ xgw = 0
+ wub = 0.0
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ igbmod = 1
+ lvoff = -2.6594942e-9
+ rbdb = 50
+ prwb = 0
+ prwg = 0
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ rbpb = 50
+ rbpd = 50
+ lvsat = -0.0057226009
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ lvth0 = -1.408097e-9
+ pbswgd = 0.8
+ pbswgs = 0.8
+ rdsw = 200
+ delta = 0.018814
+ laigc = -1.5153664e-11
+ igcmod = 1
+ rnoia = 0
+ rnoib = 0
+ pkvth0we = 0.0
+ ngate = 1.7e+20
+ ngcon = 1
+ )

.model pch_tt_7 pmos (
+ level = 54
+ voffl = 0
+ dsub = 0.5
+ dtox = 3.91e-10
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ weta0 = 0
+ ptvfbsdoff = 0
+ lpclm = -4.4240467e-8
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ eta0 = 0.18948293
+ ijthsfwd = 0.01
+ voffcv = -0.125
+ wpemod = 1
+ etab = -0.27185615
+ cgidl = 1
+ ijthsrev = 0.01
+ pbswd = 0.9
+ pbsws = 0.9
+ njtsswg = 6.489
+ tpbswg = 0.001
+ pdits = 0
+ cigsd = 0.013281
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ ppdiblc2 = 0
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.001
+ pdiblcb = 0
+ pk2we = 0.0
+ ptvoff = 0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ ags = 2.81014
+ pvfbsdoff = 0
+ tnoia = 0
+ diomod = 1
+ cjd = 0.001346
+ cit = -0.0030912222
+ cjs = 0.001346
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 4.0349e-9
+ peta0 = 0
+ k3b = 2.1176
+ pditsd = 0
+ pditsl = 0
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ bigbacc = 0.0054401
+ dwj = 0
+ cjswgd = 1.81e-10
+ pku0we = 0.0
+ cjswgs = 1.81e-10
+ tpbsw = 0.0025
+ pkvth0we = 0.0
+ keta = 0.048888889
+ cjswd = 5.1e-11
+ kvth0we = -0.00022
+ cjsws = 5.1e-11
+ la0 = -1.5788889e-7
+ jsd = 1.5e-7
+ mjswd = 0.01
+ jss = 1.5e-7
+ lat = 0.0042661578
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ kt1 = -0.090229195
+ kt2 = -0.087042222
+ lk2 = 4.3353879e-9
+ llc = 0
+ lln = 1
+ lu0 = -7.2628889e-11
+ mjd = 0.335
+ mjs = 0.335
+ lua = -4.5270917e-17
+ lub = -1.9748742e-26
+ luc = -2.161341e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ lintnoi = -5e-9
+ njd = 1.02
+ mjswgd = 0.95
+ njs = 1.02
+ mjswgs = 0.95
+ pa0 = 0
+ bigbinv = 0.00149
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ jswd = 3.69e-13
+ vtsswgd = 1.1
+ pk2 = 0
+ jsws = 3.69e-13
+ vtsswgs = 1.1
+ vfbsdoff = 0.01
+ lcit = 3.2272489e-10
+ pu0 = 0
+ tcjswg = 0.00128
+ prt = 0
+ pub = 0.0
+ pud = 0
+ kt1l = 0
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 1.0031266e-9
+ ub1 = -2.5489021e-18
+ uc1 = 1.9738889e-10
+ tpb = 0.0016
+ wa0 = 0
+ ute = -1
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 0
+ lint = 0
+ wlc = 0
+ wln = 1
+ wu0 = 0
+ xgl = -8.2e-9
+ xgw = 0
+ paramchk = 1
+ wub = 0.0
+ wud = 0
+ wwc = 0
+ lkt1 = -1.2059355e-8
+ lkt2 = 6.2681889e-10
+ wwl = 0
+ wwn = 1
+ lmax = 5.4e-8
+ lmin = 4.5e-8
+ scref = 1e-6
+ lpe0 = 6.44e-8
+ lpeb = 0
+ pigcd = 2.572
+ aigsd = 0.0063636407
+ minv = -0.33
+ lvoff = -4.1866651e-9
+ lua1 = -2.3291554e-17
+ lub1 = 9.339033e-26
+ luc1 = 5.0524444e-19
+ fprout = 200
+ ndep = 1e+18
+ lvsat = -0.00014010428
+ ijthdfwd = 0.01
+ xrcrg1 = 12
+ xrcrg2 = 1
+ lwlc = 0
+ lvth0 = -2.3166339e-9
+ moin = 5.5538
+ delta = 0.018814
+ laigc = -9.9932362e-12
+ nigc = 2.291
+ nfactor = 1
+ rnoia = 0
+ rnoib = 0
+ wtvoff = 0
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ ijthdrev = 0.01
+ ngate = 1.7e+20
+ ngcon = 1
+ wpclm = 0
+ lpdiblc2 = 0
+ capmod = 2
+ ntox = 1
+ pcit = 0.0
+ wku0we = 1.5e-11
+ pclm = 1.5127667
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ nigbacc = 10
+ a0 = 2.2222222
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = -44044.444
+ mobmod = 0
+ cf = 8.17e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.016765256
+ k3 = -2.5823
+ em = 20000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.0098022222
+ w0 = 0
+ ua = 5.4398899e-10
+ ub = 1.8214956e-18
+ uc = 4.42645e-10
+ ud = 0
+ phin = 0.15
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 6e-9
+ pkt1 = 0
+ nigbinv = 2.171
+ lkvth0we = 3e-12
+ rbdb = 50
+ prwb = 0
+ prwg = 0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ rdsw = 200
+ tvoff = 0.0051729841
+ acnqsmod = 0
+ fnoimod = 1
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ eigbinv = 1.1
+ rbodymod = 0
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = -1.7191043e-9
+ rshg = 14.1
+ letab = 1.0185157e-8
+ ppclm = 0
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ tvfbsdoff = 0.1
+ cigbacc = 0.245
+ wpdiblc2 = 0
+ tnoimod = 0
+ tnom = 25
+ dmcgt = 0
+ toxref = 3e-9
+ tcjsw = 9.34e-5
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ cigbinv = 0.006
+ bigsd = 0.0003327
+ wkvth0we = 0.0
+ version = 4.5
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ tempmod = 0
+ ltvoff = -2.2124443e-10
+ wvoff = 0
+ wcit = 0.0
+ trnqsmod = 0
+ voff = -0.092629909
+ wvsat = 0.0
+ acde = 0.5
+ wvth0 = 0.0
+ aigbacc = 0.012071
+ vsat = 89628.791
+ wint = 0
+ vth0 = -0.32163849
+ lku0we = 1.8e-11
+ wmax = 0.00090001
+ aigc = 0.0066178053
+ wmin = 9e-6
+ epsrox = 3.9
+ lketa = -6.3155556e-9
+ rgatemod = 0
+ xpart = 1
+ aigbinv = 0.009974
+ tnjtsswg = 1
+ rdsmod = 0
+ igbmod = 1
+ egidl = 0.001
+ bigc = 0.0012521
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ wwlc = 0
+ pbswgd = 0.8
+ pbswgs = 0.8
+ cdsc = 0
+ cgbo = 0
+ igcmod = 1
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigc = 0.15259
+ wtvfbsdoff = 0
+ poxedge = 1
+ binunit = 2
+ ltvfbsdoff = 0
+ pvoff = 0
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ cdscb = 0
+ cdscd = 0
+ pvsat = 0.0
+ wk2we = 0.0
+ pvth0 = 0.0
+ drout = 0.56
+ permod = 1
+ k2we = 5e-5
+ )

.model pch_tt_8 pmos (
+ level = 54
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ wkvth0we = 0.0
+ cigbacc = 0.245
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ trnqsmod = 0
+ ku0we = -0.0007
+ tnoimod = 0
+ beta0 = 13.32
+ leta0 = 2.1323128e-9
+ ntox = 1
+ letab = 3.9337702e-9
+ pcit = 0.0
+ pclm = 1.0208333
+ tpbswg = 0.001
+ cigbinv = 0.006
+ ppclm = 0
+ phin = 0.15
+ dlcig = 2.5e-9
+ tvfbsdoff = 0.1
+ bgidl = 1834800000.0
+ pkt1 = 0.0
+ rgatemod = 0
+ ptvoff = 0
+ tnjtsswg = 1
+ version = 4.5
+ tempmod = 0
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ diomod = 1
+ rbdb = 50
+ prwb = 0
+ prwg = 0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ aigbacc = 0.012071
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.81e-10
+ pku0we = 0.0
+ cjswgs = 1.81e-10
+ rdsw = 200
+ bigsd = 0.0003327
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ mjswgd = 0.95
+ mjswgs = 0.95
+ wvoff = 0
+ aigbinv = 0.009974
+ tcjswg = 0.00128
+ wvsat = 0.0
+ wvth0 = 0.0
+ rshg = 14.1
+ lketa = 8.0381778e-9
+ xpart = 1
+ poxedge = 1
+ egidl = 0.001
+ tnom = 25
+ fprout = 200
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ xrcrg1 = 12
+ xrcrg2 = 1
+ binunit = 2
+ ijthsfwd = 0.01
+ wtvoff = 0
+ ijthsrev = 0.01
+ wcit = 0.0
+ capmod = 2
+ voff = -0.10032114
+ wku0we = 1.5e-11
+ acde = 0.5
+ pvoff = 0
+ mobmod = 0
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ vsat = 122520.32
+ wint = 0
+ vth0 = -0.36838557
+ cdscb = 0
+ cdscd = 0
+ wkt1 = 0.0
+ pvsat = 0.0
+ wmax = 0.00090001
+ wk2we = 0.0
+ pvth0 = 0.0
+ aigc = 0.0065563017
+ wmin = 9e-6
+ drout = 0.56
+ ppdiblc2 = 0
+ voffl = 0
+ weta0 = 0
+ wetab = 0
+ bigc = 0.0012521
+ wwlc = 0
+ lpclm = -2.0135733e-8
+ laigsd = -2.1777787e-18
+ cdsc = 0
+ cgidl = 1
+ njtsswg = 6.489
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigc = 0.15259
+ a0 = -0.19555556
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ xtsswgd = 0.32
+ pkvth0we = 0.0
+ xtsswgs = 0.32
+ at = 76220.0
+ cf = 8.17e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.012217534
+ k3 = -2.5823
+ em = 20000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.0052977778
+ w0 = 0
+ ua = -1.1794951e-9
+ ub = 1.5005044e-18
+ uc = 5.0701667e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 6e-9
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.001
+ pbswd = 0.9
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ pbsws = 0.9
+ pdiblcb = 0
+ vfbsdoff = 0.01
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ pdits = 0
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ paramchk = 1
+ bigbacc = 0.0054401
+ k2we = 5e-5
+ ags = 1.0774289
+ dsub = 0.5
+ kvth0we = -0.00022
+ dtox = 3.91e-10
+ cjd = 0.001346
+ cit = -0.00097166667
+ pk2we = 0.0
+ cjs = 0.001346
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ dlc = 4.0349e-9
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ k3b = 2.1176
+ toxref = 3e-9
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ pvfbsdoff = 0
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ tnoia = 0
+ ijthdfwd = 0.01
+ eta0 = 0.11088258
+ etab = -0.14427684
+ la0 = -3.9417778e-8
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = -0.0016268
+ kt1 = -0.30391077
+ kt2 = -0.08425
+ lk2 = 4.1125495e-9
+ peta0 = 0
+ llc = 0
+ lln = 1
+ lu0 = 1.4808889e-10
+ petab = 0
+ mjd = 0.335
+ mjs = 0.335
+ lua = 3.9179804e-17
+ lub = -4.0201778e-27
+ luc = -2.4081867e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 0
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0.0
+ pbs = 0.75
+ tpbsw = 0.0025
+ pk2 = 0
+ pu0 = 0
+ prt = 0
+ pub = 0.0
+ pud = 0
+ cjswd = 5.1e-11
+ cjsws = 5.1e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ ltvoff = -2.4936809e-11
+ agidl = 3.2166e-9
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 1.4917512e-9
+ ub1 = -1.5908843e-18
+ uc1 = 1.6325556e-10
+ ijthdrev = 0.01
+ tpb = 0.0016
+ wa0 = 0
+ ute = -1
+ wat = 0.0
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 0
+ wlc = 0
+ wln = 1
+ lpdiblc2 = 0
+ wu0 = 0
+ xgl = -8.2e-9
+ xgw = 0
+ wub = 0.0
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ lku0we = 1.8e-11
+ epsrox = 3.9
+ nfactor = 1
+ scref = 1e-6
+ rdsmod = 0
+ pigcd = 2.572
+ aigsd = 0.0063636407
+ igbmod = 1
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ wtvfbsdoff = 0
+ lvoff = -3.8097951e-9
+ lkvth0we = 3e-12
+ pbswgd = 0.8
+ pbswgs = 0.8
+ lvsat = -0.0017517894
+ lvth0 = -2.6027058e-11
+ igcmod = 1
+ ltvfbsdoff = 0
+ delta = 0.018814
+ nigbacc = 10
+ laigc = -6.97956e-12
+ acnqsmod = 0
+ rnoia = 0
+ rnoib = 0
+ keta = -0.24404444
+ rbodymod = 0
+ ngate = 1.7e+20
+ lags = 8.4902844e-8
+ ngcon = 1
+ nigbinv = 2.171
+ wpclm = 0
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 2.1886667e-10
+ kt1l = 0
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ ptvfbsdoff = 0
+ lint = 0
+ permod = 1
+ lkt1 = -1.5889574e-9
+ lkt2 = 4.9e-10
+ lmax = 4.5e-8
+ lmin = 3.6e-8
+ fnoimod = 1
+ wpdiblc2 = 0
+ lpe0 = 6.44e-8
+ lpeb = 0
+ eigbinv = 1.1
+ minv = -0.33
+ lua1 = -4.7234158e-17
+ lub1 = 4.6447457e-26
+ luc1 = 2.1777778e-18
+ voffcv = -0.125
+ wpemod = 1
+ ndep = 1e+18
+ lwlc = 0
+ moin = 5.5538
+ tvoff = 0.0011667062
+ nigc = 2.291
+ )

.model pch_tt_9 pmos (
+ level = 54
+ vtsswgs = 1.1
+ ags = 0.82538676
+ vsat = 121084.96
+ wint = 0
+ vth0 = -0.38547733
+ pdits = 0
+ cjd = 0.001346
+ cit = 5e-6
+ cjs = 0.001346
+ clc = 1e-7
+ cle = 0.6
+ cigsd = 0.013281
+ bvd = 8.2
+ bvs = 8.2
+ wkt1 = -1.0361455e-8
+ wkt2 = -3.8769913e-9
+ dlc = 1.0572421799999999e-8
+ wmax = 9e-6
+ dvt0w = 0
+ k3b = 2.1176
+ dvt1w = 0
+ aigc = 0.0068303602
+ dvt2w = 0
+ wmin = 9e-7
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ ptvoff = 0
+ waigsd = 1.9139418e-12
+ la0 = 0
+ pk2we = 0.0
+ jsd = 1.5e-7
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ jss = 1.5e-7
+ lat = 0
+ wua1 = -3.2799159e-16
+ kt1 = -0.16992583
+ lk2 = 0
+ kt2 = -0.04703951
+ wub1 = 5.9231251e-25
+ wuc1 = -8.7396626e-17
+ llc = 0
+ lln = 1
+ lu0 = 0
+ mjd = 0.335
+ mjs = 0.335
+ lkvth0we = 3e-12
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ diomod = 1
+ pvfbsdoff = 0
+ njd = 1.02
+ bigc = 0.0012521
+ njs = 1.02
+ wute = -7.8572347e-8
+ pa0 = 0
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ wwlc = 0
+ pk2 = 0
+ tnoia = 0
+ pu0 = 0
+ pditsd = 0
+ pditsl = 0
+ prt = 0
+ pud = 0
+ cjswgd = 1.81e-10
+ pku0we = 0.0
+ cjswgs = 1.81e-10
+ rsh = 15.2
+ tcj = 0.000832
+ peta0 = 0
+ cdsc = 0
+ ua1 = 1.2333536e-9
+ ub1 = -1.432383e-18
+ uc1 = 7.8434267e-11
+ cgbo = 0
+ tpb = 0.0016
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ acnqsmod = 0
+ xtid = 3
+ xtis = 3
+ wketa = 2.2362589e-8
+ wa0 = 3.3745816e-7
+ ute = -0.99127556
+ web = 6628.3
+ wec = -16935.0
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ wk2 = -2.287053e-9
+ tpbsw = 0.0025
+ cigc = 0.15259
+ wlc = 0
+ wln = 1
+ wu0 = -8.6631049e-11
+ xgl = -8.2e-9
+ xgw = 0
+ wua = -1.124189e-16
+ wub = -6.7100784e-26
+ wuc = -2.319496e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ cjswd = 5.1e-11
+ nfactor = 1
+ cjsws = 5.1e-11
+ mjswd = 0.01
+ mjswgd = 0.95
+ mjsws = 0.01
+ mjswgs = 0.95
+ agidl = 3.2166e-9
+ rbodymod = 0
+ tcjswg = 0.00128
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ nigbacc = 10
+ scref = 1e-6
+ k2we = 5e-5
+ wpdiblc2 = 3.6469361e-10
+ pigcd = 2.572
+ dsub = 0.5
+ aigsd = 0.0063633875
+ dtox = 3.91e-10
+ fprout = 200
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ lvoff = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ nigbinv = 2.171
+ lvsat = 0
+ eta0 = 0.16744607
+ etab = -0.23671111
+ lvth0 = 0.0
+ delta = 0.018814
+ wtvoff = -9.8925647e-11
+ rnoia = 0
+ rnoib = 0
+ wkvth0we = 0.0
+ fnoimod = 1
+ ngate = 1.7e+20
+ capmod = 2
+ trnqsmod = 0
+ eigbinv = 1.1
+ ngcon = 1
+ wpclm = -3.01194e-7
+ wku0we = 1.5e-11
+ mobmod = 0
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ rgatemod = 0
+ tnjtsswg = 1
+ cigbacc = 0.245
+ tnoimod = 0
+ tvoff = 0.0026265487
+ cigbinv = 0.006
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ keta = -0.044833188
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ version = 4.5
+ jswd = 3.69e-13
+ ku0we = -0.0007
+ jsws = 3.69e-13
+ lcit = 0
+ tempmod = 0
+ beta0 = 13.32
+ leta0 = 0
+ kt1l = 0
+ ppclm = 0
+ aigbacc = 0.012071
+ lint = 6.5375218e-9
+ tvfbsdoff = 0.1
+ dlcig = 2.5e-9
+ lkt1 = 0
+ bgidl = 1834800000.0
+ lmax = 2.001e-5
+ lmin = 8.9991e-6
+ lpe0 = 6.44e-8
+ lpeb = 0
+ a0 = 2.4935296
+ a1 = 0
+ a2 = 1
+ toxref = 3e-9
+ b0 = 0
+ b1 = 0
+ at = 72000
+ cf = 8.17e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.00052197993
+ k3 = -2.5823
+ em = 20000000.0
+ aigbinv = 0.009974
+ minv = -0.33
+ ll = 0
+ lw = 0
+ u0 = 0.0098046193
+ w0 = 0
+ ua = 1.4218267e-10
+ ub = 1.1900227e-18
+ uc = 2.2715501e-11
+ ud = 0
+ dmcgt = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 6e-9
+ tcjsw = 9.34e-5
+ ndep = 1e+18
+ ijthsfwd = 0.01
+ lwlc = 0
+ moin = 5.5538
+ nigc = 2.291
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ bigsd = 0.0003327
+ ltvoff = 0
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ ijthsrev = 0.01
+ wvoff = 5.5905393e-9
+ poxedge = 1
+ wvsat = -0.0097711764
+ wvth0 = 3.080586e-9
+ ntox = 1
+ pcit = 0
+ pclm = 1.5174437
+ binunit = 2
+ lku0we = 1.8e-11
+ wtvfbsdoff = 0
+ waigc = 3.5172206e-12
+ epsrox = 3.9
+ phin = 0.15
+ lketa = 0
+ rdsmod = 0
+ ltvfbsdoff = 0
+ ppdiblc2 = 0
+ pkt1 = 0
+ xpart = 1
+ igbmod = 1
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ egidl = 0.001
+ pbswgd = 0.8
+ pbswgs = 0.8
+ rbdb = 50
+ prwb = 0
+ prwg = 0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ igcmod = 1
+ rbsb = 50
+ pvag = 2.1
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ rdsw = 200
+ ptvfbsdoff = 0
+ pkvth0we = 0.0
+ vfbsdoff = 0.01
+ rshg = 14.1
+ pvoff = 0
+ cdscb = 0
+ cdscd = 0
+ permod = 1
+ pvsat = 0
+ wk2we = 0.0
+ pvth0 = 0.0
+ paramchk = 1
+ njtsswg = 6.489
+ drout = 0.56
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ voffl = 0
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.0026324684
+ weta0 = -2.2161431e-9
+ tnom = 25
+ pdiblcb = 0
+ wetab = 6.0440267e-8
+ voffcv = -0.125
+ wpemod = 1
+ lpclm = 0
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ ijthdfwd = 0.01
+ cgidl = 1
+ bigbacc = 0.0054401
+ wags = 1.128996e-7
+ ijthdrev = 0.01
+ pbswd = 0.9
+ pbsws = 0.9
+ kvth0we = -0.00022
+ lpdiblc2 = 0
+ voff = -0.11172412
+ tpbswg = 0.001
+ acde = 0.5
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ )

.model pch_tt_10 pmos (
+ level = 54
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ lags = 3.1017116e-7
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 0
+ nfactor = 1
+ kt1l = 0
+ paramchk = 1
+ scref = 1e-6
+ pigcd = 2.572
+ aigsd = 0.0063633879
+ lint = 6.5375218e-9
+ lkt1 = -4.1907452e-8
+ lkt2 = -8.3161855e-9
+ lmax = 8.9991e-6
+ lvoff = -7.1040424e-9
+ lmin = 8.9908e-7
+ lpe0 = 6.44e-8
+ lpeb = 0
+ lvsat = 0
+ lvth0 = -4.4817588e-9
+ ijthdfwd = 0.01
+ toxref = 3e-9
+ nigbacc = 10
+ minv = -0.33
+ delta = 0.018814
+ lua1 = 2.9697696e-17
+ lub1 = 1.2607181e-25
+ luc1 = -4.744495e-18
+ laigc = -4.752933e-11
+ wtvfbsdoff = 0
+ ndep = 1e+18
+ rnoia = 0
+ rnoib = 0
+ lute = -8.6179201e-9
+ lwlc = 0
+ tvfbsdoff = 0.1
+ moin = 5.5538
+ ltvfbsdoff = 0
+ pketa = -2.2807538e-14
+ nigc = 2.291
+ ngate = 1.7e+20
+ ijthdrev = 0.01
+ nigbinv = 2.171
+ ngcon = 1
+ wpclm = -3.01194e-7
+ lpdiblc2 = 7.3300428e-9
+ ltvoff = -4.2514859e-10
+ gbmin = 1e-12
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ pags = -3.4942959e-14
+ ntox = 1
+ pcit = 0
+ pclm = 1.5174437
+ fnoimod = 1
+ wvfbsdoff = 0
+ lku0we = 1.8e-11
+ ptvfbsdoff = 0
+ eigbinv = 1.1
+ lvfbsdoff = 0
+ epsrox = 3.9
+ phin = 0.15
+ lkvth0we = 3e-12
+ pkt1 = 9.0189586e-15
+ pkt2 = -4.3236504e-15
+ rdsmod = 0
+ igbmod = 1
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ tvoff = 0.0026738399
+ pbswgd = 0.8
+ acnqsmod = 0
+ pbswgs = 0.8
+ rbdb = 50
+ pua1 = 9.6044121e-22
+ prwb = 0
+ pub1 = -1.3952204e-30
+ prwg = 0
+ puc1 = 1.1914589e-22
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ pute = 7.7612988e-14
+ igcmod = 1
+ cigbacc = 0.245
+ rdsw = 200
+ rbodymod = 0
+ tnoimod = 0
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = 0
+ cigbinv = 0.006
+ ppclm = 0
+ paigsd = 3.3403436e-20
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ rshg = 14.1
+ version = 4.5
+ wpdiblc2 = 5.6393415e-10
+ permod = 1
+ tempmod = 0
+ ags = 0.79088496
+ dmcgt = 0
+ cjd = 0.001346
+ cit = 5e-6
+ cjs = 0.001346
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ tcjsw = 9.34e-5
+ dlc = 1.0572421799999999e-8
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ aigbacc = 0.012071
+ tnom = 25
+ la0 = -3.6651331e-7
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ jsd = 1.5e-7
+ voffcv = -0.125
+ wpemod = 1
+ jss = 1.5e-7
+ lat = 0
+ kt1 = -0.16526426
+ kt2 = -0.046114462
+ lk2 = 4.5045048e-9
+ llc = 0
+ lln = 1
+ bigsd = 0.0003327
+ lu0 = -1.1944212e-10
+ mjd = 0.335
+ mjs = 0.335
+ lua = -1.1601528e-16
+ lub = 1.1870612e-25
+ luc = 1.7407612e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = -2.3980423e-13
+ wkvth0we = 0.0
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ pk2 = -1.7678537e-15
+ aigbinv = 0.009974
+ wvoff = 6.4925381e-9
+ pu0 = 1.0845918e-15
+ prt = 0
+ pua = 1.4359661e-22
+ pub = 1.4495718e-31
+ puc = -1.3724663e-23
+ pud = 0
+ trnqsmod = 0
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 1.2300502e-9
+ ub1 = -1.4464065e-18
+ uc1 = 7.8962019e-11
+ wvsat = -0.0097711764
+ tpb = 0.0016
+ wvth0 = 3.7267412e-9
+ wa0 = 3.6413271e-7
+ ute = -0.99031694
+ wags = 1.1678647e-7
+ web = 6628.3
+ wec = -16935.0
+ wk2 = -2.0904063e-9
+ wlc = 0
+ wln = 1
+ wu0 = -2.0727529e-10
+ xgl = -8.2e-9
+ waigc = 4.3868453e-12
+ xgw = 0
+ wua = -1.2839182e-16
+ wub = -8.3225053e-26
+ wuc = -2.1668301e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ voff = -0.11093391
+ acde = 0.5
+ tpbswg = 0.001
+ lketa = -1.0921036e-8
+ vsat = 121084.96
+ wint = 0
+ xpart = 1
+ vth0 = -0.3849788
+ rgatemod = 0
+ wkt1 = -1.1364676e-8
+ wkt2 = -3.3960513e-9
+ poxedge = 1
+ wmax = 9e-6
+ tnjtsswg = 1
+ aigc = 0.0068356471
+ wmin = 9e-7
+ egidl = 0.001
+ binunit = 2
+ ptvoff = -4.5667618e-16
+ waigsd = 1.9102262e-12
+ wua1 = -4.3482598e-16
+ wub1 = 7.4750944e-25
+ wuc1 = -1.0064978e-16
+ bigc = 0.0012521
+ wute = -8.7205605e-8
+ diomod = 1
+ wwlc = 0
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.81e-10
+ pku0we = 0.0
+ cjswgs = 1.81e-10
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigc = 0.15259
+ pvoff = -8.1089692e-15
+ jtsswgd = 1.75e-7
+ pvfbsdoff = 0
+ mjswgd = 0.95
+ jtsswgs = 1.75e-7
+ mjswgs = 0.95
+ cdscb = 0
+ cdscd = 0
+ tcjswg = 0.00128
+ pvsat = 0
+ wk2we = 0.0
+ pvth0 = -5.8089351e-15
+ drout = 0.56
+ paigc = -7.8179264e-18
+ a0 = 2.5342986
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 72000
+ cf = 8.17e-11
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.0010230372
+ k3 = -2.5823
+ em = 20000000.0
+ voffl = 0
+ ll = 0
+ lw = 0
+ u0 = 0.0098179054
+ w0 = 0
+ ua = 1.5508759e-10
+ ub = 1.1768184e-18
+ uc = 2.077917e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 6e-9
+ weta0 = -2.2161431e-9
+ wetab = 6.0440267e-8
+ k2we = 5e-5
+ lpclm = 0
+ dsub = 0.5
+ dtox = 3.91e-10
+ ijthsfwd = 0.01
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ njtsswg = 6.489
+ cgidl = 1
+ fprout = 200
+ xrcrg1 = 12
+ xrcrg2 = 1
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ eta0 = 0.16744607
+ etab = -0.23671111
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.0018171133
+ pdiblcb = 0
+ pbswd = 0.9
+ wtvoff = -4.8127407e-11
+ pbsws = 0.9
+ ijthsrev = 0.01
+ pdits = 0
+ capmod = 2
+ cigsd = 0.013281
+ wku0we = 1.5e-11
+ bigbacc = 0.0054401
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ mobmod = 0
+ ppdiblc2 = -1.7911725e-15
+ kvth0we = -0.00022
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ tnoia = 0
+ peta0 = 0
+ wketa = 2.4899578e-8
+ laigsd = -3.7090202e-15
+ tpbsw = 0.0025
+ pkvth0we = 0.0
+ cjswd = 5.1e-11
+ cjsws = 5.1e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ keta = -0.04361839
+ vfbsdoff = 0.01
+ )

.model pch_tt_11 pmos (
+ level = 54
+ egidl = 0.001
+ ltvfbsdoff = 0
+ toxref = 3e-9
+ ijthsfwd = 0.01
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ tnom = 25
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ ijthsrev = 0.01
+ ptvfbsdoff = 0
+ ltvoff = -2.603747e-10
+ pvfbsdoff = 0
+ wags = -5.7105665e-9
+ pvoff = 6.0510934e-15
+ cdscb = 0
+ cdscd = 0
+ pvsat = 0
+ wk2we = 0.0
+ voff = -0.10782222
+ njtsswg = 6.489
+ pvth0 = 3.2463808e-15
+ drout = 0.56
+ acde = 0.5
+ paigc = 1.0166993e-17
+ lku0we = 1.8e-11
+ xtsswgd = 0.32
+ vsat = 121084.96
+ xtsswgs = 0.32
+ wint = 0
+ ppdiblc2 = 8.932051e-16
+ vth0 = -0.38647369
+ epsrox = 3.9
+ voffl = 0
+ wkt1 = 3.9882501e-9
+ wkt2 = -1.3862366e-8
+ ckappad = 0.6
+ wmax = 9e-6
+ ckappas = 0.6
+ aigc = 0.0068328167
+ wmin = 9e-7
+ pdiblc1 = 0
+ pdiblc2 = 0.0082016634
+ pdiblcb = 0
+ weta0 = -2.2161431e-9
+ rdsmod = 0
+ wetab = 6.0440267e-8
+ igbmod = 1
+ lpclm = 0
+ wua1 = 1.0350058e-15
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ wub1 = -1.41997e-24
+ wuc1 = 5.1522417e-17
+ cgidl = 1
+ pbswgd = 0.8
+ bigc = 0.0012521
+ pbswgs = 0.8
+ wwlc = 0
+ bigbacc = 0.0054401
+ igcmod = 1
+ pkvth0we = 0.0
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ pbswd = 0.9
+ pbsws = 0.9
+ kvth0we = -0.00022
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigc = 0.15259
+ vfbsdoff = 0.01
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ pdits = 0
+ cigsd = 0.013281
+ paigsd = -3.7089273e-20
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ paramchk = 1
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ permod = 1
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ k2we = 5e-5
+ tnoia = 0
+ dsub = 0.5
+ dtox = 3.91e-10
+ ijthdfwd = 0.01
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ peta0 = 0
+ voffcv = -0.125
+ wpemod = 1
+ wketa = -2.3248862e-8
+ tpbsw = 0.0025
+ eta0 = 0.16744607
+ nfactor = 1
+ etab = -0.23671111
+ cjswd = 5.1e-11
+ cjsws = 5.1e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ ijthdrev = 0.01
+ lpdiblc2 = 1.6477933e-9
+ nigbacc = 10
+ tpbswg = 0.001
+ scref = 1e-6
+ pigcd = 2.572
+ aigsd = 0.0063633394
+ lvoff = -9.8734428e-9
+ nigbinv = 2.171
+ ptvoff = 2.6240046e-16
+ lkvth0we = 3e-12
+ waigsd = 1.9894315e-12
+ lvsat = 0
+ lvth0 = -3.1513088e-9
+ delta = 0.018814
+ diomod = 1
+ laigc = -4.5010295e-11
+ acnqsmod = 0
+ rnoia = 0
+ rnoib = 0
+ tvfbsdoff = 0.1
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.81e-10
+ pku0we = 0.0
+ cjswgs = 1.81e-10
+ fnoimod = 1
+ pketa = 2.0044574e-14
+ rbodymod = 0
+ ngate = 1.7e+20
+ eigbinv = 1.1
+ ngcon = 1
+ wpclm = -3.01194e-7
+ keta = -0.035478054
+ mjswgd = 0.95
+ mjswgs = 0.95
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ tcjswg = 0.00128
+ lags = 2.7680102e-7
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 8.2671111e-11
+ kt1l = 0
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ wpdiblc2 = -2.4522204e-9
+ lint = 6.5375218e-9
+ cigbacc = 0.245
+ lkt1 = -1.4522155e-8
+ lkt2 = -7.1896716e-9
+ lmax = 8.9908e-7
+ lmin = 4.4908e-7
+ tnoimod = 0
+ lpe0 = 6.44e-8
+ lpeb = 0
+ fprout = 200
+ minv = -0.33
+ cigbinv = 0.006
+ lua1 = 8.7159171e-17
+ lub1 = -2.6689299e-25
+ luc1 = 2.9116076e-17
+ tvoff = 0.0024887007
+ xrcrg1 = 12
+ xrcrg2 = 1
+ ndep = 1e+18
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ lwlc = 0
+ moin = 5.5538
+ wkvth0we = 0.0
+ wtvoff = -8.5607868e-10
+ nigc = 2.291
+ version = 4.5
+ a0 = 2.8862723
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ trnqsmod = 0
+ at = 72000
+ cf = 8.17e-11
+ tempmod = 0
+ ef = 1.15
+ ku0we = -0.0007
+ k1 = 0.30425
+ k2 = 0.0046668319
+ k3 = -2.5823
+ em = 20000000.0
+ ll = 0
+ lw = 0
+ beta0 = 13.32
+ u0 = 0.0098044338
+ w0 = 0
+ ua = 8.4190146e-11
+ ub = 1.1838278e-18
+ uc = 4.9200634e-11
+ ud = 0
+ leta0 = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 6e-9
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ capmod = 2
+ ppclm = 0
+ aigbacc = 0.012071
+ wku0we = 1.5e-11
+ pags = 7.4079401e-14
+ ags = 0.8283795
+ dlcig = 2.5e-9
+ mobmod = 0
+ bgidl = 1834800000.0
+ ntox = 1
+ pcit = 0
+ pclm = 1.5174437
+ cjd = 0.001346
+ cit = -8.7888889e-5
+ cjs = 0.001346
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 1.0572421799999999e-8
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ rgatemod = 0
+ tnjtsswg = 1
+ phin = 0.15
+ aigbinv = 0.009974
+ dmcgt = 0
+ la0 = -6.797699e-7
+ pkt1 = -4.6451461e-15
+ jsd = 1.5e-7
+ pkt2 = 4.9913693e-15
+ tcjsw = 9.34e-5
+ jss = 1.5e-7
+ lat = 0
+ kt1 = -0.19603426
+ kt2 = -0.047380208
+ lk2 = -5.594787e-10
+ llc = 0
+ lln = 1
+ lu0 = -1.0745246e-10
+ mjd = 0.335
+ mjs = 0.335
+ lua = -5.2916554e-17
+ lub = 1.1246778e-25
+ luc = -7.8874906e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 4.0323955e-14
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ pk2 = 1.1838025e-15
+ pu0 = -8.8186737e-16
+ laigsd = 3.9492818e-14
+ prt = 0
+ pua = -2.1071339e-22
+ pub = -4.1382897e-32
+ puc = 1.6409308e-23
+ pud = 0
+ rbdb = 50
+ pua1 = -3.4770908e-22
+ prwb = 0
+ pub1 = 5.3383631e-31
+ prwg = 0
+ rsh = 15.2
+ puc1 = -1.6287371e-23
+ tcj = 0.000832
+ ua1 = 1.1654868e-9
+ ub1 = -1.004873e-18
+ uc1 = 4.0916434e-11
+ bigsd = 0.0003327
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ tpb = 0.0016
+ wa0 = 4.9381936e-8
+ ute = -1
+ web = 6628.3
+ wec = -16935.0
+ wk2 = -5.406874e-9
+ rdsw = 200
+ wlc = 0
+ wln = 1
+ wu0 = 2.0022293e-9
+ xgl = -8.2e-9
+ wvoff = -9.4176445e-9
+ xgw = 0
+ wua = 2.6970929e-16
+ wub = 1.2614582e-25
+ wuc = -5.5526695e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ poxedge = 1
+ wvsat = -0.0097711764
+ wvth0 = -6.4477711e-9
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ binunit = 2
+ waigc = -1.5820929e-11
+ rshg = 14.1
+ lketa = -1.8165935e-8
+ xpart = 1
+ wtvfbsdoff = 0
+ )

.model pch_tt_12 pmos (
+ level = 54
+ wkvth0we = 0.0
+ pketa = 2.9922765e-15
+ ngate = 1.7e+20
+ ngcon = 1
+ cigbacc = 0.245
+ ltvoff = -1.0992228e-10
+ wpclm = -3.01194e-7
+ trnqsmod = 0
+ gbmin = 1e-12
+ tnoimod = 0
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ cigbinv = 0.006
+ lku0we = 1.8e-11
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ epsrox = 3.9
+ rgatemod = 0
+ tnjtsswg = 1
+ rdsmod = 0
+ version = 4.5
+ igbmod = 1
+ tempmod = 0
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ pbswgd = 0.8
+ pbswgs = 0.8
+ tvoff = 0.0021467634
+ aigbacc = 0.012071
+ igcmod = 1
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ ku0we = -0.0007
+ ags = 0.29253015
+ aigbinv = 0.009974
+ beta0 = 13.32
+ keta = -0.031086208
+ leta0 = 0
+ cjd = 0.001346
+ cit = -0.00056559017
+ cjs = 0.001346
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 1.38228675e-8
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ lags = 5.1257474e-7
+ ppclm = 0
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 2.9285967e-10
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ kt1l = 0
+ la0 = -1.4357692e-8
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0
+ kt1 = -0.19916819
+ kt2 = -0.054700402
+ lk2 = 1.425099e-9
+ permod = 1
+ llc = -1.18e-13
+ lln = 0.7
+ lu0 = -4.8076045e-10
+ mjd = 0.335
+ mjs = 0.335
+ lua = -1.6078561e-16
+ lub = 5.7693033e-26
+ luc = -4.8483261e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ lint = 9.7879675e-9
+ pa0 = -2.613694e-13
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ pk2 = -5.5906497e-16
+ lkt1 = -1.3143224e-8
+ lkt2 = -3.9687861e-9
+ pu0 = -2.2461433e-17
+ lmax = 4.4908e-7
+ prt = 0
+ pua = 5.4100623e-23
+ pub = -6.3187687e-32
+ puc = -3.6550877e-24
+ pud = 0
+ dmcgt = 0
+ lmin = 2.1577e-7
+ poxedge = 1
+ tcjsw = 9.34e-5
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 1.2176874e-9
+ ub1 = -1.2376668e-18
+ lpe0 = 6.44e-8
+ uc1 = 1.0272662e-10
+ lpeb = 0
+ tpb = 0.0016
+ wa0 = 7.3504866e-7
+ ijthsfwd = 0.01
+ ute = -1
+ web = 6628.3
+ wec = -16935.0
+ wk2 = -1.4458115e-9
+ binunit = 2
+ voffcv = -0.125
+ wpemod = 1
+ wlc = 0
+ wln = 1
+ minv = -0.33
+ wu0 = 4.9034036e-11
+ xgl = -8.2e-9
+ xgw = 0
+ lua1 = 6.4190903e-17
+ lub1 = -1.6446372e-25
+ wua = -3.3214073e-16
+ wub = 1.7570216e-25
+ wuc = -9.9257962e-18
+ wud = 0
+ luc1 = 1.9195943e-18
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ ndep = 1e+18
+ bigsd = 0.0003327
+ lwlc = 0
+ moin = 5.5538
+ wvoff = 6.3544834e-9
+ nigc = 2.291
+ ijthsrev = 0.01
+ wvsat = -0.0097711764
+ wvth0 = 4.1127039e-10
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ waigc = 4.9938134e-12
+ tpbswg = 0.001
+ jtsswgd = 1.75e-7
+ pags = 2.5662868e-13
+ jtsswgs = 1.75e-7
+ ntox = 1
+ pcit = -8.1677938e-17
+ lketa = -2.0098347e-8
+ pclm = 1.5174437
+ xpart = 1
+ ppdiblc2 = -1.9289508e-16
+ phin = 0.15
+ ptvoff = -6.733506e-17
+ egidl = 0.001
+ waigsd = 1.9051377e-12
+ pkt1 = 4.9381461e-16
+ pkt2 = -1.2251691e-15
+ diomod = 1
+ pditsd = 0
+ pditsl = 0
+ rbdb = 50
+ cjswgd = 1.81e-10
+ pku0we = 0.0
+ pua1 = -4.1586322e-23
+ prwb = 0
+ pub1 = 2.600258e-32
+ prwg = 0
+ cjswgs = 1.81e-10
+ puc1 = -8.5761835e-25
+ njtsswg = 6.489
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ pkvth0we = 0.0
+ rdsw = 200
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ ckappad = 0.6
+ ckappas = 0.6
+ mjswgd = 0.95
+ mjswgs = 0.95
+ pdiblc1 = 0
+ pdiblc2 = 0.01380092
+ pvfbsdoff = 0
+ pdiblcb = 0
+ vfbsdoff = 0.01
+ pvoff = -8.886429e-16
+ tcjswg = 0.00128
+ cdscb = 0
+ cdscd = 0
+ pvsat = 0
+ wk2we = 0.0
+ pvth0 = 2.2840255e-16
+ drout = 0.56
+ paramchk = 1
+ rshg = 14.1
+ paigc = 1.0085061e-18
+ bigbacc = 0.0054401
+ voffl = 0
+ weta0 = -2.2161431e-9
+ kvth0we = -0.00022
+ wetab = 6.0440267e-8
+ lpclm = 0
+ lintnoi = -5e-9
+ fprout = 200
+ ijthdfwd = 0.01
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ xrcrg1 = 12
+ xrcrg2 = 1
+ cgidl = 1
+ tnom = 25
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ wtvoff = -1.0667978e-10
+ pbswd = 0.9
+ pbsws = 0.9
+ ijthdrev = 0.01
+ lpdiblc2 = -8.1587971e-10
+ capmod = 2
+ wags = -4.2059528e-7
+ wku0we = 1.5e-11
+ wcit = 1.8563168e-10
+ pdits = 0
+ cigsd = 0.013281
+ mobmod = 0
+ voff = -0.12166106
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ acde = 0.5
+ vsat = 121084.96
+ wint = 0
+ vth0 = -0.40344281
+ nfactor = 1
+ pk2we = 0.0
+ wkt1 = -7.6912059e-9
+ wkt2 = 2.6613072e-10
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ wmax = 9e-6
+ aigc = 0.0067878654
+ wmin = 9e-7
+ lkvth0we = 3e-12
+ tnoia = 0
+ a0 = 1.3739719
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 72000
+ wua1 = 3.3927227e-16
+ cf = 8.17e-11
+ wub1 = -2.6580249e-25
+ wuc1 = 1.6454797e-17
+ ef = 1.15
+ k1 = 0.30425
+ k2 = 0.00015642806
+ k3 = -2.5823
+ em = 20000000.0
+ peta0 = 0
+ ll = -1.18e-13
+ lw = 0
+ u0 = 0.010652861
+ w0 = 0
+ ua = 3.293471e-10
+ ub = 1.3083159e-18
+ uc = 4.2293442e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ bigc = 0.0012521
+ xw = 6e-9
+ wketa = 1.5506359e-8
+ wwlc = 0
+ acnqsmod = 0
+ tpbsw = 0.0025
+ nigbacc = 10
+ cjswd = 5.1e-11
+ cjsws = 5.1e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ cdsc = 0
+ cgbo = 0
+ rbodymod = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigc = 0.15259
+ wtvfbsdoff = 0
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ nigbinv = 2.171
+ ltvfbsdoff = 0
+ scref = 1e-6
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ pigcd = 2.572
+ wpdiblc2 = 1.6189099e-11
+ aigsd = 0.0063634291
+ fnoimod = 1
+ lvoff = -3.7843526e-9
+ eigbinv = 1.1
+ k2we = 5e-5
+ toxref = 3e-9
+ lvsat = 0
+ dsub = 0.5
+ dtox = 3.91e-10
+ lvth0 = 4.3151043e-9
+ ptvfbsdoff = 0
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ delta = 0.018814
+ laigc = -2.5231709e-11
+ tvfbsdoff = 0.1
+ rnoia = 0
+ rnoib = 0
+ eta0 = 0.16744607
+ etab = -0.23671111
+ )

.model pch_tt_13 pmos (
+ level = 54
+ pags = 7.0037917e-14
+ lku0we = 1.8e-11
+ pvth0 = -7.2768891e-16
+ drout = 0.56
+ epsrox = 3.9
+ ntox = 1
+ pcit = 3.1250046e-17
+ pclm = 1.5924795
+ paigc = -7.3857349e-19
+ voffl = 0
+ rdsmod = 0
+ phin = 0.15
+ igbmod = 1
+ weta0 = -2.2161431e-9
+ wetab = 6.0440267e-8
+ lkvth0we = 3e-12
+ pkt1 = 2.8071967e-16
+ pkt2 = -8.6151083e-16
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ lpclm = -1.5832542e-8
+ pbswgd = 0.8
+ pbswgs = 0.8
+ cgidl = 1
+ igcmod = 1
+ acnqsmod = 0
+ rbdb = 50
+ pua1 = -5.7774504e-23
+ prwb = 0
+ pub1 = 1.0356474e-31
+ prwg = 0
+ puc1 = 6.0450908e-24
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ rdsw = 200
+ rbodymod = 0
+ pbswd = 0.9
+ pbsws = 0.9
+ nfactor = 1
+ pdits = 0
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ permod = 1
+ rshg = 14.1
+ nigbacc = 10
+ wpdiblc2 = -2.9527442e-9
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ tnoia = 0
+ voffcv = -0.125
+ wpemod = 1
+ nigbinv = 2.171
+ peta0 = 0
+ tnom = 25
+ wketa = 2.8638443e-8
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ tpbsw = 0.0025
+ cjswd = 5.1e-11
+ cjsws = 5.1e-11
+ mjswd = 0.01
+ wkvth0we = 0.0
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ trnqsmod = 0
+ fnoimod = 1
+ eigbinv = 1.1
+ wags = 4.6372111e-7
+ tpbswg = 0.001
+ wcit = -3.4957204e-10
+ voff = -0.13366619
+ acde = 0.5
+ scref = 1e-6
+ vsat = 116618.55
+ wint = 0
+ vth0 = -0.40791428
+ rgatemod = 0
+ pigcd = 2.572
+ aigsd = 0.0063634291
+ wkt1 = -6.6812774e-9
+ wkt2 = -1.4573681e-9
+ tnjtsswg = 1
+ ptvoff = -1.8786066e-17
+ wmax = 9e-6
+ aigc = 0.0067673585
+ wmin = 9e-7
+ lvoff = -1.2512704e-9
+ waigsd = 1.9051377e-12
+ cigbacc = 0.245
+ lvsat = 0.00094241323
+ diomod = 1
+ lvth0 = 5.2585836e-9
+ wua1 = 4.1599351e-16
+ wub1 = -6.3339564e-25
+ wuc1 = -1.6259465e-17
+ tnoimod = 0
+ delta = 0.018814
+ laigc = -2.090475e-11
+ pditsd = 0
+ pditsl = 0
+ tvfbsdoff = 0.1
+ bigc = 0.0012521
+ cjswgd = 1.81e-10
+ pku0we = 0.0
+ cjswgs = 1.81e-10
+ wwlc = 0
+ rnoia = 0
+ rnoib = 0
+ cigbinv = 0.006
+ cdsc = 0
+ pketa = 2.2140676e-16
+ ngate = 1.7e+20
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ ngcon = 1
+ mjswgd = 0.95
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ mjswgs = 0.95
+ wpclm = -3.6917638e-7
+ cigc = 0.15259
+ tcjswg = 0.00128
+ version = 4.5
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ tempmod = 0
+ jswgs = 3.69e-13
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ aigbacc = 0.012071
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ k2we = 5e-5
+ fprout = 200
+ aigbinv = 0.009974
+ dsub = 0.5
+ dtox = 3.91e-10
+ xrcrg1 = 12
+ xrcrg2 = 1
+ ijthsfwd = 0.01
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ tvoff = 0.0019304691
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ ags = 2.6061153
+ wtvoff = -3.3676979e-10
+ eta0 = 0.16744607
+ etab = -0.23671111
+ cjd = 0.001346
+ cit = 0.00047888384
+ cjs = 0.001346
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 1.38228675e-8
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ ijthsrev = 0.01
+ ku0we = -0.0007
+ beta0 = 13.32
+ capmod = 2
+ leta0 = 0
+ la0 = -4.2186937e-8
+ poxedge = 1
+ wku0we = 1.5e-11
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0.00028821144
+ kt1 = -0.23884145
+ kt2 = -0.071460529
+ lk2 = 4.3288295e-9
+ llc = -1.18e-13
+ lln = 0.7
+ lu0 = -1.8451509e-10
+ mjd = 0.335
+ ppclm = 1.4344283e-14
+ mjs = 0.335
+ lua = -2.3141614e-17
+ lub = -3.0092793e-26
+ luc = -1.1168748e-18
+ lud = 0
+ lwc = 0
+ mobmod = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = -1.7418058e-15
+ nsd = 1e+20
+ binunit = 2
+ pbd = 0.75
+ pat = -2.5956322e-9
+ pbs = 0.75
+ pk2 = -2.0925962e-16
+ dlcig = 2.5e-9
+ pu0 = 6.8306111e-19
+ bgidl = 1834800000.0
+ prt = 0
+ pua = -2.4112447e-23
+ pub = 3.4375734e-32
+ puc = -1.1236355e-25
+ pud = 0
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 2.2048659e-9
+ ub1 = -2.7884819e-18
+ ppdiblc2 = 4.3354985e-16
+ uc1 = 8.0779763e-11
+ tpb = 0.0016
+ wa0 = -4.9541389e-7
+ ute = -1
+ wat = 0.012301575
+ web = 6628.3
+ wec = -16935.0
+ wk2 = -3.1036812e-9
+ wlc = 0
+ wln = 1
+ wu0 = -6.065551e-11
+ xgl = -8.2e-9
+ xgw = 0
+ wua = 3.8537331e-17
+ wub = -2.8668372e-25
+ wuc = -2.6715958e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ wtvfbsdoff = 0
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ bigsd = 0.0003327
+ ltvfbsdoff = 0
+ pkvth0we = 0.0
+ wvoff = 5.8569161e-9
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ wvsat = -0.0057246059
+ vfbsdoff = 0.01
+ keta = -0.13181891
+ wvth0 = 4.9425095e-9
+ waigc = 1.3273811e-11
+ lags = 2.4408277e-8
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 7.2475659e-11
+ a0 = 1.505864
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ kt1l = 0
+ ptvfbsdoff = 0
+ at = 70634.069
+ paramchk = 1
+ cf = 8.17e-11
+ lketa = 1.156253e-9
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.013605325
+ k3 = -2.5823
+ em = 20000000.0
+ ll = -1.18e-13
+ lw = 0
+ u0 = 0.0092488547
+ w0 = 0
+ xpart = 1
+ ua = -3.2299413e-10
+ ub = 1.7243624e-18
+ uc = 2.4608838e-11
+ ud = 0
+ njtsswg = 6.489
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 6e-9
+ lint = 9.7879675e-9
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ lkt1 = -4.7721669e-9
+ lkt2 = -4.3239941e-10
+ egidl = 0.001
+ lmax = 2.1577e-7
+ lmin = 9e-8
+ toxref = 3e-9
+ ckappad = 0.6
+ ckappas = 0.6
+ lpe0 = 6.44e-8
+ pdiblc1 = 0
+ pdiblc2 = 0.017260131
+ lpeb = 0
+ pdiblcb = 0
+ ijthdfwd = 0.01
+ minv = -0.33
+ lua1 = -1.4410376e-16
+ lub1 = 1.6275827e-25
+ luc1 = 6.550381e-18
+ ndep = 1e+18
+ lwlc = 0
+ moin = 5.5538
+ bigbacc = 0.0054401
+ nigc = 2.291
+ ltvoff = -6.4284173e-11
+ ijthdrev = 0.01
+ pvfbsdoff = 0
+ lpdiblc2 = -1.5457732e-9
+ kvth0we = -0.00022
+ pvoff = -7.836562e-16
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ cdscb = 0
+ cdscd = 0
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ pvsat = -8.5382639e-10
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ wk2we = 0.0
+ )

.model pch_tt_14 pmos (
+ level = 54
+ cjd = 0.001346
+ poxedge = 1
+ cit = -0.00080588346
+ wua1 = -1.4703955e-15
+ cjs = 0.001346
+ clc = 1e-7
+ cle = 0.6
+ wub1 = 2.631826e-24
+ bvd = 8.2
+ wuc1 = 2.762344e-16
+ bvs = 8.2
+ igcmod = 1
+ dlc = 4.0349e-9
+ k3b = 2.1176
+ tvoff = 0.0011122833
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ bigc = 0.0012521
+ wwlc = 0
+ xjbvd = 1
+ binunit = 2
+ xjbvs = 1
+ lk2we = 0.0
+ pkvth0we = 0.0
+ la0 = -2.3326483e-7
+ jsd = 1.5e-7
+ cdsc = 0
+ jss = 1.5e-7
+ lat = -0.0065502639
+ kt1 = -0.2764195
+ kt2 = -0.075556865
+ lk2 = 3.8809157e-9
+ llc = 0
+ cgbo = 0
+ lln = 1
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ lu0 = 2.0644492e-10
+ xtid = 3
+ xtis = 3
+ mjd = 0.335
+ mjs = 0.335
+ lua = 5.4621428e-17
+ lub = 1.4388057e-26
+ luc = 1.0238844e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ cgsl = 3.0105e-11
+ njs = 1.02
+ cgso = 2.6482e-11
+ pa0 = 5.4920056e-14
+ cigc = 0.15259
+ ku0we = -0.0007
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 1.0391973e-9
+ pbs = 0.75
+ pk2 = 6.854543e-16
+ beta0 = 13.32
+ vfbsdoff = 0.01
+ pu0 = -1.2707891e-16
+ leta0 = -6.4826039e-10
+ prt = 0
+ pua = -5.2218942e-24
+ pub = -3.6833051e-32
+ puc = -9.869134e-24
+ pud = 0
+ letab = 2.0996791e-8
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 8.9078668e-10
+ ub1 = -1.404024e-18
+ uc1 = 4.4088848e-11
+ ppclm = 7.4853015e-14
+ tpb = 0.0016
+ wa0 = -1.0981997e-6
+ ute = -1
+ wat = -0.026366825
+ web = 6628.3
+ wec = -16935.0
+ wk2 = -1.2621914e-8
+ wlc = 0
+ dlcig = 2.5e-9
+ permod = 1
+ wln = 1
+ wu0 = 1.2985144e-9
+ xgl = -8.2e-9
+ xgw = 0
+ bgidl = 1834800000.0
+ wua = -1.62426e-16
+ wub = 4.7085654e-25
+ wuc = 7.7079472e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ paramchk = 1
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ k2we = 5e-5
+ voffcv = -0.125
+ wpemod = 1
+ dsub = 0.5
+ dtox = 3.91e-10
+ ijthdfwd = 0.01
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ bigsd = 0.0003327
+ eta0 = 0.17434246
+ etab = -0.46008122
+ njtsswg = 6.489
+ wvoff = -4.5993296e-9
+ ijthdrev = 0.01
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ wvsat = -0.039767366
+ wvth0 = -1.6418701e-8
+ lpdiblc2 = 0
+ ckappad = 0.6
+ tpbswg = 0.001
+ ckappas = 0.6
+ waigc = -2.1370578e-11
+ pdiblc1 = 0
+ pdiblc2 = 0.00081573526
+ pdiblcb = 0
+ lketa = 9.0137227e-9
+ xpart = 1
+ ptvoff = 1.200911e-16
+ waigsd = 1.9051377e-12
+ bigbacc = 0.0054401
+ egidl = 0.001
+ lkvth0we = 3e-12
+ diomod = 1
+ kvth0we = -0.00022
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.81e-10
+ pku0we = 0.0
+ cjswgs = 1.81e-10
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ acnqsmod = 0
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ rbodymod = 0
+ mjswgd = 0.95
+ mjswgs = 0.95
+ pvfbsdoff = 0
+ tcjswg = 0.00128
+ keta = -0.21540901
+ pvoff = 1.9923089e-16
+ cdscb = 0
+ cdscd = 0
+ lags = -3.1969346e-8
+ pvsat = 2.3461931e-9
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ wk2we = 0.0
+ pvth0 = 1.2802649e-15
+ lcit = 1.9324378e-10
+ drout = 0.56
+ kt1l = 0
+ paigc = 2.5179991e-18
+ voffl = 0
+ wpdiblc2 = 1.6594883e-9
+ lint = 0
+ lkt1 = -1.2398309e-9
+ lkt2 = -4.7343777e-11
+ weta0 = 4.241971e-8
+ nfactor = 1
+ lmax = 9e-8
+ wetab = 1.3144359e-7
+ fprout = 200
+ lmin = 5.4e-8
+ lpclm = -1.0675035e-7
+ xrcrg1 = 12
+ xrcrg2 = 1
+ lpe0 = 6.44e-8
+ lpeb = 0
+ cgidl = 1
+ minv = -0.33
+ lua1 = -2.0580314e-17
+ lub1 = 3.261922e-26
+ luc1 = 9.999327e-18
+ wtvoff = -1.8141864e-9
+ ndep = 1e+18
+ lwlc = 0
+ moin = 5.5538
+ wkvth0we = 0.0
+ nigbacc = 10
+ pbswd = 0.9
+ nigc = 2.291
+ pbsws = 0.9
+ capmod = 2
+ trnqsmod = 0
+ wku0we = 1.5e-11
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ mobmod = 0
+ pdits = 0
+ nigbinv = 2.171
+ cigsd = 0.013281
+ pags = 2.8964227e-14
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ wtvfbsdoff = 0
+ ntox = 1
+ pcit = -6.9565404e-17
+ pclm = 2.5596902
+ rgatemod = 0
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ tnjtsswg = 1
+ ltvfbsdoff = 0
+ phin = 0.15
+ pkt1 = 7.7820041e-17
+ pkt2 = 1.7971063e-15
+ fnoimod = 1
+ tnoia = 0
+ eigbinv = 1.1
+ peta0 = -4.1957702e-15
+ petab = -6.6743123e-15
+ wketa = 8.0928346e-8
+ tpbsw = 0.0025
+ rbdb = 50
+ pua1 = 1.1954606e-22
+ prwb = 0
+ pub1 = -2.033661e-31
+ prwg = 0
+ puc1 = -2.1449333e-23
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ cjswd = 5.1e-11
+ pvag = 2.1
+ cjsws = 5.1e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ rdsw = 200
+ ptvfbsdoff = 0
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ cigbacc = 0.245
+ tnoimod = 0
+ rshg = 14.1
+ scref = 1e-6
+ pigcd = 2.572
+ cigbinv = 0.006
+ aigsd = 0.0063634291
+ lvoff = -2.6816163e-9
+ toxref = 3e-9
+ lvsat = -0.0059831154
+ lvth0 = -1.5502539e-9
+ version = 4.5
+ ijthsfwd = 0.01
+ delta = 0.018814
+ tvfbsdoff = 0.1
+ tempmod = 0
+ laigc = -1.5433256e-11
+ tnom = 25
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ rnoia = 0
+ rnoib = 0
+ aigbacc = 0.012071
+ ltvoff = 1.2625293e-11
+ pketa = -4.6938441e-15
+ a0 = 3.5386076
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ ngate = 1.7e+20
+ at = 143383.81
+ cf = 8.17e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.0088402851
+ k3 = -2.5823
+ ijthsrev = 0.01
+ em = 20000000.0
+ ngcon = 1
+ ll = 0
+ lw = 0
+ u0 = 0.0050897056
+ wpclm = -1.0128863e-6
+ w0 = 0
+ ua = -1.1502605e-9
+ ub = 1.2511619e-18
+ uc = -9.619668e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 6e-9
+ gbmin = 1e-12
+ wags = 9.0067526e-7
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ aigbinv = 0.009974
+ wcit = 7.2293275e-10
+ lku0we = 1.8e-11
+ wvfbsdoff = 0
+ epsrox = 3.9
+ lvfbsdoff = 0
+ voff = -0.11844975
+ acde = 0.5
+ vsat = 190294.39
+ ppdiblc2 = 0
+ rdsmod = 0
+ wint = 0
+ vth0 = -0.33547984
+ igbmod = 1
+ wkt1 = -4.5227706e-9
+ wkt2 = -2.9740529e-8
+ wmax = 9e-6
+ aigc = 0.0067091511
+ wmin = 9e-7
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ pbswgd = 0.8
+ ags = 3.2058772
+ pbswgs = 0.8
+ )

.model pch_tt_15 pmos (
+ level = 54
+ keta = 0.054978601
+ fnoimod = 1
+ pdits = 0
+ eigbinv = 1.1
+ cigsd = 0.013281
+ permod = 1
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 3.30566e-10
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ kt1l = 0
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ lint = 0
+ lkt1 = -1.3608112e-8
+ lkt2 = 1.0752811e-9
+ lmax = 5.4e-8
+ lmin = 4.5e-8
+ voffcv = -0.125
+ wpemod = 1
+ tnoia = 0
+ lpe0 = 6.44e-8
+ lpeb = 0
+ ijthsfwd = 0.01
+ cigbacc = 0.245
+ peta0 = 5.9496569e-15
+ petab = -1.9628815e-15
+ minv = -0.33
+ lua1 = -1.9488641e-18
+ lub1 = 6.8003561e-26
+ wketa = -5.4843946e-8
+ luc1 = -2.115524e-18
+ tpbsw = 0.0025
+ ndep = 1e+18
+ tnoimod = 0
+ cjswd = 5.1e-11
+ lwlc = 0
+ cjsws = 5.1e-11
+ moin = 5.5538
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ nigc = 2.291
+ cigbinv = 0.006
+ ijthsrev = 0.01
+ tpbswg = 0.001
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ version = 4.5
+ tempmod = 0
+ ntox = 1
+ pcit = -7.0617065e-17
+ pclm = 1.3082183
+ scref = 1e-6
+ ptvoff = 9.8606268e-17
+ ppdiblc2 = 0
+ pigcd = 2.572
+ aigsd = 0.0063634291
+ waigsd = 1.9051377e-12
+ aigbacc = 0.012071
+ phin = 0.15
+ lvoff = -4.1725981e-9
+ diomod = 1
+ pkt1 = 1.3948109e-14
+ pkt2 = -4.0388508e-15
+ lvsat = -0.00019489408
+ lvth0 = -2.0426855e-9
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.81e-10
+ pku0we = 0.0
+ cjswgs = 1.81e-10
+ tvfbsdoff = 0.1
+ delta = 0.018814
+ aigbinv = 0.009974
+ laigc = -9.3796225e-12
+ rnoia = 0
+ rnoib = 0
+ rbdb = 50
+ pua1 = -1.9221227e-22
+ prwb = 0
+ pub1 = 2.2863324e-31
+ prwg = 0
+ puc1 = 2.3602641e-23
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ pkvth0we = 0.0
+ rbsb = 50
+ pvag = 2.1
+ mjswgd = 0.95
+ mjswgs = 0.95
+ rdsw = 200
+ pketa = 3.1809489e-15
+ ngate = 1.7e+20
+ ngcon = 1
+ tcjswg = 0.00128
+ wpclm = 1.8421624e-6
+ vfbsdoff = 0.01
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ poxedge = 1
+ paramchk = 1
+ rshg = 14.1
+ binunit = 2
+ ags = 2.6546816
+ cjd = 0.001346
+ cit = -0.0031735079
+ cjs = 0.001346
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 4.0349e-9
+ fprout = 200
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ ijthdfwd = 0.01
+ la0 = -1.5436392e-7
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0.0043243403
+ kt1 = -0.063173267
+ kt2 = -0.094912467
+ lk2 = 4.2787193e-9
+ llc = 0
+ tvoff = 0.0053332949
+ lln = 1
+ lu0 = -6.1856189e-11
+ wtvoff = -1.4437583e-9
+ tnom = 25
+ mjd = 0.335
+ mjs = 0.335
+ lua = -3.3837758e-17
+ lub = -3.4072549e-26
+ luc = -2.4014309e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = -3.174587e-14
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ xjbvd = 1
+ xjbvs = 1
+ nsd = 1e+20
+ pbd = 0.75
+ pat = -5.2399134e-10
+ lk2we = 0.0
+ pbs = 0.75
+ pk2 = 5.1035691e-16
+ pu0 = -9.701894e-17
+ prt = 0
+ pua = -1.0296702e-22
+ pub = 1.290002e-31
+ puc = 2.16225e-23
+ pud = 0
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ rsh = 15.2
+ wtvfbsdoff = 0
+ tcj = 0.000832
+ ua1 = 5.6955479e-10
+ ub1 = -2.0140988e-18
+ uc1 = 2.5296559e-10
+ ijthdrev = 0.01
+ capmod = 2
+ tpb = 0.0016
+ wa0 = 3.9604044e-7
+ ute = -1
+ wat = 0.00058470362
+ ku0we = -0.0007
+ web = 6628.3
+ wec = -16935.0
+ wk2 = -9.6029938e-9
+ wku0we = 1.5e-11
+ wlc = 0
+ beta0 = 13.32
+ wln = 1
+ wu0 = 7.8023907e-10
+ xgl = -8.2e-9
+ xgw = 0
+ lpdiblc2 = 0
+ wua = 1.5228349e-15
+ wub = -2.3883374e-24
+ leta0 = -2.3797369e-9
+ wuc = -4.6587973e-16
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ letab = 1.0403109e-8
+ ltvfbsdoff = 0
+ mobmod = 0
+ wags = 1.4000585e-6
+ ppclm = -9.0739811e-14
+ wcit = 7.4106483e-10
+ voff = -0.092743162
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ acde = 0.5
+ vsat = 90497.467
+ wint = 0
+ vth0 = -0.32698964
+ wkt1 = -2.4366569e-7
+ wkt2 = 7.087942e-8
+ wmax = 9e-6
+ aigc = 0.0066047781
+ wmin = 9e-7
+ njtsswg = 6.489
+ dmcgt = 0
+ lkvth0we = 3e-12
+ tcjsw = 9.34e-5
+ ptvfbsdoff = 0
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ wua1 = 3.9047481e-15
+ wub1 = -4.8164385e-24
+ wuc1 = -5.0052376e-16
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.00081573526
+ pdiblcb = 0
+ bigc = 0.0012521
+ acnqsmod = 0
+ wwlc = 0
+ bigsd = 0.0003327
+ cdsc = 0
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ wvoff = 1.0199556e-9
+ rbodymod = 0
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigc = 0.15259
+ wvsat = -0.0078232946
+ bigbacc = 0.0054401
+ wvth0 = 4.8192399e-8
+ waigc = 1.173226e-10
+ kvth0we = -0.00022
+ lintnoi = -5e-9
+ lketa = -6.6687589e-9
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ xpart = 1
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ wpdiblc2 = 1.6594883e-9
+ toxref = 3e-9
+ egidl = 0.001
+ k2we = 5e-5
+ dsub = 0.5
+ dtox = 3.91e-10
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ eta0 = 0.2041955
+ etab = -0.27743155
+ ltvoff = -2.3219338e-10
+ wkvth0we = 0.0
+ pvfbsdoff = 0
+ trnqsmod = 0
+ nfactor = 1
+ pvoff = -1.2668765e-16
+ lku0we = 1.8e-11
+ cdscb = 0
+ cdscd = 0
+ epsrox = 3.9
+ pvsat = 4.9343693e-10
+ wk2we = 0.0
+ pvth0 = -2.4671789e-15
+ drout = 0.56
+ paigc = -5.5262052e-18
+ rdsmod = 0
+ igbmod = 1
+ rgatemod = 0
+ voffl = 0
+ tnjtsswg = 1
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ nigbacc = 10
+ weta0 = -1.3250145e-7
+ wetab = 5.0212024e-8
+ pbswgd = 0.8
+ pbswgs = 0.8
+ lpclm = -3.4164983e-8
+ a0 = 2.1782471
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = -44109.368
+ cf = 8.17e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.015698968
+ k3 = -2.5823
+ em = 20000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.0097155868
+ w0 = 0
+ igcmod = 1
+ ua = 3.7489785e-10
+ ub = 2.0866896e-18
+ uc = 4.9437493e-10
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 6e-9
+ cgidl = 1
+ nigbinv = 2.171
+ pbswd = 0.9
+ pbsws = 0.9
+ )

.model pch_tt_16 pmos (
+ level = 54
+ wpdiblc2 = 1.6594883e-9
+ voffcv = -0.125
+ wpemod = 1
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ bigbacc = 0.0054401
+ tnom = 25
+ kvth0we = -0.00022
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ bigsd = 0.0003327
+ lintnoi = -5e-9
+ wkvth0we = 0.0
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ wvoff = -9.7608128e-9
+ trnqsmod = 0
+ wvsat = -0.0020201595
+ tpbswg = 0.001
+ wvth0 = 7.6331233e-9
+ wags = 3.1454838e-6
+ waigc = -1.1150212e-11
+ wcit = -4.2593599e-9
+ voff = -0.099237323
+ acde = 0.5
+ lketa = 8.2510741e-9
+ ptvoff = -1.3565734e-16
+ xpart = 1
+ waigsd = 2.0479558e-12
+ vsat = 122744.64
+ wint = 0
+ rgatemod = 0
+ vth0 = -0.36923313
+ wkt1 = 3.1251908e-7
+ wkt2 = -1.0928272e-8
+ tnjtsswg = 1
+ wmax = 9e-6
+ aigc = 0.0065575398
+ wmin = 9e-7
+ diomod = 1
+ egidl = 0.001
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.81e-10
+ pku0we = 0.0
+ cjswgs = 1.81e-10
+ nfactor = 1
+ wua1 = -3.8771176e-15
+ wub1 = 4.4904637e-24
+ wuc1 = 9.3089203e-17
+ bigc = 0.0012521
+ wwlc = 0
+ mjswgd = 0.95
+ mjswgs = 0.95
+ pvfbsdoff = 0
+ cdsc = 0
+ tcjswg = 0.00128
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigc = 0.15259
+ nigbacc = 10
+ pvoff = 4.0157e-16
+ cdscb = 0
+ cdscd = 0
+ pvsat = 2.0908331e-10
+ wk2we = 0.0
+ pvth0 = -4.797744e-16
+ drout = 0.56
+ paigc = 7.6896258e-19
+ nigbinv = 2.171
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ voffl = 0
+ dmdg = 0
+ fprout = 200
+ weta0 = 4.9304045e-9
+ xrcrg1 = 12
+ xrcrg2 = 1
+ wetab = 3.974597e-8
+ wtvfbsdoff = 0
+ lpclm = -2.1829165e-8
+ k2we = 5e-5
+ dsub = 0.5
+ dtox = 3.91e-10
+ ijthsfwd = 0.01
+ wtvoff = 3.3371317e-9
+ cgidl = 1
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ fnoimod = 1
+ ltvfbsdoff = 0
+ eigbinv = 1.1
+ eta0 = 0.11033512
+ etab = -0.14869011
+ capmod = 2
+ pbswd = 0.9
+ pbsws = 0.9
+ ijthsrev = 0.01
+ wku0we = 1.5e-11
+ mobmod = 0
+ pdits = 0
+ cigsd = 0.013281
+ ptvfbsdoff = 0
+ cigbacc = 0.245
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ ppdiblc2 = 0
+ tnoimod = 0
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ laigsd = 7.7486946e-16
+ cigbinv = 0.006
+ tnoia = 0
+ peta0 = -7.8450381e-16
+ petab = -1.4500449e-15
+ wketa = 4.9202854e-8
+ version = 4.5
+ tpbsw = 0.0025
+ tempmod = 0
+ cjswd = 5.1e-11
+ pkvth0we = 0.0
+ cjsws = 5.1e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ agidl = 3.2166e-9
+ aigbacc = 0.012071
+ vfbsdoff = 0.01
+ keta = -0.24950779
+ lags = 9.4399385e-8
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 1.9950138e-10
+ aigbinv = 0.009974
+ kt1l = 0
+ paramchk = 1
+ scref = 1e-6
+ pigcd = 2.572
+ aigsd = 0.0063634133
+ toxref = 3e-9
+ lint = 0
+ lvoff = -3.8543842e-9
+ lkt1 = -1.1161514e-10
+ lkt2 = 4.9336152e-10
+ lmax = 4.5e-8
+ lmin = 3.6e-8
+ lpe0 = 6.44e-8
+ lvsat = -0.0017750054
+ lpeb = 0
+ tvfbsdoff = 0.1
+ lvth0 = 2.7245694e-11
+ ijthdfwd = 0.01
+ delta = 0.018814
+ laigc = -7.0649434e-12
+ minv = -0.33
+ lua1 = -6.8231177e-17
+ lub1 = 7.1697841e-26
+ luc1 = 2.786749e-18
+ poxedge = 1
+ rnoia = 0
+ rnoib = 0
+ ndep = 1e+18
+ ltvoff = -9.8738127e-12
+ lwlc = 0
+ moin = 5.5538
+ binunit = 2
+ pketa = -1.9173443e-15
+ ngate = 1.7e+20
+ nigc = 2.291
+ ijthdrev = 0.01
+ ngcon = 1
+ wpclm = -3.2091624e-7
+ lpdiblc2 = 0
+ gbmin = 1e-12
+ lku0we = 1.8e-11
+ noff = 2.2684
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ epsrox = 3.9
+ ags = 0.72816353
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ cjd = 0.001346
+ cit = -0.00049871975
+ cjs = 0.001346
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ pags = -8.5525843e-14
+ dlc = 4.0349e-9
+ k3b = 2.1176
+ rdsmod = 0
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ ntox = 1
+ pcit = 1.7440375e-16
+ pclm = 1.0564669
+ igbmod = 1
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ la0 = -3.7737017e-8
+ jsd = 1.5e-7
+ phin = 0.15
+ jss = 1.5e-7
+ lat = -0.0019151022
+ jtsswgd = 1.75e-7
+ kt1 = -0.33861198
+ kt2 = -0.083036557
+ lk2 = 4.0583258e-9
+ jtsswgs = 1.75e-7
+ llc = 0
+ lln = 1
+ pbswgd = 0.8
+ pbswgs = 0.8
+ lu0 = 1.5317989e-10
+ mjd = 0.335
+ mjs = 0.335
+ lua = 2.9640356e-17
+ lub = 1.5163389e-26
+ luc = -2.5002144e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ lkvth0we = 3e-12
+ njd = 1.02
+ njs = 1.02
+ pa0 = -1.5136929e-14
+ pkt1 = -1.3304944e-14
+ pkt2 = -3.0273858e-17
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 2.5964497e-9
+ pbs = 0.75
+ pk2 = 4.883387e-16
+ igcmod = 1
+ pu0 = -4.5849539e-17
+ prt = 0
+ pua = 8.5912273e-23
+ pub = -1.727672e-31
+ puc = 8.2880171e-25
+ pud = 0
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 1.9222551e-9
+ ub1 = -2.0894923e-18
+ uc1 = 1.529192e-10
+ tvoff = 0.00079616085
+ tpb = 0.0016
+ wa0 = 5.7082474e-8
+ acnqsmod = 0
+ xjbvd = 1
+ ute = -1
+ wat = -0.063097766
+ xjbvs = 1
+ web = 6628.3
+ wec = -16935.0
+ rbdb = 50
+ wk2 = -9.1536426e-9
+ pua1 = 1.8909915e-22
+ prwb = 0
+ lk2we = 0.0
+ pub1 = -2.2740497e-31
+ prwg = 0
+ puc1 = -5.4843946e-24
+ wlc = 0
+ wln = 1
+ wu0 = -2.6403442e-10
+ xgl = -8.2e-9
+ rbpb = 50
+ rbpd = 50
+ xgw = 0
+ rbps = 50
+ rbsb = 50
+ wua = -2.3318447e-15
+ pvag = 2.1
+ wub = 3.770181e-24
+ wuc = -4.1518546e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ rdsw = 200
+ rbodymod = 0
+ paigsd = -6.9980875e-21
+ ku0we = -0.0007
+ beta0 = 13.32
+ njtsswg = 6.489
+ leta0 = 2.2194218e-9
+ letab = 4.094779e-9
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ ppclm = 1.5251044e-14
+ permod = 1
+ a0 = -0.20189383
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ ckappad = 0.6
+ at = 83226.192
+ cf = 8.17e-11
+ ckappas = 0.6
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.01120114
+ k3 = -2.5823
+ em = 20000000.0
+ dlcig = 2.5e-9
+ pdiblc1 = 0
+ pdiblc2 = 0.00081573526
+ ll = 0
+ lw = 0
+ bgidl = 1834800000.0
+ u0 = 0.0053270954
+ w0 = 0
+ pdiblcb = 0
+ ua = -9.2057386e-10
+ ub = 1.0818745e-18
+ uc = 5.5311765e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 6e-9
+ rshg = 14.1
+ )

.model pch_tt_17 pmos (
+ level = 54
+ tpbsw = 0.0025
+ aigbinv = 0.009974
+ eta0 = 0.191845
+ cjswd = 5.1e-11
+ cjsws = 5.1e-11
+ etab = -0.18516667
+ a0 = 2.6112
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ at = 72000
+ cf = 8.17e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.0045864754
+ k3 = -2.5823
+ em = 20000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.0097059667
+ w0 = 0
+ ua = 1.9119717e-10
+ ub = 1.0765761e-18
+ uc = -8.28048e-12
+ ud = 0
+ ijthdrev = 0.01
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 6e-9
+ tpbswg = 0.001
+ lpdiblc2 = 0
+ ptvoff = 0
+ waigsd = 1.9350626e-12
+ scref = 1e-6
+ poxedge = 1
+ pigcd = 2.572
+ aigsd = 0.0063633642
+ diomod = 1
+ binunit = 2
+ lvoff = 0
+ pditsd = 0
+ lkvth0we = 3e-12
+ pditsl = 0
+ cjswgd = 1.81e-10
+ pku0we = 0.0
+ cjswgs = 1.81e-10
+ tvfbsdoff = 0.1
+ lvsat = 0
+ lvth0 = 0
+ delta = 0.018814
+ acnqsmod = 0
+ rnoia = 0
+ rnoib = 0
+ mjswgd = 0.95
+ mjswgs = 0.95
+ tcjswg = 0.00128
+ ngate = 1.7e+20
+ rbodymod = 0
+ ags = 0.98525249
+ ngcon = 1
+ wpclm = -5.08417e-8
+ cjd = 0.001346
+ cit = 5e-6
+ cjs = 0.001346
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ dlc = 1.0572421799999999e-8
+ k3b = 2.1176
+ dwb = 0
+ keta = -0.016063969
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ gbmin = 1e-12
+ wvfbsdoff = 0
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ lvfbsdoff = 0
+ wtvfbsdoff = 0
+ la0 = 0
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0
+ lcit = 0
+ kt1 = -0.18299632
+ lk2 = 0
+ kt2 = -0.042133438
+ llc = 0
+ lln = 1
+ lu0 = 0
+ mjd = 0.335
+ kt1l = 0
+ mjs = 0.335
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 0
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ ltvfbsdoff = 0
+ pk2 = 0
+ wpdiblc2 = -1.7580235e-10
+ fprout = 200
+ pu0 = 0
+ prt = 0
+ pud = 0
+ lint = 6.5375218e-9
+ xrcrg1 = 12
+ xrcrg2 = 1
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 1.45515e-9
+ ub1 = -1.5029257e-18
+ uc1 = -4.3667733e-11
+ lkt1 = 0
+ lmax = 2.001e-5
+ tpb = 0.0016
+ wa0 = 2.308488e-7
+ lmin = 8.9991e-6
+ ute = -0.96728333
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 1.3953799e-9
+ njtsswg = 6.489
+ lpe0 = 6.44e-8
+ wlc = 0
+ wln = 1
+ wu0 = 2.7482e-12
+ xgl = -8.2e-9
+ lpeb = 0
+ xgw = 0
+ wua = -1.5682603e-16
+ wub = 3.5681818e-26
+ wuc = 4.8873989e-18
+ wud = 0
+ wtvoff = -7.2458121e-11
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ tvoff = 0.0025973351
+ minv = -0.33
+ xjbvd = 1
+ xjbvs = 1
+ ckappad = 0.6
+ ckappas = 0.6
+ lk2we = 0.0
+ ndep = 1e+18
+ pdiblc1 = 0
+ pdiblc2 = 0.0032290423
+ pdiblcb = 0
+ lwlc = 0
+ ptvfbsdoff = 0
+ capmod = 2
+ wkvth0we = 0.0
+ moin = 5.5538
+ wku0we = 1.5e-11
+ nigc = 2.291
+ trnqsmod = 0
+ mobmod = 0
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = 0
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ bigbacc = 0.0054401
+ ppclm = 0
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ kvth0we = -0.00022
+ ntox = 1
+ pcit = 0
+ pclm = 1.2411167
+ rgatemod = 0
+ lintnoi = -5e-9
+ tnjtsswg = 1
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ phin = 0.15
+ vtsswgs = 1.1
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ pkt1 = 0
+ bigsd = 0.0003327
+ rbdb = 50
+ prwb = 0
+ prwg = 0
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ rdsw = 200
+ wvoff = 3.276885e-9
+ wvsat = -0.017628054
+ wvth0 = 1.0594256e-9
+ waigc = -7.2361068e-12
+ nfactor = 1
+ lketa = 0
+ rshg = 14.1
+ xpart = 1
+ toxref = 3e-9
+ egidl = 0.001
+ nigbacc = 10
+ ijthsfwd = 0.01
+ tnom = 25
+ ltvoff = 0
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ pvfbsdoff = 0
+ nigbinv = 2.171
+ ijthsrev = 0.01
+ lku0we = 1.8e-11
+ pvoff = 0
+ epsrox = 3.9
+ wags = -3.1938756e-8
+ cdscb = 0
+ cdscd = 0
+ pvsat = 0
+ wk2we = 0.0
+ rdsmod = 0
+ pvth0 = 0
+ fnoimod = 1
+ drout = 0.56
+ voff = -0.10917042
+ igbmod = 1
+ acde = 0.5
+ eigbinv = 1.1
+ ppdiblc2 = 0
+ vsat = 129757.01
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ wint = 0
+ voffl = 0
+ vth0 = -0.38324647
+ wkt1 = 1.4804073e-9
+ wkt2 = -8.3218931e-9
+ pbswgd = 0.8
+ pbswgs = 0.8
+ wmax = 9e-7
+ aigc = 0.0068422292
+ wmin = 5.4e-7
+ weta0 = -2.432157e-8
+ wetab = 1.3741e-8
+ igcmod = 1
+ lpclm = 0
+ wua1 = -5.289391e-16
+ wub1 = 6.5622425e-25
+ wuc1 = 2.3227786e-17
+ cgidl = 1
+ bigc = 0.0012521
+ wute = -1.003093e-7
+ cigbacc = 0.245
+ wwlc = 0
+ pkvth0we = 0.0
+ cdsc = 0
+ tnoimod = 0
+ pbswd = 0.9
+ pbsws = 0.9
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigc = 0.15259
+ vfbsdoff = 0.01
+ cigbinv = 0.006
+ permod = 1
+ pdits = 0
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ paramchk = 1
+ version = 4.5
+ tempmod = 0
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ voffcv = -0.125
+ wpemod = 1
+ aigbacc = 0.012071
+ k2we = 5e-5
+ tnoia = 0
+ dsub = 0.5
+ dtox = 3.91e-10
+ ijthdfwd = 0.01
+ peta0 = 0
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ wketa = -3.7023239e-9
+ )

.model pch_tt_18 pmos (
+ level = 54
+ waigc = -9.2878513e-12
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ nigbacc = 10
+ ptvoff = 6.0745993e-16
+ pags = -1.6587566e-14
+ waigsd = 1.93751e-12
+ lketa = -8.0782883e-8
+ ntox = 1
+ pcit = 0
+ pclm = 1.2411167
+ xpart = 1
+ ppdiblc2 = 2.0750737e-15
+ diomod = 1
+ nigbinv = 2.171
+ phin = 0.15
+ egidl = 0.001
+ pditsd = 0
+ pditsl = 0
+ a0 = 2.6572474
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ cjswgd = 1.81e-10
+ pku0we = 0.0
+ cjswgs = 1.81e-10
+ at = 72000
+ cf = 8.17e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.0050849127
+ k3 = -2.5823
+ em = 20000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.0095857581
+ pkt1 = 7.4878862e-15
+ pkt2 = 7.624365e-15
+ w0 = 0
+ ua = 1.8022848e-10
+ ub = 1.0497212e-18
+ uc = -5.9216956e-12
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 6e-9
+ mjswgd = 0.95
+ mjswgs = 0.95
+ rbdb = 50
+ pua1 = 3.0135942e-22
+ prwb = 0
+ pub1 = -6.7644414e-31
+ prwg = 0
+ fnoimod = 1
+ puc1 = -4.7294542e-23
+ pvfbsdoff = 0
+ wtvfbsdoff = 0
+ tcjswg = 0.00128
+ pkvth0we = 0.0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ eigbinv = 1.1
+ pute = 3.5290383e-14
+ rdsw = 200
+ ltvfbsdoff = 0
+ vfbsdoff = 0.01
+ pvoff = 7.9887382e-16
+ cdscb = 0
+ cdscd = 0
+ pvsat = 0
+ wk2we = 0.0
+ pvth0 = -1.1664924e-15
+ drout = 0.56
+ paramchk = 1
+ paigc = 1.8445184e-17
+ rshg = 14.1
+ cigbacc = 0.245
+ fprout = 200
+ voffl = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ tnoimod = 0
+ ptvfbsdoff = 0
+ weta0 = -2.432157e-8
+ wetab = 1.3741e-8
+ lpclm = 0
+ wtvoff = -1.4002875e-10
+ cigbinv = 0.006
+ ijthdfwd = 0.01
+ cgidl = 1
+ tnom = 25
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ capmod = 2
+ version = 4.5
+ wku0we = 1.5e-11
+ tempmod = 0
+ pbswd = 0.9
+ pbsws = 0.9
+ ijthdrev = 0.01
+ mobmod = 0
+ lpdiblc2 = 3.0626629e-9
+ aigbacc = 0.012071
+ wags = -3.0093643e-8
+ pdits = 0
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ voff = -0.10728654
+ acde = 0.5
+ vsat = 129757.01
+ aigbinv = 0.009974
+ wint = 0
+ vth0 = -0.38217796
+ laigsd = 5.7445099e-14
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ wkt1 = 6.4749443e-10
+ wkt2 = -9.1699871e-9
+ wmax = 9e-7
+ aigc = 0.0068507406
+ wmin = 5.4e-7
+ lkvth0we = 3e-12
+ tnoia = 0
+ peta0 = 0
+ wua1 = -5.6246072e-16
+ wub1 = 7.3146831e-25
+ wuc1 = 2.8488581e-17
+ wketa = -8.2059163e-9
+ bigc = 0.0012521
+ wute = -1.0423482e-7
+ acnqsmod = 0
+ tpbsw = 0.0025
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ wwlc = 0
+ cjswd = 5.1e-11
+ cjsws = 5.1e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ poxedge = 1
+ cdsc = 0
+ rbodymod = 0
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigc = 0.15259
+ binunit = 2
+ toxref = 3e-9
+ scref = 1e-6
+ pigcd = 2.572
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ wpdiblc2 = -4.0662257e-10
+ aigsd = 0.0063633578
+ dmdg = 0
+ lvoff = -1.6936099e-8
+ tvfbsdoff = 0.1
+ k2we = 5e-5
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ lvsat = 0
+ lvth0 = -9.6058678e-9
+ dsub = 0.5
+ dtox = 3.91e-10
+ delta = 0.018814
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ laigc = -7.651731e-11
+ ltvoff = -1.5996918e-9
+ ags = 0.95300429
+ rnoia = 0
+ rnoib = 0
+ cjd = 0.001346
+ cit = 5e-6
+ cjs = 0.001346
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 1.0572421799999999e-8
+ k3b = 2.1176
+ eta0 = 0.191845
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ etab = -0.18516667
+ dwj = 0
+ wkvth0we = 0.0
+ pketa = 4.0487295e-14
+ ngate = 1.7e+20
+ ngcon = 1
+ wpclm = -5.08417e-8
+ trnqsmod = 0
+ la0 = -4.1396638e-7
+ lku0we = 1.8e-11
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0
+ kt1 = -0.17852273
+ kt2 = -0.039741464
+ lk2 = 4.4809517e-9
+ llc = 0
+ lln = 1
+ epsrox = 3.9
+ lu0 = 1.0806753e-9
+ mjd = 0.335
+ wvfbsdoff = 0
+ mjs = 0.335
+ lua = 9.8608496e-17
+ lub = 2.4142536e-25
+ luc = -2.1205472e-17
+ lud = 0
+ gbmin = 1e-12
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ lvfbsdoff = 0
+ njd = 1.02
+ njs = 1.02
+ pa0 = -1.9681175e-13
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ pk2 = -1.7465146e-15
+ njtsswg = 6.489
+ pu0 = -2.7146448e-18
+ rdsmod = 0
+ prt = 0
+ pua = -5.0852536e-23
+ pub = 3.3773548e-32
+ puc = 2.1258791e-23
+ pud = 0
+ igbmod = 1
+ xtsswgd = 0.32
+ rsh = 15.2
+ xtsswgs = 0.32
+ tcj = 0.000832
+ ua1 = 1.3709274e-9
+ ub1 = -1.4287011e-18
+ uc1 = -6.3574807e-11
+ tpb = 0.0016
+ wa0 = 2.527411e-7
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ ute = -0.97152091
+ ckappad = 0.6
+ ckappas = 0.6
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 1.5896529e-9
+ wlc = 0
+ rgatemod = 0
+ wln = 1
+ pdiblc1 = 0
+ pdiblc2 = 0.0028883679
+ wu0 = 3.0501627e-12
+ xgl = -8.2e-9
+ xgw = 0
+ pbswgd = 0.8
+ pdiblcb = 0
+ wua = -1.5116947e-16
+ pbswgs = 0.8
+ wub = 3.1925028e-26
+ wuc = 2.5226836e-18
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ tnjtsswg = 1
+ igcmod = 1
+ tvoff = 0.0027752763
+ bigbacc = 0.0054401
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ kvth0we = -0.00022
+ paigsd = -2.2002196e-20
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ ku0we = -0.0007
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ beta0 = 13.32
+ leta0 = 0
+ keta = -0.0070781088
+ permod = 1
+ ppclm = 0
+ lags = 2.8991134e-7
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ dlcig = 2.5e-9
+ lcit = 0
+ bgidl = 1834800000.0
+ kt1l = 0
+ voffcv = -0.125
+ wpemod = 1
+ lint = 6.5375218e-9
+ lkt1 = -4.0217527e-8
+ lkt2 = -2.1503841e-8
+ dmcgt = 0
+ lmax = 8.9991e-6
+ tcjsw = 9.34e-5
+ lmin = 8.9908e-7
+ lpe0 = 6.44e-8
+ lpeb = 0
+ ijthsfwd = 0.01
+ minv = -0.33
+ lua1 = 7.5716104e-16
+ lub1 = -6.6727951e-25
+ luc1 = 1.7896459e-16
+ nfactor = 1
+ bigsd = 0.0003327
+ ndep = 1e+18
+ lute = 3.8095772e-8
+ lwlc = 0
+ moin = 5.5538
+ wvoff = 3.1880225e-9
+ tpbswg = 0.001
+ ijthsrev = 0.01
+ nigc = 2.291
+ wvsat = -0.017628054
+ wvth0 = 1.18918e-9
+ noff = 2.2684
+ )

.model pch_tt_19 pmos (
+ level = 54
+ cjd = 0.001346
+ cit = -8.7888889e-5
+ cjs = 0.001346
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ lvsat = 0
+ dlc = 1.0572421799999999e-8
+ k3b = 2.1176
+ lvth0 = -1.6657388e-10
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ ltvfbsdoff = 0
+ wua1 = -6.1430214e-16
+ wub1 = 1.1920544e-25
+ delta = 0.018814
+ wuc1 = -4.9561039e-17
+ laigc = -1.8208261e-11
+ mjswgd = 0.95
+ mjswgs = 0.95
+ njtsswg = 6.489
+ bigc = 0.0012521
+ wute = -1.2773023e-7
+ rnoia = 0
+ rnoib = 0
+ la0 = -9.6086602e-7
+ wwlc = 0
+ tcjswg = 0.00128
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0
+ kt1 = -0.20738899
+ kt2 = -0.065812764
+ lk2 = -2.3080411e-10
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ llc = 0
+ lln = 1
+ lu0 = -1.5282408e-9
+ mjd = 0.335
+ mjs = 0.335
+ lua = -3.205013e-16
+ lub = -3.7552526e-26
+ luc = 5.1848161e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 2.9499704e-13
+ pketa = -2.8529622e-14
+ ckappad = 0.6
+ cdsc = 0
+ ckappas = 0.6
+ ngate = 1.7e+20
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ pk2 = 8.8602334e-16
+ pdiblc1 = 0
+ pdiblc2 = -8.9657994e-6
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ ngcon = 1
+ xtis = 3
+ pdiblcb = 0
+ pu0 = 4.0536683e-16
+ wpclm = -5.08417e-8
+ prt = 0
+ pua = 3.1718399e-23
+ pub = 9.4535502e-32
+ puc = -3.7711192e-23
+ pud = 0
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigc = 0.15259
+ rsh = 15.2
+ wvfbsdoff = 0
+ tcj = 0.000832
+ ua1 = 2.985915e-9
+ ub1 = -2.7037422e-18
+ uc1 = 1.5248758e-10
+ lvfbsdoff = 0
+ gbmin = 1e-12
+ tpb = 0.0016
+ wa0 = -2.9985305e-7
+ jswgd = 3.69e-13
+ ptvfbsdoff = 0
+ jswgs = 3.69e-13
+ ute = -0.85901741
+ web = 6628.3
+ wec = -16935.0
+ wk2 = -1.3682549e-9
+ a0 = 3.2717414
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ wlc = 0
+ wln = 1
+ wu0 = -4.5546835e-10
+ at = 72000
+ cf = 8.17e-11
+ xgl = -8.2e-9
+ ef = 1.15
+ k1 = 0.30425
+ k2 = 0.00020919492
+ xgw = 0
+ k3 = -2.5823
+ em = 20000000.0
+ wua = -2.439458e-16
+ wub = -3.6346832e-26
+ wuc = 6.8781092e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ ll = 0
+ lw = 0
+ u0 = 0.012517124
+ w0 = 0
+ ua = 6.5113837e-10
+ ub = 1.3631795e-18
+ uc = -8.8004429e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 6e-9
+ bigbacc = 0.0054401
+ fprout = 200
+ xrcrg1 = 12
+ xrcrg2 = 1
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ kvth0we = -0.00022
+ lintnoi = -5e-9
+ wtvoff = 9.9743807e-10
+ bigbinv = 0.00149
+ k2we = 5e-5
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ dsub = 0.5
+ dtox = 3.91e-10
+ ijthsfwd = 0.01
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ tvoff = 0.00044287651
+ capmod = 2
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ wku0we = 1.5e-11
+ eta0 = 0.191845
+ etab = -0.18516667
+ mobmod = 0
+ ijthsrev = 0.01
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = 0
+ ppclm = 0
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ nfactor = 1
+ laigsd = -3.6354984e-15
+ ppdiblc2 = -2.7249029e-15
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ nigbacc = 10
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ bigsd = 0.0003327
+ pkvth0we = 0.0
+ wvoff = 1.2743983e-8
+ nigbinv = 2.171
+ wvsat = -0.017628054
+ vfbsdoff = 0.01
+ wvth0 = -7.3071142e-10
+ keta = -0.13767457
+ waigc = 2.7297355e-11
+ lags = 8.1183869e-8
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 8.2671111e-11
+ toxref = 3e-9
+ paramchk = 1
+ lketa = 3.5447968e-8
+ kt1l = 0
+ xpart = 1
+ fnoimod = 1
+ eigbinv = 1.1
+ lint = 6.5375218e-9
+ egidl = 0.001
+ lkt1 = -1.4526561e-8
+ lkt2 = 1.6996159e-9
+ lmax = 8.9908e-7
+ lmin = 4.4908e-7
+ lpe0 = 6.44e-8
+ lpeb = 0
+ ijthdfwd = 0.01
+ ltvoff = 4.7614406e-10
+ minv = -0.33
+ lua1 = -6.8017788e-16
+ lub1 = 4.6750711e-25
+ luc1 = -1.3330934e-17
+ pvfbsdoff = 0
+ ndep = 1e+18
+ lute = -6.2032341e-8
+ lwlc = 0
+ moin = 5.5538
+ cigbacc = 0.245
+ ijthdrev = 0.01
+ nigc = 2.291
+ lku0we = 1.8e-11
+ epsrox = 3.9
+ tnoimod = 0
+ lpdiblc2 = 5.64129e-9
+ pvoff = -7.7059313e-15
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ rdsmod = 0
+ cdscb = 0
+ cdscd = 0
+ cigbinv = 0.006
+ igbmod = 1
+ pvsat = 0
+ wk2we = 0.0
+ pvth0 = 5.4221102e-16
+ drout = 0.56
+ pags = 2.5130854e-13
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ paigc = -1.411565e-17
+ ntox = 1
+ pcit = 0
+ pclm = 1.2411167
+ pbswgd = 0.8
+ pbswgs = 0.8
+ voffl = 0
+ version = 4.5
+ igcmod = 1
+ phin = 0.15
+ tempmod = 0
+ weta0 = -2.432157e-8
+ wetab = 1.3741e-8
+ lkvth0we = 3e-12
+ lpclm = 0
+ pkt1 = -4.6411548e-15
+ pkt2 = -3.0623252e-15
+ aigbacc = 0.012071
+ cgidl = 1
+ acnqsmod = 0
+ rbdb = 50
+ pua1 = 3.4749829e-22
+ prwb = 0
+ pub1 = -1.3153018e-31
+ prwg = 0
+ puc1 = 2.216962e-23
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ paigsd = 1.9849821e-21
+ rbsb = 50
+ pvag = 2.1
+ pute = 5.6201301e-14
+ rdsw = 200
+ rbodymod = 0
+ pbswd = 0.9
+ pbsws = 0.9
+ aigbinv = 0.009974
+ permod = 1
+ pdits = 0
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ rshg = 14.1
+ voffcv = -0.125
+ wpemod = 1
+ wpdiblc2 = 4.9866096e-9
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ poxedge = 1
+ tnoia = 0
+ binunit = 2
+ peta0 = 0
+ wketa = 6.9341182e-8
+ tnom = 25
+ tpbsw = 0.0025
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ cjswd = 5.1e-11
+ cjsws = 5.1e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ wkvth0we = 0.0
+ agidl = 3.2166e-9
+ tpbswg = 0.001
+ trnqsmod = 0
+ wags = -3.311005e-7
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ ptvoff = -4.0488554e-16
+ waigsd = 1.9105581e-12
+ voff = -0.13228318
+ acde = 0.5
+ scref = 1e-6
+ diomod = 1
+ vsat = 129757.01
+ pigcd = 2.572
+ rgatemod = 0
+ wint = 0
+ aigsd = 0.0063634264
+ vth0 = -0.39278391
+ tnjtsswg = 1
+ wkt1 = 1.4275631e-8
+ wkt2 = 2.8375299e-9
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.81e-10
+ pku0we = 0.0
+ wmax = 9e-7
+ wtvfbsdoff = 0
+ cjswgs = 1.81e-10
+ aigc = 0.0067852248
+ lvoff = 5.3109112e-9
+ wmin = 5.4e-7
+ ags = 1.1875295
+ tvfbsdoff = 0.1
+ )

.model pch_tt_20 pmos (
+ level = 54
+ cjd = 0.001346
+ cit = -0.00041212495
+ cjs = 0.001346
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ lvsat = 0
+ dlc = 1.38228675e-8
+ k3b = 2.1176
+ lvth0 = 6.5054743e-9
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ ltvfbsdoff = 0
+ wua1 = 2.4012676e-16
+ wub1 = -6.2487918e-26
+ delta = 0.018814
+ wuc1 = -3.9943707e-17
+ laigc = -2.2400472e-11
+ mjswgd = 0.95
+ mjswgs = 0.95
+ njtsswg = 6.489
+ bigc = 0.0012521
+ rnoia = 0
+ rnoib = 0
+ la0 = -7.2511148e-8
+ wwlc = 0
+ tcjswg = 0.00128
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0
+ kt1 = -0.20886849
+ kt2 = -0.049681978
+ lk2 = 1.2117426e-9
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ llc = -1.18e-13
+ lln = 0.7
+ lu0 = -4.8095715e-10
+ mjd = 0.335
+ mjs = 0.335
+ lua = -5.9775833e-17
+ lub = -8.2990392e-26
+ luc = -8.4878869e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = -2.0868237e-13
+ pketa = -1.8963071e-15
+ ckappad = 0.6
+ cdsc = 0
+ ckappas = 0.6
+ ngate = 1.7e+20
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ pk2 = -3.6576402e-16
+ pdiblc1 = 0
+ pdiblc2 = 0.01788848
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ ngcon = 1
+ xtis = 3
+ pdiblcb = 0
+ pu0 = -2.2283222e-17
+ wpclm = -5.08417e-8
+ prt = 0
+ pua = -3.7414239e-23
+ pub = 6.4271496e-32
+ puc = -3.5764571e-25
+ pud = 0
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigc = 0.15259
+ rsh = 15.2
+ wvfbsdoff = 0
+ tcj = 0.000832
+ ua1 = 1.3271195e-9
+ ub1 = -1.4620758e-18
+ uc1 = 1.6497662e-10
+ lvfbsdoff = 0
+ gbmin = 1e-12
+ tpb = 0.0016
+ wa0 = 8.4487289e-7
+ jswgd = 3.69e-13
+ ptvfbsdoff = 0
+ jswgs = 3.69e-13
+ ute = -1
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 1.4767164e-9
+ a0 = 1.2527531
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ wlc = 0
+ wln = 1
+ wu0 = 5.1646359e-10
+ at = 72000
+ cf = 8.17e-11
+ xgl = -8.2e-9
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.0030693202
+ xgw = 0
+ k3 = -2.5823
+ em = 20000000.0
+ wua = -8.6826164e-17
+ wub = 3.2435001e-26
+ wuc = -1.6113333e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ ll = -1.18e-13
+ lw = 0
+ u0 = 0.010136934
+ w0 = 0
+ ua = 5.8580479e-11
+ ub = 1.4664474e-18
+ uc = 4.9122952e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 6e-9
+ bigbacc = 0.0054401
+ fprout = 200
+ xrcrg1 = 12
+ xrcrg2 = 1
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ kvth0we = -0.00022
+ lintnoi = -5e-9
+ wtvoff = -3.604609e-11
+ bigbinv = 0.00149
+ k2we = 5e-5
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ dsub = 0.5
+ dtox = 3.91e-10
+ ijthsfwd = 0.01
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ tvoff = 0.0020688013
+ capmod = 2
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ wku0we = 1.5e-11
+ eta0 = 0.191845
+ etab = -0.18516667
+ mobmod = 0
+ ijthsrev = 0.01
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = 0
+ ppclm = 0
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ nfactor = 1
+ ppdiblc2 = 1.0915468e-15
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ nigbacc = 10
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ bigsd = 0.0003327
+ pkvth0we = 0.0
+ wvoff = -5.0330429e-9
+ nigbinv = 2.171
+ wvsat = -0.017628054
+ vfbsdoff = 0.01
+ wvth0 = 4.4926608e-9
+ keta = -0.023696099
+ waigc = -1.2459534e-12
+ lags = 6.5053339e-7
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 2.2533498e-10
+ toxref = 3e-9
+ paramchk = 1
+ lketa = -1.4702559e-8
+ kt1l = 0
+ xpart = 1
+ fnoimod = 1
+ eigbinv = 1.1
+ lint = 9.7879675e-9
+ egidl = 0.001
+ lkt1 = -1.3875579e-8
+ lkt2 = -5.3979298e-9
+ lmax = 4.4908e-7
+ lmin = 2.1577e-7
+ lpe0 = 6.44e-8
+ lpeb = 0
+ ijthdfwd = 0.01
+ ltvoff = -2.3926284e-10
+ minv = -0.33
+ lua1 = 4.9692128e-17
+ lub1 = -7.8826099e-26
+ luc1 = -1.8826114e-17
+ pvfbsdoff = 0
+ ndep = 1e+18
+ lwlc = 0
+ moin = 5.5538
+ cigbacc = 0.245
+ ijthdrev = 0.01
+ nigc = 2.291
+ lku0we = 1.8e-11
+ epsrox = 3.9
+ tnoimod = 0
+ lpdiblc2 = -2.233586e-9
+ pvoff = 1.1596021e-16
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ rdsmod = 0
+ cdscb = 0
+ cdscd = 0
+ cigbinv = 0.006
+ igbmod = 1
+ pvsat = 0
+ wk2we = 0.0
+ pvth0 = -1.7560727e-15
+ drout = 0.56
+ pags = 1.3163813e-13
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ paigc = -1.5565945e-18
+ ntox = 1
+ pcit = -2.0500564e-17
+ pclm = 1.2411167
+ pbswgd = 0.8
+ pbswgs = 0.8
+ voffl = 0
+ version = 4.5
+ igcmod = 1
+ phin = 0.15
+ tempmod = 0
+ weta0 = -2.432157e-8
+ wetab = 1.3741e-8
+ lkvth0we = 3e-12
+ lpclm = 0
+ pkt1 = 1.1573276e-15
+ pkt2 = 6.9635068e-17
+ aigbacc = 0.012071
+ cgidl = 1
+ acnqsmod = 0
+ rbdb = 50
+ pua1 = -2.8450432e-23
+ prwb = 0
+ pub1 = -5.1585101e-32
+ prwg = 0
+ puc1 = 1.7937993e-23
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ rdsw = 200
+ rbodymod = 0
+ pbswd = 0.9
+ pbsws = 0.9
+ aigbinv = 0.009974
+ permod = 1
+ pdits = 0
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ rshg = 14.1
+ voffcv = -0.125
+ wpemod = 1
+ wpdiblc2 = -3.6871397e-9
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ poxedge = 1
+ tnoia = 0
+ binunit = 2
+ peta0 = 0
+ wketa = 8.8109206e-9
+ tnom = 25
+ tpbsw = 0.0025
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ cjswd = 5.1e-11
+ cjsws = 5.1e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ wkvth0we = 0.0
+ agidl = 3.2166e-9
+ tpbswg = 0.001
+ trnqsmod = 0
+ wags = -5.9122303e-8
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ ptvoff = 4.9847489e-17
+ wcit = 4.6592191e-11
+ waigsd = 1.9150694e-12
+ voff = -0.10909205
+ acde = 0.5
+ scref = 1e-6
+ diomod = 1
+ vsat = 129757.01
+ pigcd = 2.572
+ rgatemod = 0
+ wint = 0
+ aigsd = 0.0063634182
+ vth0 = -0.40794766
+ tnjtsswg = 1
+ wkt1 = 1.0972613e-9
+ wkt2 = -4.2805615e-9
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.81e-10
+ pku0we = 0.0
+ wmax = 9e-7
+ wtvfbsdoff = 0
+ cjswgs = 1.81e-10
+ aigc = 0.0067947526
+ lvoff = -4.893186e-9
+ wmin = 5.4e-7
+ ags = -0.10644665
+ tvfbsdoff = 0.1
+ )

.model pch_tt_21 pmos (
+ level = 54
+ rbodymod = 0
+ version = 4.5
+ tempmod = 0
+ keta = -0.074839654
+ pvoff = 2.797289e-16
+ cdscb = 0
+ cdscd = 0
+ lags = 2.5597727e-7
+ pvsat = 0
+ aigbacc = 0.012071
+ wk2we = 0.0
+ pvth0 = 4.2710494e-16
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ drout = 0.56
+ fprout = 200
+ lcit = 1.4712816e-10
+ kt1l = 0
+ paigc = 3.3660127e-18
+ xrcrg1 = 12
+ xrcrg2 = 1
+ voffl = 0
+ wpdiblc2 = 2.1803424e-9
+ lint = 9.7879675e-9
+ weta0 = -2.432157e-8
+ wtvoff = -4.3702924e-10
+ aigbinv = 0.009974
+ wetab = 1.3741e-8
+ lkt1 = -6.1643471e-9
+ lkt2 = -3.8990903e-9
+ lmax = 2.1577e-7
+ lpclm = 5.4900145e-8
+ lmin = 9e-8
+ lpe0 = 6.44e-8
+ lpeb = 0
+ cgidl = 1
+ minv = -0.33
+ capmod = 2
+ lua1 = -2.9544713e-16
+ lub1 = 3.7855773e-25
+ luc1 = 4.6029572e-17
+ wku0we = 1.5e-11
+ a0 = 0.98313605
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ ndep = 1e+18
+ at = 41320.114
+ cf = 8.17e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.016096302
+ k3 = -2.5823
+ em = 20000000.0
+ ll = -1.18e-13
+ lwlc = 0
+ lw = 0
+ u0 = 0.008686993
+ mobmod = 0
+ w0 = 0
+ wkvth0we = 0.0
+ ua = 2.7312462e-10
+ ub = 6.1180894e-19
+ uc = 6.0007215e-11
+ ud = 0
+ moin = 5.5538
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 6e-9
+ pbswd = 0.9
+ pbsws = 0.9
+ nigc = 2.291
+ trnqsmod = 0
+ poxedge = 1
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ binunit = 2
+ pdits = 0
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ pags = -1.3976359e-13
+ ntox = 1
+ pcit = -3.638512e-17
+ pclm = 0.98092641
+ rgatemod = 0
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ tnjtsswg = 1
+ phin = 0.15
+ pkt1 = 1.542035e-15
+ pkt2 = 2.2793112e-15
+ tnoia = 0
+ peta0 = 0
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ wketa = -2.2984762e-8
+ tpbsw = 0.0025
+ rbdb = 50
+ pua1 = 7.9342593e-23
+ prwb = 0
+ pub1 = -9.194958e-32
+ prwg = 0
+ puc1 = -2.9723056e-23
+ cjswd = 5.1e-11
+ cjsws = 5.1e-11
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ mjswd = 0.01
+ rbsb = 50
+ pvag = 2.1
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ rdsw = 200
+ toxref = 3e-9
+ njtsswg = 6.489
+ ags = 1.7634876
+ scref = 1e-6
+ rshg = 14.1
+ cjd = 0.001346
+ cit = -4.1476524e-5
+ cjs = 0.001346
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ xtsswgd = 0.32
+ pigcd = 2.572
+ xtsswgs = 0.32
+ dlc = 1.38228675e-8
+ aigsd = 0.0063634182
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ tvfbsdoff = 0.1
+ ckappad = 0.6
+ ckappas = 0.6
+ lvoff = -2.4249846e-9
+ pdiblc1 = 0
+ pdiblc2 = 0.011594472
+ pdiblcb = 0
+ la0 = -1.5621959e-8
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0.006473456
+ lvsat = 0
+ kt1 = -0.24541461
+ kt2 = -0.056785482
+ lk2 = 3.9604228e-9
+ llc = -1.18e-13
+ lvth0 = 3.9839767e-9
+ lln = 0.7
+ ltvoff = -2.3342435e-10
+ lu0 = -1.7501951e-10
+ mjd = 0.335
+ mjs = 0.335
+ lua = -1.0504465e-16
+ ijthsfwd = 0.01
+ lub = 9.7338322e-26
+ luc = -1.0784466e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ delta = 0.018814
+ pa0 = -2.5809676e-14
+ nsd = 1e+20
+ laigc = -2.5435198e-11
+ pbd = 0.75
+ pat = -8.1994638e-9
+ pbs = 0.75
+ pk2 = 1.2451684e-16
+ tnom = 25
+ pu0 = -7.9199366e-18
+ prt = 0
+ pua = 5.00917e-23
+ pub = -8.1076857e-32
+ puc = 8.6464743e-24
+ pud = 0
+ rnoia = 0
+ rnoib = 0
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 2.9628506e-9
+ ub1 = -3.6297717e-18
+ uc1 = -1.423963e-10
+ bigbacc = 0.0054401
+ tpb = 0.0016
+ wa0 = -2.1822352e-8
+ pketa = 4.8125819e-15
+ ute = -1
+ wat = 0.038860018
+ ngate = 1.7e+20
+ web = 6628.3
+ wec = -16935.0
+ lku0we = 1.8e-11
+ wk2 = -8.468563e-10
+ wlc = 0
+ wln = 1
+ ijthsrev = 0.01
+ wu0 = 4.4839114e-10
+ xgl = -8.2e-9
+ ngcon = 1
+ xgw = 0
+ epsrox = 3.9
+ wua = -5.0154626e-16
+ wub = 7.2128975e-25
+ wuc = -5.8786887e-17
+ wud = 0
+ wpclm = 1.8489068e-7
+ wwc = 0
+ kvth0we = -0.00022
+ wwl = 0
+ wwn = 1
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ gbmin = 1e-12
+ lintnoi = -5e-9
+ rdsmod = 0
+ jswgd = 3.69e-13
+ bigbinv = 0.00149
+ jswgs = 3.69e-13
+ wags = 1.2271418e-6
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ igbmod = 1
+ wcit = 1.2187445e-10
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ voff = -0.12078969
+ acde = 0.5
+ pbswgd = 0.8
+ pbswgs = 0.8
+ ppdiblc2 = -1.4649193e-16
+ vsat = 129757.01
+ wint = 0
+ vth0 = -0.39599743
+ igcmod = 1
+ wkt1 = -7.259963e-10
+ wkt2 = -1.475296e-8
+ wmax = 9e-7
+ aigc = 0.0068091352
+ wmin = 5.4e-7
+ wua1 = -2.7074066e-16
+ wub1 = 1.2881293e-25
+ wuc1 = 1.8593804e-16
+ tvoff = 0.0020411307
+ bigc = 0.0012521
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ wwlc = 0
+ pkvth0we = 0.0
+ nfactor = 1
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ permod = 1
+ ku0we = -0.0007
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigc = 0.15259
+ beta0 = 13.32
+ vfbsdoff = 0.01
+ leta0 = 0
+ ppclm = -4.9739531e-14
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ nigbacc = 10
+ paramchk = 1
+ voffcv = -0.125
+ wpemod = 1
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ nigbinv = 2.171
+ k2we = 5e-5
+ dsub = 0.5
+ ijthdfwd = 0.01
+ dtox = 3.91e-10
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ bigsd = 0.0003327
+ eta0 = 0.191845
+ tpbswg = 0.001
+ etab = -0.18516667
+ wvoff = -5.8091978e-9
+ fnoimod = 1
+ ijthdrev = 0.01
+ eigbinv = 1.1
+ wvsat = -0.017628054
+ wvth0 = -5.8541529e-9
+ lpdiblc2 = -9.0555048e-10
+ wtvfbsdoff = 0
+ ptvoff = 1.3445493e-16
+ waigc = -2.4575845e-11
+ waigsd = 1.9150694e-12
+ ltvfbsdoff = 0
+ lketa = -3.9112692e-9
+ diomod = 1
+ xpart = 1
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.81e-10
+ pku0we = 0.0
+ cjswgs = 1.81e-10
+ cigbacc = 0.245
+ egidl = 0.001
+ lkvth0we = 3e-12
+ tnoimod = 0
+ mjswgd = 0.95
+ mjswgs = 0.95
+ cigbinv = 0.006
+ tcjswg = 0.00128
+ pvfbsdoff = 0
+ ptvfbsdoff = 0
+ acnqsmod = 0
+ )

.model pch_tt_22 pmos (
+ level = 54
+ xrcrg1 = 12
+ xrcrg2 = 1
+ paramchk = 1
+ rshg = 14.1
+ nfactor = 1
+ wtvoff = 2.0697628e-9
+ ijthdfwd = 0.01
+ capmod = 2
+ tvoff = -0.0031746364
+ tnom = 25
+ wku0we = 1.5e-11
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ mobmod = 0
+ nigbacc = 10
+ ijthdrev = 0.01
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = -1.0051895e-8
+ lpdiblc2 = 0
+ letab = 1.4778454e-8
+ nigbinv = 2.171
+ wags = -2.597049e-7
+ ppclm = 2.5985382e-14
+ wcit = -2.4970451e-10
+ dlcig = 2.5e-9
+ laigsd = 2.2969081e-18
+ bgidl = 1834800000.0
+ voff = -0.11952627
+ acde = 0.5
+ vsat = 226790.48
+ wint = 0
+ vth0 = -0.36144588
+ a0 = 2.9368155
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ wkt1 = -1.289882e-8
+ wkt2 = 2.7006409e-8
+ at = 192293.99
+ cf = 8.17e-11
+ wmax = 9e-7
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.02088367
+ k3 = -2.5823
+ em = 20000000.0
+ fnoimod = 1
+ aigc = 0.0066428307
+ wmin = 5.4e-7
+ ll = 0
+ lw = 0
+ u0 = 0.0082835417
+ dmcgt = 0
+ w0 = 0
+ ua = -1.5734149e-9
+ ub = 3.4167628e-18
+ uc = -1.3540772e-10
+ ud = 0
+ tcjsw = 9.34e-5
+ wl = 0
+ lkvth0we = 3e-12
+ wr = 1
+ xj = 1.1e-7
+ eigbinv = 1.1
+ xl = 4e-9
+ ww = 0
+ xw = 6e-9
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ wua1 = 6.2697239e-16
+ wub1 = -9.8389336e-25
+ wuc1 = -5.3295995e-16
+ bigc = 0.0012521
+ acnqsmod = 0
+ bigsd = 0.0003327
+ wwlc = 0
+ wvoff = -3.6240027e-9
+ cdsc = 0
+ rbodymod = 0
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigbacc = 0.245
+ wvsat = -0.072832829
+ cigc = 0.15259
+ wvth0 = 7.1065364e-9
+ waigc = 3.8715701e-11
+ tnoimod = 0
+ toxref = 3e-9
+ lketa = 1.7736502e-8
+ cigbinv = 0.006
+ xpart = 1
+ wpdiblc2 = 6.2191766e-10
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ egidl = 0.001
+ version = 4.5
+ ltvoff = 2.5685776e-10
+ k2we = 5e-5
+ tempmod = 0
+ dsub = 0.5
+ dtox = 3.91e-10
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ pvfbsdoff = 0
+ aigbacc = 0.012071
+ eta0 = 0.29878005
+ etab = -0.34238426
+ wkvth0we = 0.0
+ lku0we = 1.8e-11
+ epsrox = 3.9
+ trnqsmod = 0
+ rdsmod = 0
+ aigbinv = 0.009974
+ pvoff = 7.4320558e-17
+ igbmod = 1
+ cdscb = 0
+ cdscd = 0
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ pvsat = 5.1892488e-9
+ wk2we = 0.0
+ pvth0 = -7.9119985e-16
+ drout = 0.56
+ pbswgd = 0.8
+ pbswgs = 0.8
+ paigc = -2.5833927e-18
+ igcmod = 1
+ voffl = 0
+ rgatemod = 0
+ tnjtsswg = 1
+ weta0 = -7.0320749e-8
+ wetab = 2.4810139e-8
+ lpclm = -5.2812564e-8
+ poxedge = 1
+ cgidl = 1
+ binunit = 2
+ paigsd = -2.080997e-24
+ pbswd = 0.9
+ pbsws = 0.9
+ permod = 1
+ keta = -0.30513509
+ pdits = 0
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ jtsswgd = 1.75e-7
+ lcit = 1.1806861e-10
+ jtsswgs = 1.75e-7
+ voffcv = -0.125
+ wpemod = 1
+ kt1l = 0
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ lint = 0
+ lkt1 = -4.1189262e-9
+ lkt2 = 3.753071e-9
+ lmax = 9e-8
+ lmin = 5.4e-8
+ tnoia = 0
+ lpe0 = 6.44e-8
+ lpeb = 0
+ ijthsfwd = 0.01
+ peta0 = 4.3239229e-15
+ petab = -1.0404991e-15
+ wketa = 1.6222018e-7
+ minv = -0.33
+ wtvfbsdoff = 0
+ lua1 = 1.1693458e-16
+ lub1 = -2.0580342e-25
+ luc1 = -5.5456179e-17
+ tpbsw = 0.0025
+ tpbswg = 0.001
+ ndep = 1e+18
+ cjswd = 5.1e-11
+ njtsswg = 6.489
+ cjsws = 5.1e-11
+ mjswd = 0.01
+ lwlc = 0
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ moin = 5.5538
+ ltvfbsdoff = 0
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ ijthsrev = 0.01
+ nigc = 2.291
+ ckappad = 0.6
+ ckappas = 0.6
+ ags = 4.48665
+ pdiblc1 = 0
+ pdiblc2 = 0.0019609567
+ ptvoff = -1.0118352e-16
+ pdiblcb = 0
+ cjd = 0.001346
+ cit = 0.00026766759
+ waigsd = 1.9150916e-12
+ cjs = 0.001346
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ noff = 2.2684
+ bvs = 8.2
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ dlc = 4.0349e-9
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ diomod = 1
+ scref = 1e-6
+ ntox = 1
+ pcit = -1.4566987e-18
+ pclm = 2.1268063
+ la0 = -1.9926782e-7
+ pditsd = 0
+ pditsl = 0
+ ppdiblc2 = 0
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = -0.0077180887
+ cjswgd = 1.81e-10
+ pku0we = 0.0
+ pigcd = 2.572
+ kt1 = -0.26717441
+ cjswgs = 1.81e-10
+ kt2 = -0.13819145
+ lk2 = 4.4104354e-9
+ aigsd = 0.0063634181
+ bigbacc = 0.0054401
+ llc = 0
+ ptvfbsdoff = 0
+ lln = 1
+ lu0 = -1.3709508e-10
+ mjd = 0.335
+ mjs = 0.335
+ lua = 6.8530064e-17
+ lub = -1.6632734e-25
+ luc = 7.5845372e-18
+ lud = 0
+ tvfbsdoff = 0.1
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 2.4118768e-14
+ phin = 0.15
+ lvoff = -2.5437461e-9
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 2.0972465e-9
+ pbs = 0.75
+ pk2 = 2.0570947e-16
+ pu0 = 1.8416833e-16
+ kvth0we = -0.00022
+ prt = 0
+ pua = -1.7823119e-23
+ pub = 1.268951e-31
+ puc = -7.4643321e-24
+ pud = 0
+ pkt1 = 2.6862803e-15
+ pkt2 = -1.6460695e-15
+ lvsat = -0.009121146
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = -1.4241889e-9
+ ub1 = 2.5868363e-18
+ mjswgd = 0.95
+ lvth0 = 7.3613109e-10
+ uc1 = 9.3723935e-10
+ mjswgs = 0.95
+ lintnoi = -5e-9
+ tpb = 0.0016
+ wa0 = -5.5297601e-7
+ delta = 0.018814
+ bigbinv = 0.00149
+ ute = -1
+ vtsswgd = 1.1
+ wat = -0.070679454
+ laigc = -9.8025804e-12
+ vtsswgs = 1.1
+ tcjswg = 0.00128
+ web = 6628.3
+ wec = -16935.0
+ wk2 = -1.7106076e-9
+ wlc = 0
+ wln = 1
+ wu0 = -1.5951011e-9
+ xgl = -8.2e-9
+ xgw = 0
+ wua = 2.2095182e-16
+ wub = -1.4911779e-24
+ wuc = 1.1260467e-16
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ rnoia = 0
+ rnoib = 0
+ rbdb = 50
+ pua1 = -5.0424332e-24
+ prwb = 0
+ pub1 = 1.2644812e-32
+ prwg = 0
+ puc1 = 3.7853356e-23
+ pkvth0we = 0.0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ pketa = -1.2596682e-14
+ ngate = 1.7e+20
+ rdsw = 200
+ ngcon = 1
+ wvfbsdoff = 0
+ wpclm = -6.2069351e-7
+ lvfbsdoff = 0
+ vfbsdoff = 0.01
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ fprout = 200
+ )

.model pch_tt_23 pmos (
+ level = 54
+ ijthsfwd = 0.01
+ dtox = 3.91e-10
+ cgidl = 1
+ wku0we = 1.5e-11
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ mobmod = 0
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ eta0 = 7.956713e-6
+ etab = -0.26192508
+ pbswd = 0.9
+ pbsws = 0.9
+ ijthsrev = 0.01
+ pdits = 0
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ ppdiblc2 = 0
+ njtsswg = 6.489
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ tnoia = 0
+ ckappad = 0.6
+ ckappas = 0.6
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ pdiblc1 = 0
+ pdiblc2 = 0.0019609567
+ pdiblcb = 0
+ peta0 = -2.7992439e-15
+ petab = -1.6989745e-15
+ wketa = -4.2902456e-7
+ tpbsw = 0.0025
+ cjswd = 5.1e-11
+ cjsws = 5.1e-11
+ pkvth0we = 0.0
+ ags = 4.48665
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ cjd = 0.001346
+ cit = -0.002877963
+ cjs = 0.001346
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 4.0349e-9
+ bigbacc = 0.0054401
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ vfbsdoff = 0.01
+ a0 = 5.6551822
+ a1 = 0
+ a2 = 1
+ keta = 0.46798148
+ b0 = 0
+ b1 = 0
+ kvth0we = -0.00022
+ at = -40561.437
+ cf = 8.17e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.018874979
+ k3 = -2.5823
+ em = 20000000.0
+ la0 = -3.569331e-7
+ toxref = 3e-9
+ ll = 0
+ jsd = 1.5e-7
+ lw = 0
+ jss = 1.5e-7
+ lat = 0.0057875263
+ u0 = 0.0072884759
+ w0 = 0
+ kt1 = -0.46532049
+ kt2 = 0.0072316444
+ lk2 = 4.2939313e-9
+ ua = 5.3944309e-9
+ ub = -7.8004593e-18
+ uc = 1.0922891e-10
+ ud = 0
+ llc = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ lln = 1
+ xw = 6e-9
+ lu0 = -7.938127e-11
+ mjd = 0.335
+ lintnoi = -5e-9
+ mjs = 0.335
+ lua = -3.3560499e-16
+ lub = 4.8427154e-25
+ luc = -6.604387e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ bigbinv = 0.00149
+ njs = 1.02
+ pa0 = 1.517818e-13
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ nsd = 1e+20
+ lcit = 3.0051519e-10
+ pbd = 0.75
+ pat = -1.8496379e-9
+ pbs = 0.75
+ pk2 = 4.9657487e-16
+ paramchk = 1
+ pu0 = -8.1141216e-17
+ scref = 1e-6
+ kt1l = 0
+ prt = 0
+ pua = 1.7043409e-22
+ pub = -3.4061954e-31
+ puc = 5.8491101e-24
+ pud = 0
+ pigcd = 2.572
+ rsh = 15.2
+ aigsd = 0.0063634182
+ tcj = 0.000832
+ ua1 = 9.464156e-9
+ tvfbsdoff = 0.1
+ ub1 = -1.352433e-17
+ uc1 = -1.5339544e-9
+ tpb = 0.0016
+ wa0 = -2.7540628e-6
+ lint = 0
+ ute = -1
+ wat = -0.002629722
+ lvoff = -5.520199e-9
+ web = 6628.3
+ wec = -16935.0
+ wk2 = -6.7255282e-9
+ wlc = 0
+ wln = 1
+ lkt1 = 7.3735466e-9
+ lkt2 = -4.6814687e-9
+ wu0 = 2.9792015e-9
+ xgl = -8.2e-9
+ xgw = 0
+ ltvoff = -2.6406105e-10
+ wua = -3.0248621e-15
+ wub = 6.5694194e-24
+ wuc = -1.1693744e-16
+ wud = 0
+ lmax = 5.4e-8
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ lmin = 4.5e-8
+ lvsat = 0.0051141042
+ lpe0 = 6.44e-8
+ lvth0 = -6.7414368e-9
+ lpeb = 0
+ ijthdfwd = 0.01
+ delta = 0.018814
+ laigc = -1.6050622e-11
+ minv = -0.33
+ lua1 = -5.1458943e-16
+ lub1 = 7.2864421e-25
+ luc1 = 8.7873061e-17
+ rnoia = 0
+ rnoib = 0
+ ndep = 1e+18
+ lku0we = 1.8e-11
+ lwlc = 0
+ epsrox = 3.9
+ moin = 5.5538
+ pketa = 2.1695512e-14
+ ngate = 1.7e+20
+ wvfbsdoff = 0
+ ijthdrev = 0.01
+ lvfbsdoff = 0
+ ngcon = 1
+ nigc = 2.291
+ wpclm = -1.0386396e-6
+ nfactor = 1
+ rdsmod = 0
+ igbmod = 1
+ lpdiblc2 = 0
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ noff = 2.2684
+ pscbe1 = 926400000.0
+ noia = 2.86e+42
+ pscbe2 = 1e-20
+ noib = 2.5e+24
+ noic = 31000000000.0
+ pbswgd = 0.8
+ pbswgs = 0.8
+ igcmod = 1
+ ntox = 1
+ pcit = -4.3391024e-17
+ pclm = 4.4879115
+ nigbacc = 10
+ phin = 0.15
+ lkvth0we = 3e-12
+ pkt1 = -5.0612736e-15
+ pkt2 = 1.1767646e-15
+ nigbinv = 2.171
+ tvoff = 0.0058067224
+ acnqsmod = 0
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ rbdb = 50
+ pua1 = 2.7224008e-22
+ prwb = 0
+ pub1 = -3.6990718e-31
+ prwg = 0
+ puc1 = -5.7927018e-23
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ permod = 1
+ rbodymod = 0
+ rdsw = 200
+ ku0we = -0.0007
+ beta0 = 13.32
+ fnoimod = 1
+ leta0 = 7.2768866e-9
+ letab = 1.0111821e-8
+ eigbinv = 1.1
+ ppclm = 5.0226256e-14
+ voffcv = -0.125
+ wpemod = 1
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ rshg = 14.1
+ wtvfbsdoff = 0
+ wpdiblc2 = 6.2191766e-10
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ ltvfbsdoff = 0
+ cigbacc = 0.245
+ tnoimod = 0
+ tnom = 25
+ tpbswg = 0.001
+ bigsd = 0.0003327
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ cigbinv = 0.006
+ wkvth0we = 0.0
+ wvoff = -2.1208799e-8
+ trnqsmod = 0
+ wvsat = 0.09105966
+ ptvoff = 1.2747838e-16
+ ptvfbsdoff = 0
+ wvth0 = -3.7395008e-8
+ waigsd = 1.9150557e-12
+ version = 4.5
+ waigc = -1.4751759e-11
+ wags = -2.597049e-7
+ tempmod = 0
+ wcit = 4.7330111e-10
+ diomod = 1
+ voff = -0.068208113
+ lketa = -2.7104259e-8
+ acde = 0.5
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.81e-10
+ pku0we = 0.0
+ cjswgs = 1.81e-10
+ aigbacc = 0.012071
+ xpart = 1
+ rgatemod = 0
+ vsat = -18644.867
+ wint = 0
+ vth0 = -0.2325223
+ tnjtsswg = 1
+ wkt1 = 1.206797e-7
+ wkt2 = -2.1663145e-8
+ egidl = 0.001
+ wmax = 9e-7
+ aigc = 0.0067505556
+ wmin = 5.4e-7
+ mjswgd = 0.95
+ mjswgs = 0.95
+ aigbinv = 0.009974
+ tcjswg = 0.00128
+ pvfbsdoff = 0
+ wua1 = -4.1537606e-15
+ wub1 = 5.6118307e-24
+ wuc1 = 1.1184258e-15
+ bigc = 0.0012521
+ wwlc = 0
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigc = 0.15259
+ pvoff = 1.0942388e-15
+ poxedge = 1
+ cdscb = 0
+ cdscd = 0
+ fprout = 200
+ pvsat = -4.3165155e-9
+ wk2we = 0.0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ pvth0 = 1.7898897e-15
+ drout = 0.56
+ binunit = 2
+ paigc = 5.1772001e-19
+ voffl = 0
+ dmcg = 3.1e-8
+ wtvoff = -1.8726837e-9
+ dmci = 3.1e-8
+ dmdg = 0
+ weta0 = 5.2492471e-8
+ wetab = 3.6163164e-8
+ lpclm = -1.8975667e-7
+ k2we = 5e-5
+ capmod = 2
+ dsub = 0.5
+ )

.model pch_tt_24 pmos (
+ level = 54
+ beta0 = 13.32
+ leta0 = 4.5580824e-10
+ letab = 2.8639817e-9
+ cigbacc = 0.245
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ ppclm = -6.983762e-15
+ laigsd = -1.7489044e-14
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ tnoimod = 0
+ ntox = 1
+ pcit = -2.3939875e-16
+ pclm = 0.55996802
+ rgatemod = 0
+ cigbinv = 0.006
+ tnjtsswg = 1
+ phin = 0.15
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ pkt1 = 8.0439909e-15
+ pkt2 = -6.3201272e-16
+ version = 4.5
+ tempmod = 0
+ bigsd = 0.0003327
+ rbdb = 50
+ pua1 = -2.7866327e-22
+ prwb = 0
+ pub1 = 3.2786288e-31
+ prwg = 0
+ puc1 = 2.5974765e-23
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ aigbacc = 0.012071
+ wvoff = -2.6959456e-8
+ rdsw = 200
+ wvsat = 0.037826603
+ wvth0 = -5.1175681e-9
+ toxref = 3e-9
+ waigc = -9.7737582e-11
+ aigbinv = 0.009974
+ lketa = 1.4220453e-8
+ rshg = 14.1
+ xpart = 1
+ egidl = 0.001
+ ltvoff = -2.5344658e-10
+ pvfbsdoff = 0
+ ijthsfwd = 0.01
+ poxedge = 1
+ a0 = -2.5402778
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ tnom = 25
+ at = 213109.93
+ cf = 8.17e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.022656115
+ k3 = -2.5823
+ em = 20000000.0
+ lku0we = 1.8e-11
+ ll = 0
+ lw = 0
+ u0 = 0.0013978574
+ w0 = 0
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ ua = -6.0379704e-9
+ ub = 8.1069989e-18
+ uc = -2.2784413e-10
+ ud = 0
+ binunit = 2
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ epsrox = 3.9
+ xw = 6e-9
+ ijthsrev = 0.01
+ rdsmod = 0
+ igbmod = 1
+ pvoff = 1.376021e-15
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ wags = -2.597049e-7
+ cdscb = 0
+ cdscd = 0
+ pbswgd = 0.8
+ pbswgs = 0.8
+ pvsat = -1.7080957e-9
+ wcit = 4.4734589e-9
+ wk2we = 0.0
+ pvth0 = 2.0829517e-16
+ drout = 0.56
+ igcmod = 1
+ voff = -0.080254273
+ paigc = 4.5840253e-18
+ acde = 0.5
+ ppdiblc2 = 0
+ voffl = 0
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ vsat = 78763.66
+ wint = 0
+ vth0 = -0.35515952
+ wkt1 = -1.4677468e-7
+ wkt2 = 1.5250678e-8
+ wmax = 9e-7
+ weta0 = -2.1233528e-8
+ aigc = 0.0066531108
+ wetab = 8.325777e-9
+ wmin = 5.4e-7
+ lpclm = 2.7125638e-9
+ cgidl = 1
+ paigsd = 9.5490179e-21
+ wua1 = 7.089165e-15
+ wub1 = -8.6283747e-24
+ wuc1 = -5.9385548e-16
+ bigc = 0.0012521
+ wwlc = 0
+ pkvth0we = 0.0
+ permod = 1
+ cdsc = 0
+ pbswd = 0.9
+ pbsws = 0.9
+ njtsswg = 6.489
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ wtvfbsdoff = 0
+ cigc = 0.15259
+ vfbsdoff = 0.01
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ ckappad = 0.6
+ ckappas = 0.6
+ pdits = 0
+ voffcv = -0.125
+ wpemod = 1
+ pdiblc1 = 0
+ pdiblc2 = 0.0019609567
+ cigsd = 0.013281
+ ltvfbsdoff = 0
+ pdiblcb = 0
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ paramchk = 1
+ pk2we = 0.0
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ bigbacc = 0.0054401
+ tnoia = 0
+ k2we = 5e-5
+ ags = 4.48665
+ ijthdfwd = 0.01
+ dsub = 0.5
+ dtox = 3.91e-10
+ kvth0we = -0.00022
+ peta0 = 8.1333004e-16
+ ptvfbsdoff = 0
+ petab = -3.349425e-16
+ cjd = 0.001346
+ cit = -0.010137593
+ cjs = 0.001346
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dvt0 = 3.48
+ tpbswg = 0.001
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ wketa = 1.6324308e-7
+ dlc = 4.0349e-9
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ tpbsw = 0.0025
+ dwg = 0
+ lintnoi = -5e-9
+ dwj = 0
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ cjswd = 5.1e-11
+ cjsws = 5.1e-11
+ mjswd = 0.01
+ eta0 = 0.13921364
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ etab = -0.11400999
+ la0 = 4.4644444e-8
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = -0.0066423707
+ kt1 = 0.16833478
+ kt2 = -0.11193164
+ lk2 = 4.479207e-9
+ ijthdrev = 0.01
+ llc = 0
+ lln = 1
+ lu0 = 2.0925904e-10
+ mjd = 0.335
+ ptvoff = 8.5019581e-17
+ mjs = 0.335
+ lua = 2.2458267e-16
+ lub = -2.9519392e-25
+ luc = 9.9121919e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = -8.9774533e-14
+ waigsd = 1.7201778e-12
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 6.8793549e-9
+ pbs = 0.75
+ lpdiblc2 = 0
+ pk2 = 1.0702031e-16
+ pu0 = -9.6657248e-17
+ prt = 0
+ pua = -9.0705467e-23
+ pub = 1.0841652e-31
+ puc = -1.0416838e-23
+ pud = 0
+ diomod = 1
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = -1.018181e-8
+ ub1 = 1.2390462e-17
+ uc1 = 9.111363e-10
+ tpb = 0.0016
+ wa0 = 2.1756583e-6
+ ute = -1
+ wat = -0.18077244
+ pditsd = 0
+ web = 6628.3
+ wec = -16935.0
+ pditsl = 0
+ wk2 = 1.2245648e-9
+ cjswgd = 1.81e-10
+ pku0we = 0.0
+ cjswgs = 1.81e-10
+ wlc = 0
+ wln = 1
+ wu0 = 3.2958552e-9
+ xgl = -8.2e-9
+ xgw = 0
+ scref = 1e-6
+ wua = 2.3045166e-15
+ wub = -2.5945817e-24
+ wuc = 2.150207e-16
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ tvfbsdoff = 0.1
+ pigcd = 2.572
+ aigsd = 0.0063637751
+ lvoff = -4.9299372e-9
+ mjswgd = 0.95
+ mjswgs = 0.95
+ lkvth0we = 3e-12
+ nfactor = 1
+ lvsat = 0.00034108628
+ tcjswg = 0.00128
+ lvth0 = -7.3221299e-10
+ delta = 0.018814
+ laigc = -1.1275829e-11
+ acnqsmod = 0
+ rnoia = 0
+ rnoib = 0
+ wvfbsdoff = 0
+ pketa = -7.3256019e-15
+ ngate = 1.7e+20
+ lvfbsdoff = 0
+ rbodymod = 0
+ nigbacc = 10
+ ngcon = 1
+ wpclm = 1.2891178e-7
+ gbmin = 1e-12
+ keta = -0.37538
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ fprout = 200
+ xrcrg1 = 12
+ xrcrg2 = 1
+ nigbinv = 2.171
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 6.5623704e-10
+ kt1l = 0
+ wtvoff = -1.0061777e-9
+ wpdiblc2 = 6.2191766e-10
+ lint = 0
+ lkt1 = -2.3675561e-8
+ lkt2 = 1.1575324e-9
+ lmax = 4.5e-8
+ lmin = 3.6e-8
+ capmod = 2
+ fnoimod = 1
+ lpe0 = 6.44e-8
+ lpeb = 0
+ wku0we = 1.5e-11
+ eigbinv = 1.1
+ tvoff = 0.0055901005
+ mobmod = 0
+ minv = -0.33
+ lua1 = 4.4806289e-16
+ lub1 = -5.4118058e-25
+ luc1 = -3.1936385e-17
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ ndep = 1e+18
+ wkvth0we = 0.0
+ lwlc = 0
+ moin = 5.5538
+ nigc = 2.291
+ trnqsmod = 0
+ ku0we = -0.0007
+ )

.model pch_tt_25 pmos (
+ level = 54
+ wint = 0
+ ags = 0.93810347
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ vth0 = -0.37798248
+ wkt1 = -1.5318394e-9
+ wkt2 = 2.21858e-9
+ cjd = 0.001346
+ cit = 5e-6
+ cjs = 0.001346
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ wmax = 5.4e-7
+ bvs = 8.2
+ aigc = 0.0068215676
+ wmin = 2.7e-7
+ dlc = 1.0572421799999999e-8
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ k3b = 2.1176
+ lkvth0we = 3e-12
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ tnoia = 0
+ peta0 = 0
+ la0 = 0
+ wua1 = 1.6452204e-16
+ wub1 = -6.9710259e-26
+ wuc1 = 2.1709154e-17
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0
+ wketa = 2.2687563e-8
+ kt1 = -0.17747938
+ lk2 = 0
+ kt2 = -0.061438333
+ llc = 0
+ lln = 1
+ lu0 = 0
+ tpbsw = 0.0025
+ acnqsmod = 0
+ mjd = 0.335
+ bigc = 0.0012521
+ mjs = 0.335
+ wute = 3.2371733e-8
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ wwlc = 0
+ pa0 = 0
+ cjswd = 5.1e-11
+ nsd = 1e+20
+ cjsws = 5.1e-11
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ pk2 = 0
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ pu0 = 0
+ prt = 0
+ pud = 0
+ rbodymod = 0
+ cdsc = 0
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 1.8507467e-10
+ ub1 = -1.7337534e-19
+ uc1 = -4.0886356e-11
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ tpb = 0.0016
+ wa0 = -1.5013787e-7
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigc = 0.15259
+ ute = -1.2102889
+ toxref = 3e-9
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 4.440518e-10
+ wlc = 0
+ wln = 1
+ wu0 = 3.7953067e-11
+ xgl = -8.2e-9
+ xgw = 0
+ nfactor = 1
+ wua = -1.5196107e-16
+ wub = 9.0507286e-26
+ wuc = 5.3799588e-18
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ scref = 1e-6
+ tvfbsdoff = 0.1
+ pigcd = 2.572
+ aigsd = 0.0063632886
+ wpdiblc2 = -7.7579138e-11
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ ltvoff = 0
+ lvoff = 0
+ nigbacc = 10
+ lvsat = 0
+ k2we = 5e-5
+ lvth0 = 0
+ dsub = 0.5
+ dtox = 3.91e-10
+ delta = 0.018814
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ lku0we = 1.8e-11
+ rnoia = 0
+ rnoib = 0
+ epsrox = 3.9
+ nigbinv = 2.171
+ eta0 = 0.17962267
+ wvfbsdoff = 0
+ wkvth0we = 0.0
+ etab = -0.19577778
+ lvfbsdoff = 0
+ ngate = 1.7e+20
+ rdsmod = 0
+ ngcon = 1
+ igbmod = 1
+ wpclm = -1.1447315e-8
+ trnqsmod = 0
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ pbswgd = 0.8
+ pbswgs = 0.8
+ fnoimod = 1
+ eigbinv = 1.1
+ igcmod = 1
+ a0 = 3.3089778
+ a1 = 0
+ a2 = 1
+ rgatemod = 0
+ b0 = 0
+ b1 = 0
+ at = 72000
+ cf = 8.17e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.0028441163
+ k3 = -2.5823
+ em = 20000000.0
+ tnjtsswg = 1
+ ll = 0
+ lw = 0
+ u0 = 0.0096414889
+ w0 = 0
+ ua = 1.8228697e-10
+ ub = 9.7616315e-19
+ uc = -9.1826044e-12
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 6e-9
+ wtvfbsdoff = 0
+ cigbacc = 0.245
+ tvoff = 0.0026578776
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ permod = 1
+ ltvfbsdoff = 0
+ tnoimod = 0
+ cigbinv = 0.006
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = 0
+ keta = -0.064397096
+ voffcv = -0.125
+ wpemod = 1
+ ppclm = 0
+ version = 4.5
+ dlcig = 2.5e-9
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ bgidl = 1834800000.0
+ lcit = 0
+ tempmod = 0
+ ptvfbsdoff = 0
+ kt1l = 0
+ aigbacc = 0.012071
+ lint = 6.5375218e-9
+ dmcgt = 0
+ lkt1 = 0
+ tcjsw = 9.34e-5
+ lmax = 2.001e-5
+ lmin = 8.9991e-6
+ lpe0 = 6.44e-8
+ lpeb = 0
+ ijthsfwd = 0.01
+ tpbswg = 0.001
+ minv = -0.33
+ aigbinv = 0.009974
+ bigsd = 0.0003327
+ ndep = 1e+18
+ lwlc = 0
+ moin = 5.5538
+ wvoff = 2.5521431e-9
+ ptvoff = 0
+ ijthsrev = 0.01
+ nigc = 2.291
+ waigsd = 1.9763167e-12
+ wvsat = 0.0034765009
+ wvth0 = -1.8147147e-9
+ diomod = 1
+ waigc = 4.045116e-12
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.81e-10
+ pku0we = 0.0
+ cjswgs = 1.81e-10
+ poxedge = 1
+ lketa = 0
+ ntox = 1
+ xpart = 1
+ pcit = 0
+ pclm = 1.1689658
+ ppdiblc2 = 0
+ binunit = 2
+ egidl = 0.001
+ mjswgd = 0.95
+ mjswgs = 0.95
+ phin = 0.15
+ tcjswg = 0.00128
+ pkt1 = 0
+ pvfbsdoff = 0
+ rbdb = 50
+ prwb = 0
+ prwg = 0
+ pkvth0we = 0.0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ jtsswgd = 1.75e-7
+ rdsw = 200
+ jtsswgs = 1.75e-7
+ vfbsdoff = 0.01
+ fprout = 200
+ pvoff = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ cdscb = 0
+ cdscd = 0
+ pvsat = 0
+ wk2we = 0.0
+ pvth0 = 0
+ drout = 0.56
+ paramchk = 1
+ wtvoff = -1.0551434e-10
+ rshg = 14.1
+ voffl = 0
+ weta0 = -1.7648176e-8
+ wetab = 1.9534667e-8
+ njtsswg = 6.489
+ capmod = 2
+ lpclm = 0
+ wku0we = 1.5e-11
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ ijthdfwd = 0.01
+ cgidl = 1
+ mobmod = 0
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.0030491463
+ tnom = 25
+ pdiblcb = 0
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ pbswd = 0.9
+ pbsws = 0.9
+ ijthdrev = 0.01
+ lpdiblc2 = 0
+ bigbacc = 0.0054401
+ wags = -6.1953916e-9
+ pdits = 0
+ cigsd = 0.013281
+ kvth0we = -0.00022
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ voff = -0.10784306
+ acde = 0.5
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ vsat = 91103.982
+ pk2we = 0.0
+ )

.model pch_tt_26 pmos (
+ level = 54
+ bigsd = 0.0003327
+ poxedge = 1
+ pkvth0we = 0.0
+ wvoff = 2.9007224e-9
+ binunit = 2
+ toxref = 3e-9
+ wvsat = 0.0034765009
+ wvth0 = -1.8762892e-9
+ vfbsdoff = 0.01
+ keta = -0.06875265
+ waigc = 4.3476029e-12
+ lags = 1.0877241e-7
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 0
+ lketa = 3.9156432e-8
+ paramchk = 1
+ kt1l = 0
+ xpart = 1
+ ltvoff = -4.4286369e-10
+ egidl = 0.001
+ lint = 6.5375218e-9
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ lkt1 = -3.4853729e-8
+ lkt2 = -1.4641311e-8
+ lmax = 8.9991e-6
+ pvfbsdoff = 0
+ lmin = 8.9908e-7
+ lpe0 = 6.44e-8
+ ijthdfwd = 0.01
+ lpeb = 0
+ lku0we = 1.8e-11
+ minv = -0.33
+ epsrox = 3.9
+ lua1 = 1.4818924e-15
+ lub1 = -2.0711788e-24
+ luc1 = 2.2491171e-16
+ ndep = 1e+18
+ lute = 1.330224e-7
+ rdsmod = 0
+ lwlc = 0
+ moin = 5.5538
+ igbmod = 1
+ ijthdrev = 0.01
+ nigc = 2.291
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ lpdiblc2 = 8.2033961e-9
+ njtsswg = 6.489
+ pbswgd = 0.8
+ pvoff = -3.1337282e-15
+ pbswgs = 0.8
+ noff = 2.2684
+ cdscb = 0
+ cdscd = 0
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ igcmod = 1
+ pvsat = 0
+ wk2we = 0.0
+ pvth0 = 5.5355474e-16
+ drout = 0.56
+ ckappad = 0.6
+ ckappas = 0.6
+ pags = 8.2314292e-14
+ wtvfbsdoff = 0
+ pdiblc1 = 0
+ pdiblc2 = 0.002136644
+ paigc = -2.7193569e-18
+ pdiblcb = 0
+ ntox = 1
+ pcit = 0
+ pclm = 1.1689658
+ voffl = 0
+ ltvfbsdoff = 0
+ weta0 = -1.7648176e-8
+ phin = 0.15
+ wetab = 1.9534667e-8
+ lkvth0we = 3e-12
+ lpclm = 0
+ paigsd = -4.5957918e-20
+ pkt1 = 4.5592526e-15
+ pkt2 = 3.8774237e-15
+ bigbacc = 0.0054401
+ cgidl = 1
+ permod = 1
+ acnqsmod = 0
+ kvth0we = -0.00022
+ rbdb = 50
+ pua1 = -9.4343892e-23
+ prwb = 0
+ pub1 = 9.0084871e-32
+ prwg = 0
+ puc1 = -7.238167e-23
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ lintnoi = -5e-9
+ pute = -1.6539558e-14
+ bigbinv = 0.00149
+ rbodymod = 0
+ pbswd = 0.9
+ pbsws = 0.9
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ rdsw = 200
+ ptvfbsdoff = 0
+ a0 = 3.4253346
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 72000
+ cf = 8.17e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.0024652651
+ k3 = -2.5823
+ em = 20000000.0
+ ll = 0
+ voffcv = -0.125
+ lw = 0
+ wpemod = 1
+ u0 = 0.0095254275
+ w0 = 0
+ ua = 1.8429003e-10
+ ub = 9.3982253e-19
+ uc = -1.1498405e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 6e-9
+ pdits = 0
+ cigsd = 0.013281
+ ags = 0.9260042
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ cjd = 0.001346
+ cit = 5e-6
+ cjs = 0.001346
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 1.0572421799999999e-8
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ rshg = 14.1
+ wpdiblc2 = 3.818702e-12
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ la0 = -1.0460478e-6
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0
+ kt1 = -0.17360244
+ kt2 = -0.059809712
+ lk2 = -3.4058721e-9
+ llc = 0
+ lln = 1
+ lu0 = 1.0433917e-9
+ mjd = 0.335
+ mjs = 0.335
+ lua = -1.8007487e-17
+ lub = 3.2670219e-25
+ luc = 2.0819042e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ tnoia = 0
+ njd = 1.02
+ njs = 1.02
+ pa0 = 1.483047e-13
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ tpbswg = 0.001
+ pk2 = 2.5596912e-15
+ pu0 = 1.7642195e-17
+ nfactor = 1
+ peta0 = 0
+ prt = 0
+ pua = 1.2819791e-23
+ pub = -1.2787603e-32
+ puc = -1.6865938e-24
+ pud = 0
+ wketa = 2.5468383e-8
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 2.0236805e-11
+ ub1 = 5.7011626e-20
+ uc1 = -6.5904343e-11
+ tnom = 25
+ tpbsw = 0.0025
+ tpb = 0.0016
+ wa0 = -1.666345e-7
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ ute = -1.2250856
+ cjswd = 5.1e-11
+ cjsws = 5.1e-11
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 1.5932531e-10
+ mjswd = 0.01
+ wlc = 0
+ mjsws = 0.01
+ wln = 1
+ agidl = 3.2166e-9
+ wu0 = 3.5990642e-11
+ wkvth0we = 0.0
+ xgl = -8.2e-9
+ xgw = 0
+ wua = -1.5338707e-16
+ wub = 9.1929712e-26
+ wuc = 5.5675666e-18
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ ptvoff = -2.4168192e-17
+ waigsd = 1.9814288e-12
+ trnqsmod = 0
+ nigbacc = 10
+ diomod = 1
+ wags = -1.5351598e-8
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.81e-10
+ pku0we = 0.0
+ cjswgs = 1.81e-10
+ tvfbsdoff = 0.1
+ voff = -0.10676035
+ scref = 1e-6
+ acde = 0.5
+ nigbinv = 2.171
+ pigcd = 2.572
+ rgatemod = 0
+ aigsd = 0.0063632773
+ vsat = 91103.982
+ wint = 0
+ vth0 = -0.37656355
+ tnjtsswg = 1
+ mjswgd = 0.95
+ mjswgs = 0.95
+ wkt1 = -2.0389865e-9
+ wkt2 = 1.7872759e-9
+ lvoff = -9.7335308e-9
+ wmax = 5.4e-7
+ aigc = 0.0068257672
+ wmin = 2.7e-7
+ tcjswg = 0.00128
+ lvsat = 0
+ lvth0 = -1.2756137e-8
+ delta = 0.018814
+ laigc = -3.7754415e-11
+ wua1 = 1.7501635e-16
+ wub1 = -7.9730823e-26
+ wuc1 = 2.9760508e-17
+ fnoimod = 1
+ rnoia = 0
+ rnoib = 0
+ bigc = 0.0012521
+ eigbinv = 1.1
+ wute = 3.4211506e-8
+ wwlc = 0
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ pketa = -2.4999571e-14
+ ngate = 1.7e+20
+ cdsc = 0
+ ngcon = 1
+ cgbo = 0
+ wpclm = -1.1447315e-8
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ fprout = 200
+ cigc = 0.15259
+ gbmin = 1e-12
+ xrcrg1 = 12
+ xrcrg2 = 1
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ cigbacc = 0.245
+ wtvoff = -1.02826e-10
+ tnoimod = 0
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ capmod = 2
+ cigbinv = 0.006
+ wku0we = 1.5e-11
+ k2we = 5e-5
+ mobmod = 0
+ ijthsfwd = 0.01
+ dsub = 0.5
+ dtox = 3.91e-10
+ tvoff = 0.0027071394
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ xjbvd = 1
+ xjbvs = 1
+ version = 4.5
+ lk2we = 0.0
+ tempmod = 0
+ eta0 = 0.17962267
+ etab = -0.19577778
+ ijthsrev = 0.01
+ ku0we = -0.0007
+ aigbacc = 0.012071
+ beta0 = 13.32
+ leta0 = 0
+ laigsd = 1.0132005e-13
+ ppclm = 0
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ aigbinv = 0.009974
+ ppdiblc2 = -7.3176658e-16
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ )

.model pch_tt_27 pmos (
+ level = 54
+ tvfbsdoff = 0.1
+ fnoimod = 1
+ scref = 1e-6
+ eigbinv = 1.1
+ rshg = 14.1
+ ltvoff = -3.7535707e-10
+ pigcd = 2.572
+ aigsd = 0.0063633912
+ lvoff = -1.1639377e-8
+ lvsat = 0
+ lvth0 = 1.0506701e-9
+ ijthsfwd = 0.01
+ lku0we = 1.8e-11
+ delta = 0.018814
+ laigc = -5.5983746e-11
+ epsrox = 3.9
+ tnom = 25
+ rnoia = 0
+ rnoib = 0
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ cigbacc = 0.245
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ rdsmod = 0
+ igbmod = 1
+ pketa = 5.6398736e-15
+ ngate = 1.7e+20
+ wtvfbsdoff = 0
+ ijthsrev = 0.01
+ ngcon = 1
+ tnoimod = 0
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ wpclm = -1.1447315e-8
+ pbswgd = 0.8
+ pbswgs = 0.8
+ gbmin = 1e-12
+ cigbinv = 0.006
+ jswgd = 3.69e-13
+ ltvfbsdoff = 0
+ jswgs = 3.69e-13
+ igcmod = 1
+ wags = 3.4820603e-7
+ voff = -0.10461895
+ acde = 0.5
+ version = 4.5
+ ppdiblc2 = 9.4893758e-16
+ vsat = 91103.982
+ tempmod = 0
+ wint = 0
+ vth0 = -0.39207682
+ wkt1 = 1.4552168e-8
+ wkt2 = 6.9668931e-9
+ wmax = 5.4e-7
+ aigc = 0.0068462496
+ wmin = 2.7e-7
+ aigbacc = 0.012071
+ ptvfbsdoff = 0
+ tvoff = 0.0026312893
+ wua1 = 1.777316e-16
+ wub1 = 1.5048515e-26
+ wuc1 = -3.1929257e-17
+ permod = 1
+ xjbvd = 1
+ xjbvs = 1
+ bigc = 0.0012521
+ wute = 6.965504e-8
+ lk2we = 0.0
+ wwlc = 0
+ pkvth0we = 0.0
+ aigbinv = 0.009974
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ ku0we = -0.0007
+ beta0 = 13.32
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ voffcv = -0.125
+ wpemod = 1
+ cigc = 0.15259
+ vfbsdoff = 0.01
+ leta0 = 0
+ ppclm = 0
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ paramchk = 1
+ poxedge = 1
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ binunit = 2
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ tpbswg = 0.001
+ k2we = 5e-5
+ ijthdfwd = 0.01
+ dsub = 0.5
+ dtox = 3.91e-10
+ a0 = 2.4559917
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 72000
+ cf = 8.17e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.0065510297
+ k3 = -2.5823
+ em = 20000000.0
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ ll = 0
+ lw = 0
+ u0 = 0.011059968
+ w0 = 0
+ ua = 2.2475737e-10
+ ub = 1.3971204e-18
+ uc = 8.9671176e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 6e-9
+ bigsd = 0.0003327
+ ptvoff = 6.0034078e-17
+ eta0 = 0.17962267
+ etab = -0.19577778
+ waigsd = 1.9297907e-12
+ wvoff = -2.3606869e-9
+ ijthdrev = 0.01
+ wvsat = 0.0034765009
+ diomod = 1
+ wvth0 = -1.1167848e-9
+ lpdiblc2 = -1.0873556e-9
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ waigc = -6.0221967e-12
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.81e-10
+ pku0we = 0.0
+ cjswgs = 1.81e-10
+ lketa = -2.7133526e-8
+ xpart = 1
+ mjswgd = 0.95
+ mjswgs = 0.95
+ egidl = 0.001
+ tcjswg = 0.00128
+ pvfbsdoff = 0
+ lkvth0we = 3e-12
+ njtsswg = 6.489
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ acnqsmod = 0
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.012575691
+ pdiblcb = 0
+ rbodymod = 0
+ fprout = 200
+ xrcrg1 = 12
+ xrcrg2 = 1
+ pvoff = 1.5489261e-15
+ keta = 0.0057304489
+ cdscb = 0
+ cdscd = 0
+ pvsat = 0
+ bigbacc = 0.0054401
+ lags = 9.833094e-7
+ wk2we = 0.0
+ pvth0 = -1.2240418e-16
+ wtvoff = -1.9743529e-10
+ drout = 0.56
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 8.2671111e-11
+ paigc = 6.5097646e-18
+ kt1l = 0
+ kvth0we = -0.00022
+ voffl = 0
+ wpdiblc2 = -1.8846129e-9
+ lintnoi = -5e-9
+ capmod = 2
+ lint = 6.5375218e-9
+ bigbinv = 0.00149
+ weta0 = -1.7648176e-8
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ wetab = 1.9534667e-8
+ wku0we = 1.5e-11
+ lkt1 = -4.3329349e-9
+ lkt2 = -2.567581e-9
+ lpclm = 0
+ lmax = 8.9908e-7
+ lmin = 4.4908e-7
+ mobmod = 0
+ lpe0 = 6.44e-8
+ lpeb = 0
+ cgidl = 1
+ minv = -0.33
+ lua1 = 1.3348283e-16
+ lub1 = 2.1611253e-25
+ luc1 = 5.928335e-17
+ ndep = 1e+18
+ lute = 1.2896693e-7
+ wkvth0we = 0.0
+ lwlc = 0
+ moin = 5.5538
+ pbswd = 0.9
+ pbsws = 0.9
+ ags = -0.056621626
+ nigc = 2.291
+ trnqsmod = 0
+ cjd = 0.001346
+ cit = -8.7888889e-5
+ cjs = 0.001346
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 1.0572421799999999e-8
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ pdits = 0
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ cigsd = 0.013281
+ nfactor = 1
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ la0 = -1.8333262e-7
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0
+ pags = -2.41252e-13
+ kt1 = -0.20789546
+ kt2 = -0.0733757
+ lk2 = 2.3045842e-10
+ llc = 0
+ lln = 1
+ lu0 = -3.2234965e-10
+ mjd = 0.335
+ mjs = 0.335
+ lua = -5.402342e-17
+ lub = -8.029291e-26
+ luc = -6.9221885e-17
+ lud = 0
+ ntox = 1
+ lwc = 0
+ lwl = 0
+ pcit = 0
+ lwn = 1
+ pclm = 1.1689658
+ njd = 1.02
+ njs = 1.02
+ pa0 = -1.295362e-13
+ rgatemod = 0
+ nsd = 1e+20
+ pbd = 0.75
+ pk2we = 0.0
+ pat = 0
+ pbs = 0.75
+ pk2 = 6.34174e-16
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ tnjtsswg = 1
+ pu0 = -2.5304972e-16
+ prt = 0
+ pua = -1.1377853e-22
+ pub = 1.1787175e-31
+ puc = 2.8393052e-23
+ pud = 0
+ phin = 0.15
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 1.5353037e-9
+ ub1 = -2.5129786e-18
+ uc1 = 1.2019494e-10
+ tpb = 0.0016
+ tnoia = 0
+ wa0 = 1.4554629e-7
+ pkt1 = -1.0206874e-14
+ pkt2 = -7.3243565e-16
+ ute = -1.2205289
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 2.3228278e-9
+ nigbacc = 10
+ wlc = 0
+ wln = 1
+ wu0 = 3.4013886e-10
+ xgl = -8.2e-9
+ xgw = 0
+ peta0 = 0
+ wua = -1.1141771e-17
+ wub = -5.4878553e-26
+ wuc = -2.8229789e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ wketa = -8.9579586e-9
+ tpbsw = 0.0025
+ cjswd = 5.1e-11
+ cjsws = 5.1e-11
+ rbdb = 50
+ pua1 = -9.6760461e-23
+ prwb = 0
+ pub1 = 5.7312604e-33
+ prwg = 0
+ puc1 = -1.747778e-23
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ nigbinv = 2.171
+ pute = -4.8084303e-14
+ rdsw = 200
+ toxref = 3e-9
+ )

.model pch_tt_28 pmos (
+ level = 54
+ wtvfbsdoff = 0
+ lku0we = 1.8e-11
+ k2we = 5e-5
+ epsrox = 3.9
+ dsub = 0.5
+ dtox = 3.91e-10
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ ltvfbsdoff = 0
+ bigbacc = 0.0054401
+ rdsmod = 0
+ igbmod = 1
+ wkvth0we = 0.0
+ eta0 = 0.17962267
+ etab = -0.19577778
+ kvth0we = -0.00022
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ trnqsmod = 0
+ pbswgd = 0.8
+ lintnoi = -5e-9
+ pbswgs = 0.8
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ pvoff = -2.2654209e-16
+ igcmod = 1
+ cdscb = 0
+ cdscd = 0
+ pvsat = 0
+ wk2we = 0.0
+ pvth0 = -6.9676914e-16
+ ptvfbsdoff = 0
+ drout = 0.56
+ paigc = -3.9499473e-18
+ voffl = 0
+ rgatemod = 0
+ tnjtsswg = 1
+ weta0 = -1.7648176e-8
+ wetab = 1.9534667e-8
+ lpclm = 0
+ cgidl = 1
+ permod = 1
+ ags = -1.2539967
+ nfactor = 1
+ cjd = 0.001346
+ cit = -0.00036538451
+ cjs = 0.001346
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 1.38228675e-8
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ pbswd = 0.9
+ pbsws = 0.9
+ voffcv = -0.125
+ wpemod = 1
+ la0 = -4.7253353e-7
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0
+ kt1 = -0.16257215
+ kt2 = -0.066291072
+ lk2 = 9.2447077e-10
+ llc = -1.18e-13
+ lln = 0.7
+ lu0 = -5.4290454e-10
+ keta = -0.0061234738
+ mjd = 0.335
+ mjs = 0.335
+ lua = -1.0290148e-16
+ lub = -5.3060964e-27
+ luc = -4.0794824e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pdits = 0
+ pa0 = 9.7298482e-15
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ cigsd = 0.013281
+ pk2 = -2.0891363e-16
+ nigbacc = 10
+ lags = 1.5101544e-6
+ pu0 = 1.1540053e-17
+ dvt0w = 0
+ dvt1w = 0
+ prt = 0
+ dvt2w = 0
+ pua = -1.3867635e-23
+ pub = 2.1855871e-32
+ puc = -2.7646346e-24
+ pud = 0
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 2.0476918e-10
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 1.7313241e-9
+ ub1 = -1.3316629e-18
+ uc1 = 2.2670111e-10
+ kt1l = 0
+ tpb = 0.0016
+ wa0 = -1.7096745e-7
+ ute = -0.86054925
+ web = 6628.3
+ wec = -16935.0
+ pk2we = 0.0
+ wk2 = 4.238936e-9
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ wlc = 0
+ wln = 1
+ wu0 = -2.6120153e-10
+ xgl = -8.2e-9
+ xgw = 0
+ wua = -2.3821198e-16
+ wub = 1.6333936e-25
+ wuc = 4.2583136e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ nigbinv = 2.171
+ lint = 9.7879675e-9
+ tpbswg = 0.001
+ lkt1 = -2.4275192e-8
+ lkt2 = -5.6848171e-9
+ lmax = 4.4908e-7
+ tnoia = 0
+ lmin = 2.1577e-7
+ lpe0 = 6.44e-8
+ ijthsfwd = 0.01
+ lpeb = 0
+ peta0 = 0
+ wketa = -7.8373297e-10
+ minv = -0.33
+ tpbsw = 0.0025
+ lua1 = 4.723388e-17
+ lub1 = -3.0366637e-25
+ luc1 = 1.2420632e-17
+ ptvoff = 5.0195791e-17
+ cjswd = 5.1e-11
+ cjsws = 5.1e-11
+ ndep = 1e+18
+ fnoimod = 1
+ mjswd = 0.01
+ lute = -2.9424109e-8
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ waigsd = 1.9297907e-12
+ lwlc = 0
+ eigbinv = 1.1
+ moin = 5.5538
+ ijthsrev = 0.01
+ nigc = 2.291
+ diomod = 1
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.81e-10
+ pku0we = 0.0
+ cjswgs = 1.81e-10
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ tvfbsdoff = 0.1
+ pags = -3.3771496e-13
+ scref = 1e-6
+ a0 = 3.1132665
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 72000
+ cf = 8.17e-11
+ ntox = 1
+ mjswgd = 0.95
+ ef = 1.15
+ mjswgs = 0.95
+ k1 = 0.30425
+ k2 = -0.0081283305
+ k3 = -2.5823
+ pcit = -9.2716403e-18
+ em = 20000000.0
+ ppdiblc2 = -3.8737293e-16
+ pclm = 1.1689658
+ pigcd = 2.572
+ cigbacc = 0.245
+ ll = -1.18e-13
+ aigsd = 0.0063633912
+ lw = 0
+ u0 = 0.01156123
+ w0 = 0
+ ua = 3.3584387e-10
+ ub = 1.2266958e-18
+ uc = -5.8379738e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 6e-9
+ tcjswg = 0.00128
+ lvoff = -4.2658924e-9
+ phin = 0.15
+ tnoimod = 0
+ lvsat = 0
+ pkt1 = 6.8355166e-15
+ pkt2 = 2.2627554e-16
+ lvth0 = 4.5653579e-9
+ cigbinv = 0.006
+ delta = 0.018814
+ laigc = -1.8017042e-11
+ wvfbsdoff = 0
+ rnoia = 0
+ rnoib = 0
+ lvfbsdoff = 0
+ rbdb = 50
+ pua1 = -2.7108228e-23
+ pkvth0we = 0.0
+ prwb = 0
+ pub1 = 7.1177686e-32
+ prwg = 0
+ puc1 = 8.7727027e-25
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ pketa = 2.0432143e-15
+ version = 4.5
+ ngate = 1.7e+20
+ pute = 1.6065563e-14
+ fprout = 200
+ rdsw = 200
+ ngcon = 1
+ tempmod = 0
+ wpclm = -1.1447315e-8
+ xrcrg1 = 12
+ xrcrg2 = 1
+ vfbsdoff = 0.01
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ aigbacc = 0.012071
+ wtvoff = -1.7507555e-10
+ paramchk = 1
+ rshg = 14.1
+ capmod = 2
+ aigbinv = 0.009974
+ wku0we = 1.5e-11
+ mobmod = 0
+ ijthdfwd = 0.01
+ tvoff = 0.002323434
+ tnom = 25
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ poxedge = 1
+ ijthdrev = 0.01
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = 0
+ lpdiblc2 = 4.7505822e-10
+ binunit = 2
+ ppclm = 0
+ wags = 5.6744004e-7
+ wcit = 2.107191e-11
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ voff = -0.12137687
+ acde = 0.5
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ vsat = 91103.982
+ wint = 0
+ vth0 = -0.40006475
+ wkt1 = -2.4180539e-8
+ wkt2 = 4.7880041e-9
+ wmax = 5.4e-7
+ dmcgt = 0
+ aigc = 0.0067599617
+ wmin = 2.7e-7
+ tcjsw = 9.34e-5
+ lkvth0we = 3e-12
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ wua1 = 1.9431072e-17
+ wub1 = -1.3369336e-25
+ wuc1 = -7.3645279e-17
+ acnqsmod = 0
+ bigc = 0.0012521
+ bigsd = 0.0003327
+ wute = -7.6140111e-8
+ wwlc = 0
+ wvoff = 1.674468e-9
+ toxref = 3e-9
+ rbodymod = 0
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ wvsat = 0.0034765009
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ wvth0 = 1.885901e-10
+ cigc = 0.15259
+ waigc = 1.7749876e-11
+ njtsswg = 6.489
+ lketa = -2.19178e-8
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ ltvoff = -2.3990075e-10
+ xpart = 1
+ ckappad = 0.6
+ wpdiblc2 = 1.1524564e-9
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.0090247504
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ pdiblcb = 0
+ egidl = 0.001
+ pvfbsdoff = 0
+ )

.model pch_tt_29 pmos (
+ level = 54
+ ijthdrev = 0.01
+ ngcon = 1
+ pbswgd = 0.8
+ pbswgs = 0.8
+ wpclm = -1.2079184e-7
+ aigbinv = 0.009974
+ nigc = 2.291
+ igcmod = 1
+ lpdiblc2 = -1.1954251e-9
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ ntox = 1
+ pcit = -8.1298391e-18
+ pclm = 1.5407845
+ poxedge = 1
+ phin = 0.15
+ lkvth0we = 3e-12
+ pkt1 = -1.21482e-15
+ pkt2 = -1.4992738e-15
+ binunit = 2
+ permod = 1
+ tvoff = 0.00085372815
+ acnqsmod = 0
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ rbdb = 50
+ pua1 = 1.9617826e-23
+ prwb = 0
+ pub1 = -3.1346313e-32
+ prwg = 0
+ puc1 = 1.1713402e-23
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ rbodymod = 0
+ voffcv = -0.125
+ wpemod = 1
+ rdsw = 200
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = 0
+ ppclm = 2.3071337e-14
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ rshg = 14.1
+ wpdiblc2 = -7.3926191e-10
+ tpbswg = 0.001
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ njtsswg = 6.489
+ ptvoff = -3.132788e-17
+ tnom = 25
+ bigsd = 0.0003327
+ waigsd = 1.9297907e-12
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ wkvth0we = 0.0
+ wvoff = 3.1859801e-10
+ diomod = 1
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.016941733
+ trnqsmod = 0
+ pdiblcb = 0
+ wvsat = 0.0032472346
+ pditsd = 0
+ wvth0 = -4.9669425e-9
+ pditsl = 0
+ cjswgd = 1.81e-10
+ pku0we = 0.0
+ cjswgs = 1.81e-10
+ waigc = -1.7260908e-11
+ wags = -1.0331048e-6
+ wcit = 1.566053e-11
+ lketa = 7.1935383e-9
+ voff = -0.13201276
+ mjswgd = 0.95
+ mjswgs = 0.95
+ bigbacc = 0.0054401
+ acde = 0.5
+ xpart = 1
+ rgatemod = 0
+ tcjswg = 0.00128
+ vsat = 91523.884
+ wint = 0
+ tnjtsswg = 1
+ vth0 = -0.39762236
+ pvfbsdoff = 0
+ kvth0we = -0.00022
+ egidl = 0.001
+ wkt1 = 1.3972715e-8
+ wkt2 = 1.2965963e-8
+ wmax = 5.4e-7
+ aigc = 0.0067957378
+ wmin = 2.7e-7
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ wua1 = -2.0201942e-16
+ wub1 = 3.5220237e-25
+ wuc1 = -1.2500135e-16
+ bigc = 0.0012521
+ wwlc = 0
+ fprout = 200
+ cdsc = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ a0 = 1.1444157
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ at = 108550.2
+ xtid = 3
+ cf = 8.17e-11
+ xtis = 3
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.025395241
+ k3 = -2.5823
+ em = 20000000.0
+ ll = -1.18e-13
+ lw = 0
+ u0 = 0.0099217592
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ w0 = 0
+ ua = -3.1599722e-11
+ ub = 1.4008434e-18
+ uc = -1.6299488e-10
+ ud = 0
+ cigc = 0.15259
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 6e-9
+ pvoff = 5.9546471e-17
+ wtvoff = 2.1129256e-10
+ cdscb = 0
+ cdscd = 0
+ pvsat = 4.83709e-11
+ wk2we = 0.0
+ pvth0 = 3.9104824e-16
+ drout = 0.56
+ paigc = 3.4373281e-18
+ nfactor = 1
+ capmod = 2
+ voffl = 0
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ wku0we = 1.5e-11
+ dmdg = 0
+ weta0 = -1.7648176e-8
+ wetab = 1.9534667e-8
+ mobmod = 0
+ ags = 5.9031333
+ lpclm = -7.8453093e-8
+ cjd = 0.001346
+ cit = 0.00015305446
+ cjs = 0.001346
+ clc = 1e-7
+ cle = 0.6
+ k2we = 5e-5
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 1.38228675e-8
+ ijthsfwd = 0.01
+ k3b = 2.1176
+ dsub = 0.5
+ cgidl = 1
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ dtox = 3.91e-10
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ nigbacc = 10
+ la0 = -5.7105222e-8
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = -0.0077120921
+ kt1 = -0.27233533
+ kt2 = -0.10755274
+ lk2 = 4.5677889e-9
+ eta0 = 0.17962267
+ llc = -1.18e-13
+ lln = 0.7
+ lu0 = -1.969763e-10
+ etab = -0.19577778
+ mjd = 0.335
+ mjs = 0.335
+ lua = -2.5370884e-17
+ lub = -4.2051244e-26
+ luc = 1.7994313e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ pbswd = 0.9
+ pbsws = 0.9
+ njd = 1.02
+ njs = 1.02
+ pa0 = -3.159814e-15
+ ijthsrev = 0.01
+ nsd = 1e+20
+ pbd = 0.75
+ pat = -4.5415452e-10
+ pbs = 0.75
+ pk2 = -2.0710507e-16
+ pu0 = 4.0684676e-18
+ prt = 0
+ pua = 6.5898257e-24
+ pub = -4.9701536e-33
+ puc = -7.066739e-24
+ pud = 0
+ nigbinv = 2.171
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 2.8369875e-9
+ ub1 = -4.0389099e-18
+ uc1 = 4.2708978e-10
+ tpb = 0.0016
+ wa0 = -1.0988104e-7
+ pdits = 0
+ ute = -1
+ wat = 0.0021523911
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 4.2303646e-9
+ cigsd = 0.013281
+ wlc = 0
+ wln = 1
+ wu0 = -2.2579117e-10
+ xgl = -8.2e-9
+ xgw = 0
+ wua = -3.3516677e-16
+ dvt0w = 0
+ wub = 2.9047692e-25
+ wuc = 6.2972257e-17
+ wud = 0
+ dvt1w = 0
+ dvt2w = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ ppdiblc2 = 1.1779633e-17
+ pk2we = 0.0
+ fnoimod = 1
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ eigbinv = 1.1
+ tnoia = 0
+ peta0 = 0
+ wketa = 1.4826965e-8
+ tpbsw = 0.0025
+ cjswd = 5.1e-11
+ cjsws = 5.1e-11
+ pkvth0we = 0.0
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ toxref = 3e-9
+ cigbacc = 0.245
+ vfbsdoff = 0.01
+ tnoimod = 0
+ keta = -0.1440919
+ tvfbsdoff = 0.1
+ wtvfbsdoff = 0
+ cigbinv = 0.006
+ ltvoff = 7.0207177e-11
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 9.537856e-11
+ paramchk = 1
+ scref = 1e-6
+ kt1l = 0
+ pigcd = 2.572
+ aigsd = 0.0063633912
+ ltvfbsdoff = 0
+ version = 4.5
+ lvoff = -2.0217201e-9
+ lint = 9.7879675e-9
+ tempmod = 0
+ lkt1 = -1.1151622e-9
+ lkt2 = 3.021395e-9
+ lku0we = 1.8e-11
+ lmax = 2.1577e-7
+ lvsat = -8.85914e-5
+ lmin = 9e-8
+ epsrox = 3.9
+ lvth0 = 4.0500147e-9
+ lpe0 = 6.44e-8
+ ijthdfwd = 0.01
+ lpeb = 0
+ delta = 0.018814
+ laigc = -2.5565813e-11
+ aigbacc = 0.012071
+ wvfbsdoff = 0
+ rdsmod = 0
+ lvfbsdoff = 0
+ minv = -0.33
+ rnoia = 0
+ rnoib = 0
+ lua1 = -1.8606111e-16
+ lub1 = 2.6756274e-25
+ luc1 = -2.9861377e-17
+ igbmod = 1
+ ndep = 1e+18
+ ptvfbsdoff = 0
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ lwlc = 0
+ pketa = -1.250643e-15
+ ngate = 1.7e+20
+ moin = 5.5538
+ )

.model pch_tt_30 pmos (
+ level = 54
+ ijthdrev = 0.01
+ ngcon = 1
+ pbswgd = 0.8
+ pbswgs = 0.8
+ wpclm = 4.9341412e-7
+ aigbinv = 0.009974
+ nigc = 2.291
+ igcmod = 1
+ lpdiblc2 = 0
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ ntox = 1
+ pcit = -6.178865e-18
+ pclm = 0.08631615
+ paigsd = 8.4526218e-25
+ poxedge = 1
+ phin = 0.15
+ lkvth0we = 3e-12
+ pkt1 = -1.7124191e-15
+ pkt2 = 2.1480498e-17
+ binunit = 2
+ permod = 1
+ tvoff = 0.0012365685
+ acnqsmod = 0
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ rbdb = 50
+ pua1 = 4.1792962e-25
+ prwb = 0
+ pub1 = 6.1746384e-33
+ prwg = 0
+ puc1 = 2.9246063e-24
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ rbodymod = 0
+ voffcv = -0.125
+ wpemod = 1
+ rdsw = 200
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = -8.5658832e-9
+ letab = 1.7579973e-8
+ ppclm = -3.4664022e-14
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ rshg = 14.1
+ wpdiblc2 = -6.1394667e-10
+ tpbswg = 0.001
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ njtsswg = 6.489
+ ptvoff = 2.0376593e-17
+ tnom = 25
+ bigsd = 0.0003327
+ waigsd = 1.9297817e-12
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ wkvth0we = 0.0
+ wvoff = -2.8254962e-9
+ diomod = 1
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.0042244444
+ trnqsmod = 0
+ pdiblcb = 0
+ wvsat = 0.017016245
+ pditsd = 0
+ wvth0 = -3.8031861e-9
+ pditsl = 0
+ cjswgd = 1.81e-10
+ pku0we = 0.0
+ cjswgs = 1.81e-10
+ waigc = 7.1461687e-12
+ wags = -1.0331048e-6
+ wcit = -5.09452e-12
+ lketa = -1.1878561e-8
+ voff = -0.12098873
+ mjswgd = 0.95
+ mjswgs = 0.95
+ bigbacc = 0.0054401
+ acde = 0.5
+ xpart = 1
+ rgatemod = 0
+ tcjswg = 0.00128
+ vsat = 62231.739
+ wint = 0
+ tnjtsswg = 1
+ vth0 = -0.34146471
+ pvfbsdoff = 0
+ kvth0we = -0.00022
+ egidl = 0.001
+ wkt1 = 1.9266322e-8
+ wkt2 = -3.2122744e-9
+ wmax = 5.4e-7
+ aigc = 0.0067006504
+ wmin = 2.7e-7
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ wua1 = 2.2347963e-18
+ wub1 = -4.6956688e-26
+ wuc1 = -3.1503526e-17
+ bigc = 0.0012521
+ wwlc = 0
+ fprout = 200
+ cdsc = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ a0 = 3.9744452
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ at = 69068.642
+ xtid = 3
+ cf = 8.17e-11
+ xtis = 3
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.022825095
+ k3 = -2.5823
+ em = 20000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.0040856963
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ w0 = 0
+ ua = -9.2439852e-11
+ ub = -1.6232125e-18
+ uc = 5.3507127e-11
+ ud = 0
+ cigc = 0.15259
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 6e-9
+ pvoff = 3.5509132e-16
+ wtvoff = -3.3875503e-10
+ cdscb = 0
+ cdscd = 0
+ pvsat = -1.2459161e-9
+ wk2we = 0.0
+ pvth0 = 2.8165514e-16
+ drout = 0.56
+ paigc = 1.1430629e-18
+ nfactor = 1
+ capmod = 2
+ voffl = 0
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ wku0we = 1.5e-11
+ dmdg = 0
+ weta0 = -5.5015839e-8
+ wetab = 4.6876459e-8
+ mobmod = 0
+ ags = 5.9031333
+ lpclm = 5.8266931e-8
+ cjd = 0.001346
+ cit = -0.00018033605
+ cjs = 0.001346
+ clc = 1e-7
+ cle = 0.6
+ k2we = 5e-5
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 4.0349e-9
+ ijthsfwd = 0.01
+ k3b = 2.1176
+ dsub = 0.5
+ cgidl = 1
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ dtox = 3.91e-10
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ nigbacc = 10
+ la0 = -3.23128e-7
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = -0.0040008257
+ kt1 = -0.32608492
+ kt2 = -0.08284588
+ lk2 = 4.3261952e-9
+ eta0 = 0.27074908
+ llc = 0
+ lln = 1
+ lu0 = 3.5161362e-10
+ etab = -0.38279877
+ mjd = 0.335
+ mjs = 0.335
+ lua = -1.9651912e-17
+ lub = 2.4221001e-25
+ luc = -2.356876e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ pbswd = 0.9
+ pbsws = 0.9
+ njd = 1.02
+ njs = 1.02
+ pa0 = 9.1746422e-14
+ laigsd = -3.0625433e-18
+ ijthsrev = 0.01
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 6.7620954e-11
+ pbs = 0.75
+ pk2 = 2.5170462e-16
+ pu0 = -8.2666616e-17
+ prt = 0
+ pua = 3.032424e-23
+ pub = -9.6166295e-32
+ puc = -2.0363205e-24
+ pud = 0
+ nigbinv = 2.171
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = -2.7998083e-10
+ ub1 = 8.7083504e-19
+ uc1 = 1.8820988e-11
+ tpb = 0.0016
+ wa0 = -1.1195219e-6
+ pdits = 0
+ ute = -1
+ wat = -0.0033984119
+ web = 6628.3
+ wec = -16935.0
+ wk2 = -6.5058945e-10
+ cigsd = 0.013281
+ wlc = 0
+ wln = 1
+ wu0 = 6.9692249e-10
+ xgl = -8.2e-9
+ xgw = 0
+ wua = -5.8766054e-16
+ dvt0w = 0
+ wub = 1.2606486e-24
+ wuc = 9.4571662e-18
+ wud = 0
+ dvt1w = 0
+ dvt2w = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ ppdiblc2 = 0
+ pk2we = 0.0
+ fnoimod = 1
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ eigbinv = 1.1
+ tnoia = 0
+ peta0 = 3.5125603e-15
+ petab = -2.5701285e-15
+ wketa = -3.6489897e-8
+ tpbsw = 0.0025
+ cjswd = 5.1e-11
+ cjsws = 5.1e-11
+ pkvth0we = 0.0
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ toxref = 3e-9
+ cigbacc = 0.245
+ vfbsdoff = 0.01
+ tnoimod = 0
+ keta = 0.058802768
+ tvfbsdoff = 0.1
+ wtvfbsdoff = 0
+ cigbinv = 0.006
+ ltvoff = 3.4220189e-11
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 1.2671727e-10
+ paramchk = 1
+ scref = 1e-6
+ kt1l = 0
+ pigcd = 2.572
+ aigsd = 0.0063633912
+ ltvfbsdoff = 0
+ version = 4.5
+ lvoff = -3.0579783e-9
+ lint = 0
+ tempmod = 0
+ lkt1 = 3.9372999e-9
+ lkt2 = 6.989501e-10
+ lku0we = 1.8e-11
+ lmax = 9e-8
+ lvsat = 0.0026648703
+ lmin = 5.4e-8
+ epsrox = 3.9
+ lvth0 = -1.2288048e-9
+ lpe0 = 6.44e-8
+ ijthdfwd = 0.01
+ lpeb = 0
+ delta = 0.018814
+ laigc = -1.6627591e-11
+ aigbacc = 0.012071
+ wvfbsdoff = 0
+ rdsmod = 0
+ lvfbsdoff = 0
+ minv = -0.33
+ rnoia = 0
+ rnoib = 0
+ lua1 = 1.0693391e-16
+ lub1 = -1.9395329e-25
+ luc1 = 8.5158894e-18
+ igbmod = 1
+ ndep = 1e+18
+ ptvfbsdoff = 0
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ lwlc = 0
+ pketa = 3.573142e-15
+ ngate = 1.7e+20
+ moin = 5.5538
+ )

.model pch_tt_31 pmos (
+ level = 54
+ paigc = -3.8652128e-18
+ voff = -0.11425646
+ nigbacc = 10
+ ags = 5.9031333
+ acde = 0.5
+ ppdiblc2 = 0
+ voffl = 0
+ cjd = 0.001346
+ cit = -0.0023632098
+ cjs = 0.001346
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ vsat = 205509.49
+ dlc = 4.0349e-9
+ wint = 0
+ k3b = 2.1176
+ vth0 = -0.32141972
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ weta0 = 4.5569198e-8
+ wkt1 = -9.053012e-8
+ wkt2 = -4.5663135e-8
+ wetab = 2.1214781e-8
+ wmax = 5.4e-7
+ aigc = 0.0065523001
+ wmin = 2.7e-7
+ lpclm = -1.6067206e-7
+ permod = 1
+ nigbinv = 2.171
+ la0 = 2.2449695e-9
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = -0.00094527867
+ kt1 = -0.078489325
+ kt2 = 0.051187672
+ lk2 = 5.4231101e-9
+ llc = 0
+ lln = 1
+ cgidl = 1
+ lu0 = -6.4149203e-10
+ mjd = 0.335
+ mjs = 0.335
+ lua = -5.2618623e-17
+ lub = -3.080728e-25
+ luc = -2.0280652e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ wua1 = 2.8402308e-15
+ njs = 1.02
+ wub1 = -3.9062366e-24
+ wuc1 = 2.0276364e-16
+ pa0 = -4.432942e-14
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 1.8264736e-9
+ pbs = 0.75
+ pk2 = -1.1995676e-16
+ pu0 = 2.2577126e-16
+ bigc = 0.0012521
+ prt = 0
+ pua = 1.5923531e-23
+ pub = 9.2000466e-32
+ puc = 3.3504384e-24
+ pud = 0
+ wwlc = 0
+ pkvth0we = 0.0
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = -3.345352e-9
+ ub1 = 3.9080279e-18
+ uc1 = 1.4308247e-10
+ tpb = 0.0016
+ voffcv = -0.125
+ wpemod = 1
+ pbswd = 0.9
+ pbsws = 0.9
+ wa0 = 1.2266134e-6
+ cdsc = 0
+ ute = -1
+ wat = -0.033723458
+ web = 6628.3
+ wec = -16935.0
+ fnoimod = 1
+ wk2 = 5.7573654e-9
+ wlc = 0
+ cgbo = 0
+ wln = 1
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ wu0 = -4.6209719e-9
+ xtid = 3
+ xgl = -8.2e-9
+ xtis = 3
+ xgw = 0
+ wua = -3.3937245e-16
+ wub = -1.9836059e-24
+ wuc = -8.3417988e-17
+ wud = 0
+ eigbinv = 1.1
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ vfbsdoff = 0.01
+ cigc = 0.15259
+ pdits = 0
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ paramchk = 1
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ tpbswg = 0.001
+ cigbacc = 0.245
+ tnoia = 0
+ k2we = 5e-5
+ tnoimod = 0
+ ijthdfwd = 0.01
+ peta0 = -2.3213718e-15
+ dsub = 0.5
+ petab = -1.0817512e-15
+ dtox = 3.91e-10
+ wketa = 7.0696889e-8
+ ptvoff = -1.3332507e-17
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ tpbsw = 0.0025
+ waigsd = 1.9297962e-12
+ cigbinv = 0.006
+ cjswd = 5.1e-11
+ cjsws = 5.1e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ eta0 = 0.012687945
+ etab = -0.23454709
+ diomod = 1
+ ijthdrev = 0.01
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.81e-10
+ pku0we = 0.0
+ version = 4.5
+ cjswgs = 1.81e-10
+ lpdiblc2 = 0
+ tempmod = 0
+ tvfbsdoff = 0.1
+ aigbacc = 0.012071
+ mjswgd = 0.95
+ mjswgs = 0.95
+ scref = 1e-6
+ tcjswg = 0.00128
+ pigcd = 2.572
+ aigsd = 0.0063633912
+ lvoff = -3.4484499e-9
+ lkvth0we = 3e-12
+ aigbinv = 0.009974
+ lvsat = -0.0056452393
+ lvth0 = -2.3914143e-9
+ delta = 0.018814
+ wvfbsdoff = 0
+ laigc = -8.0232722e-12
+ lvfbsdoff = 0
+ rnoia = 0
+ rnoib = 0
+ acnqsmod = 0
+ fprout = 200
+ pketa = -2.6436916e-15
+ ngate = 1.7e+20
+ xrcrg1 = 12
+ xrcrg2 = 1
+ rbodymod = 0
+ ngcon = 1
+ wpclm = -6.9641486e-7
+ poxedge = 1
+ gbmin = 1e-12
+ wtvoff = 2.4243635e-10
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ keta = -0.44725926
+ binunit = 2
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 2.5332395e-10
+ capmod = 2
+ kt1l = 0
+ wku0we = 1.5e-11
+ wpdiblc2 = -6.1394667e-10
+ mobmod = 0
+ lint = 0
+ lkt1 = -1.0423245e-8
+ lkt2 = -7.0749959e-9
+ lmax = 5.4e-8
+ lmin = 4.5e-8
+ a0 = -1.6354335
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 16386.797
+ cf = 8.17e-11
+ lpe0 = 6.44e-8
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.041737421
+ k3 = -2.5823
+ em = 20000000.0
+ lpeb = 0
+ ll = 0
+ lw = 0
+ u0 = 0.021208207
+ w0 = 0
+ tvoff = 0.0019328761
+ ua = 4.7595173e-10
+ ub = 7.8644222e-18
+ uc = 4.7837975e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 6e-9
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ minv = -0.33
+ xjbvd = 1
+ xjbvs = 1
+ lua1 = 2.8472544e-16
+ lub1 = -3.7011047e-25
+ lk2we = 0.0
+ luc1 = 1.3087235e-18
+ ndep = 1e+18
+ wkvth0we = 0.0
+ lwlc = 0
+ moin = 5.5538
+ ku0we = -0.0007
+ trnqsmod = 0
+ nigc = 2.291
+ beta0 = 13.32
+ leta0 = 6.4016629e-9
+ letab = 8.9813755e-9
+ ppclm = 3.4346058e-14
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ njtsswg = 6.489
+ ntox = 1
+ pcit = -1.762461e-17
+ pclm = 3.8611263
+ rgatemod = 0
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ tnjtsswg = 1
+ dmcgt = 0
+ ckappad = 0.6
+ phin = 0.15
+ ckappas = 0.6
+ tcjsw = 9.34e-5
+ pdiblc1 = 0
+ pdiblc2 = 0.0042244444
+ pdiblcb = 0
+ pkt1 = 4.6557745e-15
+ pkt2 = 2.4836304e-15
+ bigsd = 0.0003327
+ toxref = 3e-9
+ rbdb = 50
+ pua1 = -1.6418584e-22
+ prwb = 0
+ pub1 = 2.3001287e-31
+ prwg = 0
+ puc1 = -1.0662889e-23
+ wtvfbsdoff = 0
+ bigbacc = 0.0054401
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ wvoff = 3.9335999e-9
+ rdsw = 200
+ wvsat = -0.031328619
+ kvth0we = -0.00022
+ ltvfbsdoff = 0
+ wvth0 = 1.1142981e-8
+ waigc = 9.3495749e-11
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ ltvoff = -6.1656569e-12
+ lketa = 1.7473037e-8
+ xpart = 1
+ rshg = 14.1
+ pvfbsdoff = 0
+ egidl = 0.001
+ ptvfbsdoff = 0
+ lku0we = 1.8e-11
+ epsrox = 3.9
+ ijthsfwd = 0.01
+ rdsmod = 0
+ igbmod = 1
+ tnom = 25
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ nfactor = 1
+ pbswgd = 0.8
+ pbswgs = 0.8
+ ijthsrev = 0.01
+ igcmod = 1
+ pvoff = -3.6936248e-17
+ cdscb = 0
+ cdscd = 0
+ wags = -1.0331048e-6
+ pvsat = 1.5580861e-9
+ wk2we = 0.0
+ pvth0 = -5.8522254e-16
+ wcit = 1.9224593e-10
+ drout = 0.56
+ )

.model pch_tt_32 pmos (
+ level = 54
+ tvoff = 0.0050068134
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ voffcv = -0.125
+ wpemod = 1
+ njtsswg = 6.489
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = 2.7114638e-9
+ ckappad = 0.6
+ letab = 1.8240871e-9
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.0042244444
+ pdiblcb = 0
+ keta = -0.10111506
+ ppclm = 1.7398739e-15
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = -4.8395e-12
+ kt1l = 0
+ tpbswg = 0.001
+ bigbacc = 0.0054401
+ lint = 0
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ lkt1 = -1.3409032e-8
+ lkt2 = 2.2261728e-10
+ lmax = 4.5e-8
+ kvth0we = -0.00022
+ lmin = 3.6e-8
+ lpe0 = 6.44e-8
+ ijthsfwd = 0.01
+ lpeb = 0
+ ptvoff = 3.2244316e-17
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ waigsd = 1.9257033e-12
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ minv = -0.33
+ bigsd = 0.0003327
+ lua1 = -1.7116539e-16
+ lub1 = 1.8549471e-25
+ luc1 = 2.2025561e-17
+ ndep = 1e+18
+ diomod = 1
+ lwlc = 0
+ wvoff = 1.094003e-8
+ moin = 5.5538
+ ijthsrev = 0.01
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.81e-10
+ pku0we = 0.0
+ cjswgs = 1.81e-10
+ nigc = 2.291
+ wvsat = -0.018712604
+ wvth0 = 1.5582333e-8
+ waigc = 1.753535e-10
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ mjswgd = 0.95
+ mjswgs = 0.95
+ lketa = 5.1197136e-10
+ tcjswg = 0.00128
+ xpart = 1
+ ntox = 1
+ ppdiblc2 = 0
+ pcit = 1.2154904e-16
+ pclm = 0.85281474
+ pvfbsdoff = 0
+ nfactor = 1
+ egidl = 0.001
+ phin = 0.15
+ pkt1 = 2.438466e-15
+ pkt2 = -1.2154904e-16
+ fprout = 200
+ pkvth0we = 0.0
+ rbdb = 50
+ pua1 = 5.9435365e-23
+ prwb = 0
+ pub1 = -6.8901825e-32
+ prwg = 0
+ puc1 = -3.4884574e-24
+ xrcrg1 = 12
+ xrcrg2 = 1
+ nigbacc = 10
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ rdsw = 200
+ wtvoff = -6.8770288e-10
+ vfbsdoff = 0.01
+ pvoff = -3.8025133e-16
+ ags = 5.9031333
+ nigbinv = 2.171
+ cdscb = 0
+ cdscd = 0
+ cjd = 0.001346
+ cit = 0.0029054321
+ cjs = 0.001346
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ pvsat = 9.3990127e-10
+ dlc = 4.0349e-9
+ wk2we = 0.0
+ pvth0 = -8.027508e-16
+ k3b = 2.1176
+ dwb = 0
+ drout = 0.56
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ capmod = 2
+ paramchk = 1
+ paigc = -7.8762427e-18
+ wku0we = 1.5e-11
+ rshg = 14.1
+ voffl = 0
+ la0 = -2.1218621e-7
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0.010508083
+ mobmod = 0
+ kt1 = -0.017554887
+ kt2 = -0.09774321
+ lk2 = 4.0572258e-9
+ llc = 0
+ lln = 1
+ lu0 = -2.435917e-10
+ mjd = 0.335
+ mjs = 0.335
+ lua = 4.1444844e-17
+ lub = -1.5666965e-25
+ luc = -1.4956542e-17
+ lud = 0
+ lwc = 0
+ weta0 = 6.7301382e-9
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ wetab = -5.613608e-9
+ njs = 1.02
+ pa0 = 5.0455005e-14
+ fnoimod = 1
+ nsd = 1e+20
+ pbd = 0.75
+ pat = -2.4847929e-9
+ pbs = 0.75
+ pk2 = 3.3742201e-16
+ lpclm = -1.3264792e-8
+ pu0 = 1.5059926e-16
+ eigbinv = 1.1
+ prt = 0
+ pua = 9.2877876e-24
+ pub = 3.2782262e-32
+ puc = 3.1614905e-24
+ pud = 0
+ ijthdfwd = 0.01
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 5.9585425e-9
+ ub1 = -7.4308533e-18
+ uc1 = -2.7971012e-10
+ cgidl = 1
+ tpb = 0.0016
+ wa0 = -7.0776268e-7
+ ute = -1
+ wat = 0.054261574
+ web = 6628.3
+ wec = -16935.0
+ wk2 = -3.5768953e-9
+ wlc = 0
+ wln = 1
+ wu0 = -3.0868494e-9
+ tnom = 25
+ xgl = -8.2e-9
+ xgw = 0
+ wua = -2.0394912e-16
+ wub = -7.7507108e-25
+ wuc = -7.9561907e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ laigsd = -3.6731852e-16
+ pbswd = 0.9
+ pbsws = 0.9
+ ijthdrev = 0.01
+ cigbacc = 0.245
+ lpdiblc2 = 0
+ pdits = 0
+ wags = -1.0331048e-6
+ cigsd = 0.013281
+ tnoimod = 0
+ dvt0w = 0
+ dvt1w = 0
+ wcit = -2.6480326e-9
+ dvt2w = 0
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ a0 = 2.7407131
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = -217355.29
+ cf = 8.17e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.013862232
+ k3 = -2.5823
+ em = 20000000.0
+ voff = -0.14966725
+ ll = 0
+ lw = 0
+ u0 = 0.013087793
+ w0 = 0
+ cigbinv = 0.006
+ acde = 0.5
+ ua = -1.4437109e-9
+ ub = 4.7745619e-18
+ uc = 3.1168444e-10
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 6e-9
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ vsat = 182315.32
+ wint = 0
+ vth0 = -0.39307143
+ wkt1 = -4.5278925e-8
+ wkt2 = 7.5037926e-9
+ wtvfbsdoff = 0
+ wmax = 5.4e-7
+ aigc = 0.006152944
+ wmin = 2.7e-7
+ lkvth0we = 3e-12
+ tnoia = 0
+ version = 4.5
+ tempmod = 0
+ peta0 = -4.1825789e-16
+ ltvfbsdoff = 0
+ petab = 2.3283989e-16
+ wketa = 1.3494424e-8
+ wua1 = -1.7234672e-15
+ wub1 = 2.1940634e-24
+ wuc1 = 5.6346661e-17
+ tpbsw = 0.0025
+ acnqsmod = 0
+ toxref = 3e-9
+ bigc = 0.0012521
+ aigbacc = 0.012071
+ cjswd = 5.1e-11
+ cjsws = 5.1e-11
+ wwlc = 0
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ rbodymod = 0
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigc = 0.15259
+ aigbinv = 0.009974
+ tvfbsdoff = 0.1
+ ptvfbsdoff = 0
+ ltvoff = -1.5678858e-10
+ scref = 1e-6
+ pigcd = 2.572
+ aigsd = 0.0063633987
+ wpdiblc2 = -6.1394667e-10
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ lku0we = 1.8e-11
+ lvoff = -1.7133213e-9
+ epsrox = 3.9
+ lvsat = -0.0045087251
+ poxedge = 1
+ lvth0 = 1.1195196e-9
+ k2we = 5e-5
+ wvfbsdoff = 0
+ rdsmod = 0
+ lvfbsdoff = 0
+ delta = 0.018814
+ dsub = 0.5
+ dtox = 3.91e-10
+ laigc = 1.1545174e-11
+ igbmod = 1
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ binunit = 2
+ rnoia = 0
+ rnoib = 0
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ pbswgd = 0.8
+ wkvth0we = 0.0
+ pbswgs = 0.8
+ eta0 = 0.08799813
+ pketa = 1.5922924e-16
+ etab = -0.088479977
+ ngate = 1.7e+20
+ ngcon = 1
+ igcmod = 1
+ wpclm = -3.0982532e-8
+ trnqsmod = 0
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ paigsd = 2.0055591e-22
+ rgatemod = 0
+ tnjtsswg = 1
+ permod = 1
+ )

.model pch_tt_33 pmos (
+ level = 54
+ version = 4.5
+ pdits = 0
+ cigsd = 0.013281
+ tempmod = 0
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ tpbswg = 0.001
+ rshg = 14.1
+ aigbacc = 0.012071
+ wpdiblc2 = 3.3638075e-10
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ tnoia = 0
+ ptvoff = 0
+ aigbinv = 0.009974
+ peta0 = 0
+ waigsd = 1.9846811e-12
+ wketa = -1.9384664e-9
+ tpbsw = 0.0025
+ tnom = 25
+ diomod = 1
+ cjswd = 5.1e-11
+ cjsws = 5.1e-11
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ wkvth0we = 0.0
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.81e-10
+ pku0we = 0.0
+ cjswgs = 1.81e-10
+ trnqsmod = 0
+ tvfbsdoff = 0.1
+ poxedge = 1
+ mjswgd = 0.95
+ wags = 5.1942014e-9
+ mjswgs = 0.95
+ tcjswg = 0.00128
+ binunit = 2
+ scref = 1e-6
+ voff = -0.10372023
+ acde = 0.5
+ pigcd = 2.572
+ aigsd = 0.0063632583
+ rgatemod = 0
+ vsat = 108525.44
+ tnjtsswg = 1
+ wint = 0
+ vth0 = -0.37287116
+ lvoff = 0
+ wkt1 = -3.0503659e-9
+ wkt2 = -7.2833333e-10
+ wmax = 2.7e-7
+ aigc = 0.0068302204
+ wmin = 1.08e-7
+ lvsat = 0
+ lvth0 = 0
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ delta = 0.018814
+ wua1 = -5.5326541e-17
+ wub1 = -1.0689498e-25
+ wuc1 = -1.2119467e-17
+ fprout = 200
+ rnoia = 0
+ rnoib = 0
+ bigc = 0.0012521
+ wute = -7.6523556e-8
+ xrcrg1 = 12
+ xrcrg2 = 1
+ wwlc = 0
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ ngate = 1.7e+20
+ ngcon = 1
+ cdsc = 0
+ wpclm = 7.1298978e-9
+ cgbo = 0
+ cgdl = 3.0105e-11
+ wtvoff = -7.3630015e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigc = 0.15259
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ capmod = 2
+ wku0we = 1.5e-11
+ mobmod = 0
+ njtsswg = 6.489
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ k2we = 5e-5
+ ckappad = 0.6
+ ckappas = 0.6
+ ijthsfwd = 0.01
+ pdiblc1 = 0
+ pdiblc2 = 0.0015492917
+ dsub = 0.5
+ pdiblcb = 0
+ dtox = 3.91e-10
+ tvoff = 0.0025423547
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ eta0 = 0.10792519
+ etab = -0.13555556
+ ijthsrev = 0.01
+ ku0we = -0.0007
+ bigbacc = 0.0054401
+ beta0 = 13.32
+ leta0 = 0
+ wtvfbsdoff = 0
+ kvth0we = -0.00022
+ ppclm = 0
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ dlcig = 2.5e-9
+ lintnoi = -5e-9
+ bgidl = 1834800000.0
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ ltvfbsdoff = 0
+ ppdiblc2 = 0
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ toxref = 3e-9
+ bigsd = 0.0003327
+ ptvfbsdoff = 0
+ pkvth0we = 0.0
+ wvoff = 1.4142431e-9
+ a0 = 2.5876667
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 72000
+ cf = 8.17e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.015389268
+ k3 = -2.5823
+ em = 20000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.0095671852
+ w0 = 0
+ ua = -1.9215717e-10
+ ub = 1.2747184e-18
+ uc = -1.7585185e-12
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 6e-9
+ wvsat = -0.0013318206
+ nfactor = 1
+ wvth0 = -3.2254372e-9
+ vfbsdoff = 0.01
+ waigc = 1.6569661e-12
+ keta = 0.02482765
+ ltvoff = 0
+ jswd = 3.69e-13
+ lketa = 0
+ jsws = 3.69e-13
+ paramchk = 1
+ lcit = 0
+ xpart = 1
+ pvfbsdoff = 0
+ kt1l = 0
+ lku0we = 1.8e-11
+ nigbacc = 10
+ egidl = 0.001
+ epsrox = 3.9
+ lint = 6.5375218e-9
+ lkt1 = 0
+ lmax = 2.001e-5
+ lmin = 8.9991e-6
+ rdsmod = 0
+ ijthdfwd = 0.01
+ lpe0 = 6.44e-8
+ igbmod = 1
+ lpeb = 0
+ nigbinv = 2.171
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ minv = -0.33
+ pbswgd = 0.8
+ pbswgs = 0.8
+ ndep = 1e+18
+ ags = 0.89683683
+ lwlc = 0
+ igcmod = 1
+ moin = 5.5538
+ ijthdrev = 0.01
+ cjd = 0.001346
+ cit = 5e-6
+ cjs = 0.001346
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 1.0572421799999999e-8
+ nigc = 2.291
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ lpdiblc2 = 0
+ fnoimod = 1
+ pvoff = 0
+ eigbinv = 1.1
+ cdscb = 0
+ cdscd = 0
+ la0 = 0
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ jsd = 1.5e-7
+ pvsat = 0
+ jss = 1.5e-7
+ lat = 0
+ kt1 = -0.17197747
+ lk2 = 0
+ kt2 = -0.050761111
+ wk2we = 0.0
+ pvth0 = 0
+ llc = 0
+ lln = 1
+ lu0 = 0
+ drout = 0.56
+ mjd = 0.335
+ mjs = 0.335
+ lub = 0
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 0
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ pk2 = 0
+ pu0 = 0
+ ntox = 1
+ voffl = 0
+ prt = 0
+ pub = 0
+ pcit = 0
+ pud = 0
+ pclm = 1.101657
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 9.8162749e-10
+ ub1 = -3.8648101e-20
+ uc1 = 8.1681111e-11
+ tpb = 0.0016
+ weta0 = 2.1403289e-9
+ permod = 1
+ wa0 = 4.8944e-8
+ wetab = 2.9133333e-9
+ ute = -0.81574074
+ phin = 0.15
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 3.9065138e-9
+ lkvth0we = 3e-12
+ lpclm = 0
+ wlc = 0
+ wln = 1
+ wu0 = 5.8460889e-11
+ xgl = -8.2e-9
+ xgw = 0
+ wua = -4.8614483e-17
+ wub = 8.106039e-27
+ wuc = 3.3309111e-18
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ cigbacc = 0.245
+ pkt1 = 0
+ cgidl = 1
+ tnoimod = 0
+ acnqsmod = 0
+ voffcv = -0.125
+ wpemod = 1
+ rbdb = 50
+ prwb = 0
+ prwg = 0
+ rbpb = 50
+ rbpd = 50
+ cigbinv = 0.006
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ pbswd = 0.9
+ rbodymod = 0
+ pbsws = 0.9
+ rdsw = 200
+ )

.model pch_tt_34 pmos (
+ level = 54
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ nfactor = 1
+ ptvoff = -5.393716e-17
+ k2we = 5e-5
+ waigsd = 1.9861139e-12
+ ijthdfwd = 0.01
+ dsub = 0.5
+ dtox = 3.91e-10
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ diomod = 1
+ bigsd = 0.0003327
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.81e-10
+ pku0we = 0.0
+ cjswgs = 1.81e-10
+ eta0 = 0.10792519
+ wvoff = 1.3100722e-9
+ etab = -0.13555556
+ ijthdrev = 0.01
+ nigbacc = 10
+ wvsat = -0.0013318206
+ wvth0 = -3.3211131e-9
+ lpdiblc2 = 6.2970633e-9
+ waigc = 1.4905459e-12
+ mjswgd = 0.95
+ mjswgs = 0.95
+ tcjswg = 0.00128
+ nigbinv = 2.171
+ lketa = -5.5366519e-8
+ pvfbsdoff = 0
+ xpart = 1
+ egidl = 0.001
+ lkvth0we = 3e-12
+ fnoimod = 1
+ ags = 0.84380759
+ eigbinv = 1.1
+ fprout = 200
+ cjd = 0.001346
+ cit = 5e-6
+ cjs = 0.001346
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ acnqsmod = 0
+ dlc = 1.0572421799999999e-8
+ xrcrg1 = 12
+ xrcrg2 = 1
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ rbodymod = 0
+ la0 = -3.9401851e-7
+ wtvoff = -6.7630331e-11
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0
+ kt1 = -0.17107141
+ kt2 = -0.050597496
+ lk2 = 5.5319403e-9
+ llc = 0
+ lln = 1
+ lu0 = 9.9678999e-10
+ mjd = 0.335
+ mjs = 0.335
+ lua = -7.2048384e-17
+ lub = 4.3514377e-25
+ luc = 1.4270275e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = -3.1655381e-14
+ pvoff = 9.3649624e-16
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ pk2 = 9.285497e-17
+ keta = 0.030986328
+ pu0 = 3.0504276e-17
+ prt = 0
+ cdscb = 0
+ cdscd = 0
+ pua = 2.7735079e-23
+ pub = -4.2717478e-32
+ puc = 1.20866e-25
+ pud = 0
+ cigbacc = 0.245
+ capmod = 2
+ pvsat = 0
+ rsh = 15.2
+ wk2we = 0.0
+ tcj = 0.000832
+ ua1 = 8.0734953e-10
+ pvth0 = 8.6012639e-16
+ ub1 = 2.6826436e-19
+ uc1 = 8.9789043e-11
+ drout = 0.56
+ lags = 4.7673289e-7
+ wku0we = 1.5e-11
+ tpb = 0.0016
+ wa0 = 5.2465177e-8
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ ute = -0.817454
+ paigc = 1.4961177e-18
+ lcit = 0
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 3.8961851e-9
+ tnoimod = 0
+ mobmod = 0
+ wlc = 0
+ wln = 1
+ wu0 = 5.5067755e-11
+ xgl = -8.2e-9
+ xgw = 0
+ kt1l = 0
+ wua = -5.1699586e-17
+ wub = 1.2857705e-26
+ wuc = 3.3174666e-18
+ wud = 0
+ voffl = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ wpdiblc2 = 3.5925269e-10
+ cigbinv = 0.006
+ weta0 = 2.1403289e-9
+ wetab = 2.9133333e-9
+ lint = 6.5375218e-9
+ lpclm = 0
+ lkt1 = -8.1454893e-9
+ lkt2 = -1.4709041e-9
+ lmax = 8.9991e-6
+ lmin = 8.9908e-7
+ lpe0 = 6.44e-8
+ cgidl = 1
+ lpeb = 0
+ version = 4.5
+ tempmod = 0
+ minv = -0.33
+ wtvfbsdoff = 0
+ laigsd = -1.8524358e-14
+ lua1 = 1.5667589e-15
+ lub1 = -2.759143e-24
+ luc1 = -7.2890309e-17
+ ndep = 1e+18
+ wkvth0we = 0.0
+ lute = 1.5402209e-8
+ lwlc = 0
+ pbswd = 0.9
+ pbsws = 0.9
+ moin = 5.5538
+ aigbacc = 0.012071
+ ltvfbsdoff = 0
+ trnqsmod = 0
+ nigc = 2.291
+ pdits = 0
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ noff = 2.2684
+ cigsd = 0.013281
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ aigbinv = 0.009974
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ pags = -1.92428e-14
+ ntox = 1
+ pcit = 0
+ rgatemod = 0
+ pclm = 1.101657
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ ptvfbsdoff = 0
+ tnjtsswg = 1
+ phin = 0.15
+ tnoia = 0
+ pkt1 = -2.8122214e-15
+ pkt2 = 2.4239149e-16
+ peta0 = 0
+ toxref = 3e-9
+ wketa = -2.0595747e-9
+ poxedge = 1
+ tpbsw = 0.0025
+ cjswd = 5.1e-11
+ cjsws = 5.1e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ rbdb = 50
+ pua1 = -1.1776704e-22
+ binunit = 2
+ prwb = 0
+ pub1 = 2.7996299e-31
+ prwg = 0
+ puc1 = 9.811687e-24
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ pute = 1.5923616e-14
+ rdsw = 200
+ tvfbsdoff = 0.1
+ ltvoff = -3.3500511e-10
+ scref = 1e-6
+ pigcd = 2.572
+ rshg = 14.1
+ aigsd = 0.0063632604
+ lku0we = 1.8e-11
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ epsrox = 3.9
+ lvoff = -2.4480721e-8
+ a0 = 2.6314952
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ rdsmod = 0
+ wvfbsdoff = 0
+ at = 72000
+ cf = 8.17e-11
+ lvsat = 0
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.016004612
+ k3 = -2.5823
+ em = 20000000.0
+ lvfbsdoff = 0
+ lvth0 = -1.3866904e-8
+ igbmod = 1
+ ll = 0
+ lw = 0
+ u0 = 0.0094563075
+ w0 = 0
+ ua = -1.8414289e-10
+ ub = 1.2263153e-18
+ uc = -3.3458683e-12
+ ud = 0
+ ijthsfwd = 0.01
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 6e-9
+ delta = 0.018814
+ laigc = -5.3027874e-11
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ rnoia = 0
+ rnoib = 0
+ pbswgd = 0.8
+ pbswgs = 0.8
+ tnom = 25
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ igcmod = 1
+ pketa = 1.0887638e-15
+ ngate = 1.7e+20
+ ngcon = 1
+ ijthsrev = 0.01
+ wpclm = 7.1298978e-9
+ njtsswg = 6.489
+ gbmin = 1e-12
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ wags = 7.3346686e-9
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.00084883969
+ pdiblcb = 0
+ paigsd = -1.2880862e-20
+ voff = -0.10099712
+ acde = 0.5
+ ppdiblc2 = -2.0561872e-16
+ vsat = 108525.44
+ wint = 0
+ permod = 1
+ vth0 = -0.37132868
+ wkt1 = -2.7375492e-9
+ wkt2 = -7.5529568e-10
+ wmax = 2.7e-7
+ aigc = 0.0068361189
+ wmin = 1.08e-7
+ bigbacc = 0.0054401
+ tvoff = 0.0025796189
+ kvth0we = -0.00022
+ wua1 = -4.222676e-17
+ wub1 = -1.3803658e-25
+ wuc1 = -1.3210867e-17
+ xjbvd = 1
+ xjbvs = 1
+ voffcv = -0.125
+ wpemod = 1
+ lk2we = 0.0
+ lintnoi = -5e-9
+ bigc = 0.0012521
+ wute = -7.8294814e-8
+ bigbinv = 0.00149
+ pkvth0we = 0.0
+ wwlc = 0
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ cdsc = 0
+ ku0we = -0.0007
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ beta0 = 13.32
+ leta0 = 0
+ vfbsdoff = 0.01
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigc = 0.15259
+ ppclm = 0
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ paramchk = 1
+ tpbswg = 0.001
+ )

.model pch_tt_35 pmos (
+ level = 54
+ cjsws = 5.1e-11
+ cjswgd = 1.81e-10
+ pku0we = 0.0
+ cjswgs = 1.81e-10
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ ndep = 1e+18
+ lute = -1.0958354e-8
+ lwlc = 0
+ moin = 5.5538
+ ijthsrev = 0.01
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ tvfbsdoff = 0.1
+ nigc = 2.291
+ mjswgd = 0.95
+ mjswgs = 0.95
+ tcjswg = 0.00128
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ scref = 1e-6
+ pags = 1.1742809e-13
+ ppdiblc2 = -6.1367245e-16
+ pigcd = 2.572
+ ntox = 1
+ aigsd = 0.0063632396
+ pcit = 0
+ pclm = 1.101657
+ lvoff = -2.4340257e-9
+ phin = 0.15
+ wvfbsdoff = 0
+ njtsswg = 6.489
+ lvfbsdoff = 0
+ lvsat = 0
+ lvth0 = -2.799405e-11
+ pkt1 = 5.7473332e-15
+ pkt2 = -5.7270183e-16
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ delta = 0.018814
+ fprout = 200
+ laigc = -3.3884553e-11
+ xrcrg1 = 12
+ xrcrg2 = 1
+ ckappad = 0.6
+ ckappas = 0.6
+ rnoia = 0
+ rnoib = 0
+ pdiblc1 = 0
+ pdiblc2 = 0.0027845581
+ pdiblcb = 0
+ pkvth0we = 0.0
+ rbdb = 50
+ pua1 = -9.8048843e-24
+ prwb = 0
+ pub1 = -2.3189739e-32
+ prwg = 0
+ puc1 = -4.5795492e-24
+ pketa = -3.0075994e-15
+ rbpb = 50
+ rbpd = 50
+ ngate = 1.7e+20
+ rbps = 50
+ rbsb = 50
+ wtvoff = -2.2790108e-10
+ pvag = 2.1
+ pute = -9.4649237e-15
+ ngcon = 1
+ wpclm = 7.1298978e-9
+ rdsw = 200
+ vfbsdoff = 0.01
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ bigbacc = 0.0054401
+ capmod = 2
+ wku0we = 1.5e-11
+ kvth0we = -0.00022
+ mobmod = 0
+ paramchk = 1
+ lintnoi = -5e-9
+ rshg = 14.1
+ bigbinv = 0.00149
+ wtvfbsdoff = 0
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ ltvfbsdoff = 0
+ ijthdfwd = 0.01
+ tvoff = 0.0027416725
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ tnom = 25
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ ijthdrev = 0.01
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = 0
+ lpdiblc2 = 4.574275e-9
+ ptvfbsdoff = 0
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ nfactor = 1
+ ppclm = 0
+ wags = -1.4622812e-7
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ voff = -0.12576869
+ acde = 0.5
+ vsat = 108525.44
+ wint = 0
+ vth0 = -0.38687802
+ wkt1 = -1.2355026e-8
+ wkt2 = 1.605395e-10
+ dmcgt = 0
+ wmax = 2.7e-7
+ tcjsw = 9.34e-5
+ lkvth0we = 3e-12
+ aigc = 0.0068146096
+ wmin = 1.08e-7
+ nigbacc = 10
+ toxref = 3e-9
+ wua1 = -1.6353255e-16
+ wub1 = 2.0258446e-25
+ wuc1 = 2.9590615e-18
+ acnqsmod = 0
+ bigsd = 0.0003327
+ bigc = 0.0012521
+ wute = -4.9768365e-8
+ nigbinv = 2.171
+ wwlc = 0
+ wvoff = 3.4766421e-9
+ rbodymod = 0
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ wvsat = -0.0013318206
+ xtid = 3
+ xtis = 3
+ wvth0 = -2.5516532e-9
+ ltvoff = -4.7923289e-10
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigc = 0.15259
+ waigc = 2.7104678e-12
+ fnoimod = 1
+ eigbinv = 1.1
+ pvfbsdoff = 0
+ lketa = 4.197898e-9
+ xpart = 1
+ lku0we = 1.8e-11
+ epsrox = 3.9
+ wpdiblc2 = 8.1773971e-10
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ ags = 1.7348065
+ dmdg = 0
+ egidl = 0.001
+ cjd = 0.001346
+ rdsmod = 0
+ cit = -8.7888889e-5
+ cjs = 0.001346
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 1.0572421799999999e-8
+ igbmod = 1
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ k2we = 5e-5
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ dsub = 0.5
+ dtox = 3.91e-10
+ pbswgd = 0.8
+ la0 = -1.044589e-6
+ cigbacc = 0.245
+ pbswgs = 0.8
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0
+ kt1 = -0.11040563
+ kt2 = -0.048714998
+ lk2 = 3.0890726e-9
+ llc = 0
+ lln = 1
+ lu0 = -1.8172818e-9
+ mjd = 0.335
+ mjs = 0.335
+ lua = -6.2776752e-16
+ lub = 4.4518935e-25
+ luc = 5.1177769e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ igcmod = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 1.0817056e-13
+ wkvth0we = 0.0
+ nsd = 1e+20
+ pbd = 0.75
+ tnoimod = 0
+ pat = 0
+ pbs = 0.75
+ pk2 = -1.5480351e-16
+ eta0 = 0.10792519
+ etab = -0.13555556
+ pu0 = 1.5955157e-16
+ prt = 0
+ pua = 4.4574845e-23
+ pub = -2.7161351e-32
+ puc = -4.8372521e-24
+ pud = 0
+ rsh = 15.2
+ trnqsmod = 0
+ tcj = 0.000832
+ ua1 = 2.771768e-9
+ ub1 = -3.1924567e-18
+ uc1 = -6.2120134e-12
+ cigbinv = 0.006
+ tpb = 0.0016
+ wa0 = -1.0464262e-7
+ ute = -0.78783539
+ pvoff = -9.9175093e-16
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 4.174453e-9
+ wlc = 0
+ wln = 1
+ wu0 = -8.9929205e-11
+ xgl = -8.2e-9
+ xgw = 0
+ wua = -7.0620672e-17
+ wub = -4.621089e-27
+ wuc = 8.8883858e-18
+ wud = 0
+ cdscb = 0
+ cdscd = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ pvsat = 0
+ a0 = 3.3624733
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ wk2we = 0.0
+ pvth0 = 1.7530712e-16
+ at = 72000
+ cf = 8.17e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.013259817
+ k3 = -2.5823
+ em = 20000000.0
+ drout = 0.56
+ version = 4.5
+ ll = 0
+ lw = 0
+ u0 = 0.012618186
+ w0 = 0
+ ua = 4.4026063e-10
+ ub = 1.2150282e-18
+ uc = -4.4814963e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ paigc = 4.1038726e-19
+ xw = 6e-9
+ tempmod = 0
+ voffl = 0
+ rgatemod = 0
+ permod = 1
+ tnjtsswg = 1
+ weta0 = 2.1403289e-9
+ wetab = 2.9133333e-9
+ aigbacc = 0.012071
+ lpclm = 0
+ cgidl = 1
+ voffcv = -0.125
+ wpemod = 1
+ aigbinv = 0.009974
+ pbswd = 0.9
+ pbsws = 0.9
+ keta = -0.035939983
+ pdits = 0
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ lags = -3.1625612e-7
+ tpbswg = 0.001
+ poxedge = 1
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 8.2671111e-11
+ kt1l = 0
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ binunit = 2
+ lint = 6.5375218e-9
+ ptvoff = 8.8703803e-17
+ lkt1 = -6.2138035e-8
+ lkt2 = -3.1463267e-9
+ tnoia = 0
+ lmax = 8.9908e-7
+ waigsd = 1.9716411e-12
+ lmin = 4.4908e-7
+ ijthsfwd = 0.01
+ peta0 = 0
+ lpe0 = 6.44e-8
+ lpeb = 0
+ wketa = 2.5430806e-9
+ diomod = 1
+ tpbsw = 0.0025
+ minv = -0.33
+ lua1 = -1.8157361e-16
+ lub1 = 3.2089876e-25
+ luc1 = 1.2550631e-17
+ pditsd = 0
+ cjswd = 5.1e-11
+ pditsl = 0
+ )

.model pch_tt_36 pmos (
+ level = 54
+ ags = 0.79842724
+ pvfbsdoff = 0
+ wcit = 5.8162887e-11
+ lketa = -1.0850486e-8
+ cigbacc = 0.245
+ cjd = 0.001346
+ cit = -0.00049977211
+ cjs = 0.001346
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ voff = -0.11894985
+ xpart = 1
+ dlc = 1.38228675e-8
+ k3b = 2.1176
+ acde = 0.5
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ rgatemod = 0
+ tnjtsswg = 1
+ vsat = 108525.44
+ tnoimod = 0
+ wint = 0
+ vth0 = -0.39350626
+ egidl = 0.001
+ wkt1 = 8.365112e-10
+ wkt2 = -1.4765978e-9
+ la0 = -3.2362015e-7
+ wmax = 2.7e-7
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0
+ aigc = 0.0068096243
+ wmin = 1.08e-7
+ kt1 = -0.25321364
+ kt2 = -0.04359324
+ lk2 = -3.427309e-10
+ llc = -1.18e-13
+ lln = 0.7
+ cigbinv = 0.006
+ lu0 = -4.5059608e-10
+ mjd = 0.335
+ mjs = 0.335
+ lua = -1.7021816e-16
+ lub = 1.0550853e-25
+ luc = -1.2975077e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ fprout = 200
+ njs = 1.02
+ pa0 = -3.1370244e-14
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ pk2 = 1.4083403e-16
+ xrcrg1 = 12
+ xrcrg2 = 1
+ pu0 = -1.3937081e-17
+ prt = 0
+ pua = 4.7117679e-24
+ pub = -8.7289665e-33
+ puc = -3.0945045e-25
+ pud = 0
+ wua1 = -2.3000717e-16
+ wub1 = 1.2114667e-25
+ wuc1 = -1.9684753e-17
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 2.6350858e-9
+ ub1 = -2.2549964e-18
+ uc1 = 3.1191962e-11
+ bigc = 0.0012521
+ wute = -1.1762912e-7
+ version = 4.5
+ tpb = 0.0016
+ wa0 = 2.1249557e-7
+ wwlc = 0
+ ute = -0.71022675
+ wtvoff = -1.1036076e-10
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 3.5025496e-9
+ tempmod = 0
+ wlc = 0
+ wln = 1
+ wu0 = 3.0436319e-10
+ xgl = -8.2e-9
+ xgw = 0
+ wua = 1.9977231e-17
+ wub = -4.6512873e-26
+ wuc = -1.4020724e-18
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ wtvfbsdoff = 0
+ aigbacc = 0.012071
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigc = 0.15259
+ pvoff = 9.5942711e-17
+ capmod = 2
+ cdscb = 0
+ cdscd = 0
+ wku0we = 1.5e-11
+ pvsat = 0
+ wk2we = 0.0
+ pvth0 = -2.3393785e-16
+ ltvfbsdoff = 0
+ drout = 0.56
+ mobmod = 0
+ paigc = -1.759214e-19
+ aigbinv = 0.009974
+ voffl = 0
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ weta0 = 2.1403289e-9
+ wetab = 2.9133333e-9
+ lpclm = 0
+ k2we = 5e-5
+ ijthsfwd = 0.01
+ cgidl = 1
+ dsub = 0.5
+ ptvfbsdoff = 0
+ dtox = 3.91e-10
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ poxedge = 1
+ eta0 = 0.10792519
+ pbswd = 0.9
+ etab = -0.13555556
+ pbsws = 0.9
+ ijthsrev = 0.01
+ binunit = 2
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ pdits = 0
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ ppdiblc2 = 9.2177422e-17
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ tnoia = 0
+ toxref = 3e-9
+ peta0 = 0
+ wketa = -1.9938172e-9
+ tpbsw = 0.0025
+ cjswd = 5.1e-11
+ cjsws = 5.1e-11
+ pkvth0we = 0.0
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ tvfbsdoff = 0.1
+ ltvoff = -1.9203223e-10
+ vfbsdoff = 0.01
+ njtsswg = 6.489
+ keta = -0.0017391106
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ lags = 9.5750741e-8
+ lku0we = 1.8e-11
+ paramchk = 1
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ scref = 1e-6
+ ckappad = 0.6
+ ckappas = 0.6
+ lcit = 2.6389973e-10
+ pdiblc1 = 0
+ pdiblc2 = 0.016049816
+ epsrox = 3.9
+ pdiblcb = 0
+ pigcd = 2.572
+ kt1l = 0
+ aigsd = 0.0063632396
+ rdsmod = 0
+ lvoff = -5.4343156e-9
+ wvfbsdoff = 0
+ lint = 9.7879675e-9
+ igbmod = 1
+ lvfbsdoff = 0
+ lkt1 = 6.97866e-10
+ lkt2 = -5.3999005e-9
+ lvsat = 0
+ lmax = 4.4908e-7
+ lvth0 = 2.8884329e-9
+ lmin = 2.1577e-7
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ ijthdfwd = 0.01
+ lpe0 = 6.44e-8
+ delta = 0.018814
+ bigbacc = 0.0054401
+ lpeb = 0
+ pbswgd = 0.8
+ laigc = -3.1691048e-11
+ pbswgs = 0.8
+ rnoia = 0
+ rnoib = 0
+ minv = -0.33
+ igcmod = 1
+ lua1 = -1.2143343e-16
+ lub1 = -9.158653e-26
+ luc1 = -3.907118e-18
+ kvth0we = -0.00022
+ ndep = 1e+18
+ lute = -4.5106156e-8
+ pketa = -1.0113644e-15
+ ngate = 1.7e+20
+ lwlc = 0
+ lintnoi = -5e-9
+ moin = 5.5538
+ ijthdrev = 0.01
+ ngcon = 1
+ bigbinv = 0.00149
+ wpclm = 7.1298978e-9
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ nigc = 2.291
+ lpdiblc2 = -1.262443e-9
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ pags = 5.2660461e-14
+ permod = 1
+ ntox = 1
+ pcit = -2.559167e-17
+ pclm = 1.101657
+ phin = 0.15
+ lkvth0we = 3e-12
+ pkt1 = -5.70475e-17
+ pkt2 = 1.4763857e-16
+ voffcv = -0.125
+ wpemod = 1
+ tvoff = 0.0020889601
+ nfactor = 1
+ xjbvd = 1
+ acnqsmod = 0
+ xjbvs = 1
+ lk2we = 0.0
+ a0 = 1.7239078
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ rbdb = 50
+ pua1 = 1.9443948e-23
+ prwb = 0
+ pub1 = 1.2643651e-32
+ prwg = 0
+ at = 72000
+ puc1 = 5.3837292e-24
+ cf = 8.17e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.0054602636
+ k3 = -2.5823
+ em = 20000000.0
+ rbpb = 50
+ rbpd = 50
+ ll = -1.18e-13
+ lw = 0
+ rbps = 50
+ u0 = 0.009512082
+ rbsb = 50
+ pvag = 2.1
+ w0 = 0
+ rbodymod = 0
+ ua = -5.9962427e-10
+ ub = 1.98703e-18
+ uc = 1.0098696e-10
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ pute = 2.0393808e-14
+ xw = 6e-9
+ rdsw = 200
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = 0
+ nigbacc = 10
+ ppclm = 0
+ tpbswg = 0.001
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ rshg = 14.1
+ nigbinv = 2.171
+ wpdiblc2 = -7.8646151e-10
+ ptvoff = 3.6984079e-17
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ waigsd = 1.9716411e-12
+ diomod = 1
+ fnoimod = 1
+ pditsd = 0
+ pditsl = 0
+ bigsd = 0.0003327
+ cjswgd = 1.81e-10
+ pku0we = 0.0
+ tnom = 25
+ cjswgs = 1.81e-10
+ eigbinv = 1.1
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ wkvth0we = 0.0
+ wvoff = 1.0046111e-9
+ trnqsmod = 0
+ wvsat = -0.0013318206
+ mjswgd = 0.95
+ wvth0 = -1.621551e-9
+ mjswgs = 0.95
+ tcjswg = 0.00128
+ waigc = 4.0429874e-12
+ wags = 9.7102189e-10
+ )

.model pch_tt_37 pmos (
+ level = 54
+ fprout = 200
+ lvth0 = 5.5274905e-9
+ xrcrg1 = 12
+ xrcrg2 = 1
+ delta = 0.018814
+ wtvfbsdoff = 0
+ laigc = -4.357169e-12
+ rnoia = 0
+ rnoib = 0
+ acnqsmod = 0
+ wtvoff = 1.2048366e-10
+ ltvfbsdoff = 0
+ pketa = 4.1278959e-16
+ ngate = 1.7e+20
+ rbodymod = 0
+ ngcon = 1
+ wpclm = 6.8691006e-8
+ capmod = 2
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ wku0we = 1.5e-11
+ keta = -0.058692164
+ mobmod = 0
+ nfactor = 1
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 2.5291477e-11
+ ptvfbsdoff = 0
+ kt1l = 0
+ wpdiblc2 = -7.28246e-10
+ lint = 9.7879675e-9
+ lkt1 = -4.6770694e-9
+ lkt2 = -3.7791597e-9
+ lmax = 2.1577e-7
+ lmin = 9e-8
+ lpe0 = 6.44e-8
+ nigbacc = 10
+ lpeb = 0
+ tvoff = 0.0011827459
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ minv = -0.33
+ lua1 = -2.1218464e-16
+ lub1 = 2.7818737e-25
+ luc1 = 2.2554944e-17
+ ndep = 1e+18
+ wkvth0we = 0.0
+ lute = 1.5508066e-9
+ lwlc = 0
+ moin = 5.5538
+ nigbinv = 2.171
+ ku0we = -0.0007
+ trnqsmod = 0
+ beta0 = 13.32
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ nigc = 2.291
+ leta0 = 0
+ ppclm = -1.2989269e-14
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ fnoimod = 1
+ eigbinv = 1.1
+ ntox = 1
+ rgatemod = 0
+ pcit = 1.1214196e-17
+ pclm = 0.85425247
+ tnjtsswg = 1
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ phin = 0.15
+ toxref = 3e-9
+ pkt1 = -2.317336e-16
+ pkt2 = 3.7767926e-16
+ bigsd = 0.0003327
+ cigbacc = 0.245
+ rbdb = 50
+ pua1 = 2.6827919e-23
+ prwb = 0
+ pub1 = -3.4278711e-32
+ prwg = 0
+ puc1 = -2.7535024e-24
+ wvoff = 8.5374562e-10
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ pute = -4.2802262e-16
+ ltvoff = -8.1627e-13
+ rdsw = 200
+ tnoimod = 0
+ wvsat = -0.00089129698
+ ags = 1.2522222
+ wvth0 = -2.650948e-9
+ cjd = 0.001346
+ cit = 0.00063107268
+ cjs = 0.001346
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 1.38228675e-8
+ waigc = 1.4660694e-11
+ k3b = 2.1176
+ cigbinv = 0.006
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ pvfbsdoff = 0
+ lku0we = 1.8e-11
+ lketa = 1.1666086e-9
+ epsrox = 3.9
+ la0 = 6.219346e-9
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = -0.0075443287
+ xpart = 1
+ kt1 = -0.22773883
+ kt2 = -0.051274476
+ lk2 = 3.6711471e-9
+ llc = -1.18e-13
+ lln = 0.7
+ lu0 = -1.6314862e-10
+ mjd = 0.335
+ version = 4.5
+ mjs = 0.335
+ lua = 1.3101868e-17
+ lub = -8.7271368e-26
+ luc = -1.2812174e-17
+ lud = 0
+ rshg = 14.1
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = -2.0637395e-14
+ rdsmod = 0
+ nsd = 1e+20
+ pbd = 0.75
+ tempmod = 0
+ pat = -5.0045721e-10
+ pbs = 0.75
+ pk2 = 4.0368065e-17
+ egidl = 0.001
+ igbmod = 1
+ pu0 = -5.2679707e-18
+ prt = 0
+ pua = -4.0286539e-24
+ pub = 7.5106005e-33
+ puc = 1.4358513e-24
+ pud = 0
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 3.0651863e-9
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ ub1 = -4.0074881e-18
+ uc1 = -9.4220652e-11
+ tpb = 0.0016
+ aigbacc = 0.012071
+ wa0 = 1.6162969e-7
+ pbswgd = 0.8
+ pbswgs = 0.8
+ ute = -0.93134979
+ ijthsfwd = 0.01
+ wat = 0.0023718351
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 3.9786916e-9
+ wlc = 0
+ wln = 1
+ wu0 = 2.6327735e-10
+ xgl = -8.2e-9
+ xgw = 0
+ wua = 6.1401032e-17
+ wub = -1.2347765e-25
+ wuc = -9.6736445e-18
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ igcmod = 1
+ tnom = 25
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ aigbinv = 0.009974
+ ijthsrev = 0.01
+ pvoff = 1.2777532e-16
+ cdscb = 0
+ cdscd = 0
+ pvsat = -9.2948987e-11
+ wags = 2.5054667e-7
+ wk2we = 0.0
+ pvth0 = -1.6735092e-17
+ drout = 0.56
+ wcit = -1.162725e-10
+ paigc = -2.4162575e-18
+ permod = 1
+ voff = -0.1339517
+ acde = 0.5
+ ppdiblc2 = 7.9894307e-17
+ voffl = 0
+ poxedge = 1
+ vsat = 106518.57
+ wint = 0
+ vth0 = -0.40601365
+ weta0 = 2.1403289e-9
+ wetab = 2.9133333e-9
+ wkt1 = 1.664079e-9
+ wkt2 = -2.566838e-9
+ wmax = 2.7e-7
+ lpclm = 5.2201277e-8
+ binunit = 2
+ aigc = 0.0066800799
+ wmin = 1.08e-7
+ voffcv = -0.125
+ wpemod = 1
+ cgidl = 1
+ wua1 = -2.6500229e-16
+ wub1 = 3.4352994e-25
+ wuc1 = 1.8880326e-17
+ bigc = 0.0012521
+ wute = -1.8947457e-8
+ pkvth0we = 0.0
+ wwlc = 0
+ pbswd = 0.9
+ pbsws = 0.9
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ vfbsdoff = 0.01
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigc = 0.15259
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ pdits = 0
+ tpbswg = 0.001
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ paramchk = 1
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ ptvoff = -1.1725409e-17
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ a0 = 0.16068118
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ waigsd = 1.9716411e-12
+ at = 107755.11
+ cf = 8.17e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.024483382
+ k3 = -2.5823
+ em = 20000000.0
+ ll = -1.18e-13
+ lw = 0
+ u0 = 0.0081497718
+ tnoia = 0
+ w0 = 0
+ ua = -1.4684396e-9
+ ub = 2.9006788e-18
+ uc = 1.0021491e-10
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 6e-9
+ diomod = 1
+ k2we = 5e-5
+ ijthdfwd = 0.01
+ peta0 = 0
+ njtsswg = 6.489
+ dsub = 0.5
+ dtox = 3.91e-10
+ wketa = -8.743362e-9
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.81e-10
+ pku0we = 0.0
+ cjswgs = 1.81e-10
+ tpbsw = 0.0025
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ cjswd = 5.1e-11
+ cjsws = 5.1e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.01690182
+ eta0 = 0.10792519
+ pdiblcb = 0
+ etab = -0.13555556
+ tvfbsdoff = 0.1
+ ijthdrev = 0.01
+ mjswgd = 0.95
+ mjswgs = 0.95
+ lpdiblc2 = -1.4422174e-9
+ tcjswg = 0.00128
+ bigbacc = 0.0054401
+ scref = 1e-6
+ pigcd = 2.572
+ aigsd = 0.0063632396
+ kvth0we = -0.00022
+ wvfbsdoff = 0
+ lvoff = -2.268926e-9
+ lintnoi = -5e-9
+ lvfbsdoff = 0
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ lkvth0we = 3e-12
+ lvsat = 0.00042343719
+ )

.model pch_tt_38 pmos (
+ level = 54
+ poxedge = 1
+ ptvfbsdoff = 0
+ rdsw = 200
+ capmod = 2
+ vfbsdoff = 0.01
+ wku0we = 1.5e-11
+ pvoff = -1.4373467e-16
+ binunit = 2
+ cdscb = 0
+ cdscd = 0
+ mobmod = 0
+ pvsat = 1.729604e-10
+ wk2we = 0.0
+ pvth0 = 5.6763134e-17
+ drout = 0.56
+ paramchk = 1
+ paigc = -1.1563004e-18
+ voffl = 0
+ rshg = 14.1
+ weta0 = 1.2957501e-8
+ wetab = 4.1458967e-9
+ lpclm = -1.0127779e-7
+ ijthdfwd = 0.01
+ jtsswgd = 1.75e-7
+ cgidl = 1
+ jtsswgs = 1.75e-7
+ tnom = 25
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ pbswd = 0.9
+ pbsws = 0.9
+ ijthdrev = 0.01
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ lpdiblc2 = -1.4113545e-11
+ pdits = 0
+ cigsd = 0.013281
+ wags = 2.5054667e-7
+ dvt0w = 0
+ dvt1w = 0
+ njtsswg = 6.489
+ dvt2w = 0
+ wcit = 7.0487744e-11
+ xtsswgd = 0.32
+ voff = -0.14478455
+ xtsswgs = 0.32
+ acde = 0.5
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ ckappad = 0.6
+ ckappas = 0.6
+ vsat = 137363.5
+ wint = 0
+ pdiblc1 = 0
+ pdiblc2 = 0.0017092259
+ vth0 = -0.34280653
+ pdiblcb = 0
+ wkt1 = -1.350742e-8
+ wkt2 = 1.8825744e-9
+ toxref = 3e-9
+ wmax = 2.7e-7
+ lkvth0we = 3e-12
+ aigc = 0.0067219883
+ wmin = 1.08e-7
+ tnoia = 0
+ peta0 = -1.0168142e-15
+ petab = -1.1586096e-16
+ wketa = -6.6698086e-9
+ wua1 = 1.6631395e-16
+ wub1 = -2.121384e-25
+ wuc1 = 2.5860689e-17
+ tpbsw = 0.0025
+ acnqsmod = 0
+ bigbacc = 0.0054401
+ cjswd = 5.1e-11
+ bigc = 0.0012521
+ cjsws = 5.1e-11
+ wute = -6.1363432e-8
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ wwlc = 0
+ tvfbsdoff = 0.1
+ ltvoff = 3.7319947e-11
+ rbodymod = 0
+ kvth0we = -0.00022
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ lintnoi = -5e-9
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ bigbinv = 0.00149
+ cigc = 0.15259
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ lku0we = 1.8e-11
+ epsrox = 3.9
+ scref = 1e-6
+ pigcd = 2.572
+ aigsd = 0.0063632396
+ rdsmod = 0
+ wpdiblc2 = 8.0253658e-11
+ igbmod = 1
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ lvoff = -1.2506377e-9
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ lvsat = -0.0024759865
+ pbswgd = 0.8
+ pbswgs = 0.8
+ lvth0 = -4.139787e-10
+ k2we = 5e-5
+ delta = 0.018814
+ laigc = -8.2965642e-12
+ dsub = 0.5
+ igcmod = 1
+ dtox = 3.91e-10
+ rnoia = 0
+ rnoib = 0
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ nfactor = 1
+ wkvth0we = 0.0
+ pketa = 2.1787556e-16
+ ngate = 1.7e+20
+ eta0 = 0.024468866
+ etab = -0.22797789
+ ngcon = 1
+ wpclm = -1.6917696e-7
+ trnqsmod = 0
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ nigbacc = 10
+ permod = 1
+ rgatemod = 0
+ tnjtsswg = 1
+ nigbinv = 2.171
+ voffcv = -0.125
+ wpemod = 1
+ tvoff = 0.00077704148
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ fnoimod = 1
+ eigbinv = 1.1
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = 7.844894e-9
+ letab = 8.6876992e-9
+ tpbswg = 0.001
+ ppclm = 9.3703198e-15
+ keta = -0.049241031
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 1.2730569e-10
+ kt1l = 0
+ ptvoff = 1.952106e-17
+ cigbacc = 0.245
+ waigsd = 1.9716411e-12
+ dmcgt = 0
+ lint = 0
+ tcjsw = 9.34e-5
+ tnoimod = 0
+ lkt1 = -6.5946074e-9
+ lkt2 = 9.2375447e-10
+ diomod = 1
+ lmax = 9e-8
+ lmin = 5.4e-8
+ ijthsfwd = 0.01
+ lpe0 = 6.44e-8
+ pditsd = 0
+ pditsl = 0
+ lpeb = 0
+ cigbinv = 0.006
+ cjswgd = 1.81e-10
+ pku0we = 0.0
+ cjswgs = 1.81e-10
+ bigsd = 0.0003327
+ minv = -0.33
+ ags = 1.2522222
+ lua1 = 1.5814311e-16
+ lub1 = -2.3663254e-25
+ luc1 = 3.1466117e-17
+ cjd = 0.001346
+ cit = -0.00045418481
+ cjs = 0.001346
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ ndep = 1e+18
+ bvs = 8.2
+ lute = -1.2895214e-8
+ dlc = 4.0349e-9
+ wvoff = 3.7421498e-9
+ k3b = 2.1176
+ lwlc = 0
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ version = 4.5
+ moin = 5.5538
+ mjswgd = 0.95
+ mjswgs = 0.95
+ ijthsrev = 0.01
+ tempmod = 0
+ wvsat = -0.0037201203
+ nigc = 2.291
+ tcjswg = 0.00128
+ wvth0 = -3.432844e-9
+ la0 = 3.4503642e-8
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = -0.0080528059
+ kt1 = -0.20733948
+ kt2 = -0.10130548
+ lk2 = 5.547863e-9
+ waigc = 1.256895e-12
+ llc = 0
+ lln = 1
+ a0 = -0.1402156
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ lu0 = 4.580914e-11
+ mjd = 0.335
+ mjs = 0.335
+ lua = 1.1003971e-16
+ lub = -1.3258131e-25
+ luc = -1.072064e-17
+ at = 113164.44
+ lud = 0
+ cf = 8.17e-11
+ lwc = 0
+ pvfbsdoff = 0
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.044448444
+ k3 = -2.5823
+ lwl = 0
+ lwn = 1
+ em = 20000000.0
+ aigbacc = 0.012071
+ njd = 1.02
+ njs = 1.02
+ ll = 0
+ noff = 2.2684
+ pa0 = -6.959911e-15
+ lw = 0
+ u0 = 0.0059268169
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ w0 = 0
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 1.1859675e-9
+ ua = -2.4996932e-9
+ ub = 3.3826995e-18
+ uc = 7.7964547e-11
+ ud = 0
+ pbs = 0.75
+ pk2 = -8.547569e-17
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 6e-9
+ pu0 = 1.7354187e-18
+ prt = 0
+ lketa = 2.7820203e-10
+ pua = -5.4706466e-24
+ pub = 7.2761107e-33
+ puc = 2.7207836e-25
+ pud = 0
+ wtvfbsdoff = 0
+ xpart = 1
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = -8.7447052e-10
+ ub1 = 1.4693195e-18
+ uc1 = -1.8902037e-10
+ ppdiblc2 = 3.8953385e-18
+ ntox = 1
+ tpb = 0.0016
+ pcit = -6.3412667e-18
+ pclm = 2.4870084
+ wa0 = 1.612455e-8
+ ute = -0.77766872
+ wat = -0.015568853
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 5.3174549e-9
+ aigbinv = 0.009974
+ wlc = 0
+ egidl = 0.001
+ wln = 1
+ wu0 = 1.8877321e-10
+ xgl = -8.2e-9
+ xgw = 0
+ wua = 7.6741379e-17
+ wub = -1.2098307e-25
+ wuc = 2.7069183e-18
+ wud = 0
+ wwc = 0
+ ltvfbsdoff = 0
+ wwl = 0
+ wwn = 1
+ phin = 0.15
+ fprout = 200
+ xrcrg1 = 12
+ xrcrg2 = 1
+ pkt1 = 1.1943873e-15
+ pkt2 = -4.056551e-17
+ wtvoff = -2.1192558e-10
+ pkvth0we = 0.0
+ rbdb = 50
+ pua1 = -1.3715808e-23
+ prwb = 0
+ pub1 = 1.7954113e-32
+ prwg = 0
+ puc1 = -3.4096566e-24
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ pute = 3.5590791e-15
+ )

.model pch_tt_39 pmos (
+ level = 54
+ fnoimod = 1
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ eigbinv = 1.1
+ k2we = 5e-5
+ ijthsfwd = 0.01
+ tvoff = 0.00092289205
+ dsub = 0.5
+ dtox = 3.91e-10
+ xjbvd = 1
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ xjbvs = 1
+ lk2we = 0.0
+ eta0 = 0.19463541
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ etab = -0.16706384
+ ijthsrev = 0.01
+ cigbacc = 0.245
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = -2.0247657e-9
+ letab = 5.1546845e-9
+ tnoimod = 0
+ ppclm = 7.8094068e-15
+ dlcig = 2.5e-9
+ cigbinv = 0.006
+ bgidl = 1834800000.0
+ ppdiblc2 = 0
+ toxref = 3e-9
+ version = 4.5
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ tempmod = 0
+ ags = 1.2522222
+ cjd = 0.001346
+ cit = -0.0026753087
+ cjs = 0.001346
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 4.0349e-9
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ aigbacc = 0.012071
+ bigsd = 0.0003327
+ pkvth0we = 0.0
+ la0 = -1.4904033e-7
+ ltvoff = 2.8860613e-11
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0.009372509
+ kt1 = -0.53950997
+ kt2 = -0.12590838
+ lk2 = 4.2165993e-9
+ wvoff = 1.4341134e-10
+ llc = 0
+ lln = 1
+ lu0 = 4.1651089e-10
+ mjd = 0.335
+ mjs = 0.335
+ lua = 7.9060667e-17
+ lub = -2.7964918e-26
+ luc = 5.5424848e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = -2.574678e-15
+ nsd = 1e+20
+ pbd = 0.75
+ pat = -1.0212358e-9
+ wvsat = -0.0027183681
+ pbs = 0.75
+ pk2 = 2.1304022e-16
+ aigbinv = 0.009974
+ wvth0 = -2.182128e-9
+ pu0 = -6.6237547e-17
+ vfbsdoff = 0.01
+ prt = 0
+ pua = -2.0419953e-23
+ pub = 1.469069e-32
+ puc = 1.2609666e-24
+ pud = 0
+ waigc = 6.0357037e-12
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 8.3453493e-9
+ ub1 = -1.1410668e-17
+ pvfbsdoff = 0
+ uc1 = 1.6197295e-9
+ keta = -0.31465021
+ lku0we = 1.8e-11
+ tpb = 0.0016
+ wa0 = -5.9482929e-8
+ epsrox = 3.9
+ ute = -1
+ wat = 0.022486376
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 1.7062889e-10
+ wlc = 0
+ wln = 1
+ wu0 = 1.3607209e-9
+ xgl = -8.2e-9
+ xgw = 0
+ wua = 3.3448805e-16
+ wub = -2.4882066e-25
+ wuc = -1.434288e-17
+ wud = 0
+ lketa = 1.5671934e-8
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ paramchk = 1
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 2.5613086e-10
+ xpart = 1
+ rdsmod = 0
+ kt1l = 0
+ igbmod = 1
+ egidl = 0.001
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ lint = 0
+ poxedge = 1
+ pbswgd = 0.8
+ pbswgs = 0.8
+ lkt1 = 1.2671281e-8
+ lkt2 = 2.350723e-9
+ lmax = 5.4e-8
+ lmin = 4.5e-8
+ ijthdfwd = 0.01
+ igcmod = 1
+ binunit = 2
+ lpe0 = 6.44e-8
+ lpeb = 0
+ minv = -0.33
+ lua1 = -3.7660644e-16
+ lub1 = 5.1040674e-25
+ luc1 = -7.3441373e-17
+ ndep = 1e+18
+ lwlc = 0
+ ijthdrev = 0.01
+ moin = 5.5538
+ nigc = 2.291
+ lpdiblc2 = 0
+ pvoff = 6.4992158e-17
+ cdscb = 0
+ cdscd = 0
+ pvsat = 1.1485877e-10
+ noff = 2.2684
+ wk2we = 0.0
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ pvth0 = -1.5778397e-17
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ permod = 1
+ drout = 0.56
+ paigc = -1.4334713e-18
+ voffl = 0
+ ntox = 1
+ pcit = -1.8399318e-17
+ pclm = 1.8533357
+ weta0 = -4.6483037e-9
+ wetab = 2.5894049e-9
+ lpclm = -6.4524768e-8
+ lkvth0we = 3e-12
+ phin = 0.15
+ voffcv = -0.125
+ wpemod = 1
+ pkt1 = -1.7183146e-15
+ pkt2 = -1.1786798e-16
+ cgidl = 1
+ acnqsmod = 0
+ njtsswg = 6.489
+ rbdb = 50
+ pua1 = 1.8341764e-23
+ prwb = 0
+ pub1 = -1.3009877e-32
+ prwg = 0
+ puc1 = 9.9681375e-24
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ pbswd = 0.9
+ rbpb = 50
+ rbpd = 50
+ pbsws = 0.9
+ rbps = 50
+ rbodymod = 0
+ rbsb = 50
+ pvag = 2.1
+ ckappad = 0.6
+ ckappas = 0.6
+ rdsw = 200
+ pdiblc1 = 0
+ pdiblc2 = 0.0014658889
+ pdiblcb = 0
+ tpbswg = 0.001
+ pdits = 0
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ bigbacc = 0.0054401
+ ptvoff = -2.2999757e-17
+ pk2we = 0.0
+ wpdiblc2 = 1.4741467e-10
+ rshg = 14.1
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ waigsd = 1.9716411e-12
+ kvth0we = -0.00022
+ diomod = 1
+ tnoia = 0
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ pditsd = 0
+ pditsl = 0
+ vtsswgd = 1.1
+ peta0 = 4.3224906e-18
+ vtsswgs = 1.1
+ cjswgd = 1.81e-10
+ pku0we = 0.0
+ cjswgs = 1.81e-10
+ petab = -2.558443e-17
+ wketa = 3.409679e-8
+ tpbsw = 0.0025
+ tnom = 25
+ cjswd = 5.1e-11
+ cjsws = 5.1e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ tvfbsdoff = 0.1
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ wkvth0we = 0.0
+ mjswgd = 0.95
+ mjswgs = 0.95
+ wtvfbsdoff = 0
+ tcjswg = 0.00128
+ trnqsmod = 0
+ ltvfbsdoff = 0
+ wags = 2.5054667e-7
+ wcit = 2.7838518e-10
+ scref = 1e-6
+ voff = -0.1005239
+ pigcd = 2.572
+ acde = 0.5
+ aigsd = 0.0063632396
+ nfactor = 1
+ rgatemod = 0
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ tnjtsswg = 1
+ vsat = 101849.16
+ wint = 0
+ lvoff = -3.8177557e-9
+ vth0 = -0.27314034
+ fprout = 200
+ wkt1 = 3.6711578e-8
+ wkt2 = 3.2153756e-9
+ wmax = 2.7e-7
+ xrcrg1 = 12
+ xrcrg2 = 1
+ aigc = 0.0068691843
+ wmin = 1.08e-7
+ lvsat = -0.00041615496
+ lvth0 = -4.4546177e-9
+ ptvfbsdoff = 0
+ delta = 0.018814
+ laigc = -1.683393e-11
+ wtvoff = 5.2119196e-10
+ wua1 = -3.864028e-16
+ wub1 = 3.2172349e-25
+ wuc1 = -2.0479093e-16
+ rnoia = 0
+ rnoib = 0
+ a0 = 3.0243356
+ a1 = 0
+ a2 = 1
+ nigbacc = 10
+ b0 = 0
+ b1 = 0
+ at = -187272.02
+ cf = 8.17e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.021495622
+ k3 = -2.5823
+ em = 20000000.0
+ bigc = 0.0012521
+ ll = 0
+ lw = 0
+ u0 = -0.00046459259
+ w0 = 0
+ wwlc = 0
+ ua = -1.9655718e-9
+ ub = 1.5789686e-18
+ uc = -2.0243416e-10
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 6e-9
+ pketa = -2.1465872e-15
+ ngate = 1.7e+20
+ ngcon = 1
+ capmod = 2
+ wpclm = -1.4226467e-7
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ wku0we = 1.5e-11
+ xtid = 3
+ xtis = 3
+ gbmin = 1e-12
+ nigbinv = 2.171
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigc = 0.15259
+ jswgd = 3.69e-13
+ mobmod = 0
+ jswgs = 3.69e-13
+ )

.model pch_tt_40 pmos (
+ level = 54
+ fnoimod = 1
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ eigbinv = 1.1
+ laigsd = 6.1219753e-16
+ k2we = 5e-5
+ ijthsfwd = 0.01
+ tvoff = -0.00058332606
+ dsub = 0.5
+ dtox = 3.91e-10
+ xjbvd = 1
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ xjbvs = 1
+ lk2we = 0.0
+ eta0 = 0.11700471
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ etab = -0.15063456
+ ijthsrev = 0.01
+ cigbacc = 0.245
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = 1.7791389e-9
+ letab = 4.3496496e-9
+ tnoimod = 0
+ ppclm = -3.5647768e-15
+ dlcig = 2.5e-9
+ cigbinv = 0.006
+ bgidl = 1834800000.0
+ ppdiblc2 = 0
+ toxref = 3e-9
+ version = 4.5
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ tempmod = 0
+ ags = 1.2522222
+ cjd = 0.001346
+ cit = -0.0077632099
+ cjs = 0.001346
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 4.0349e-9
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ aigbacc = 0.012071
+ bigsd = 0.0003327
+ pkvth0we = 0.0
+ la0 = -3.4726683e-8
+ ltvoff = 1.026653e-10
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0.0017111307
+ kt1 = -0.31430817
+ kt2 = -0.12562663
+ lk2 = 6.2841473e-9
+ wvoff = 3.3909703e-9
+ llc = 0
+ lln = 1
+ lu0 = 5.2641728e-10
+ mjd = 0.335
+ mjs = 0.335
+ lua = 9.0470184e-17
+ lub = -1.3836274e-26
+ luc = 2.7216576e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 1.4761752e-15
+ nsd = 1e+20
+ pbd = 0.75
+ pat = -5.6834015e-11
+ wvsat = -0.010288162
+ pbs = 0.75
+ pk2 = -2.7720832e-16
+ aigbinv = 0.009974
+ wvth0 = 1.3037359e-10
+ pu0 = -6.1923224e-17
+ vfbsdoff = 0.01
+ prt = 0
+ pua = -4.2432063e-24
+ pub = -6.6397485e-33
+ puc = -1.7176927e-24
+ pud = 0
+ waigc = -4.0606639e-11
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 2.1566906e-9
+ ub1 = -3.7269546e-18
+ pvfbsdoff = 0
+ uc1 = -1.7258848e-10
+ keta = 0.15497942
+ lku0we = 1.8e-11
+ tpb = 0.0016
+ wa0 = -1.421534e-7
+ epsrox = 3.9
+ ute = -1
+ wat = 0.002804707
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 1.0175701e-8
+ wlc = 0
+ wln = 1
+ wu0 = 1.2726735e-9
+ xgl = -8.2e-9
+ xgw = 0
+ wua = 4.3503521e-18
+ wub = 1.8649442e-25
+ wuc = 4.6446086e-17
+ wud = 0
+ lketa = -7.3399177e-9
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ paramchk = 1
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 5.0543803e-10
+ xpart = 1
+ rdsmod = 0
+ kt1l = 0
+ igbmod = 1
+ egidl = 0.001
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ lint = 0
+ poxedge = 1
+ pbswgd = 0.8
+ pbswgs = 0.8
+ lkt1 = 1.6363929e-9
+ lkt2 = 2.3369169e-9
+ lmax = 4.5e-8
+ lmin = 3.6e-8
+ ijthdfwd = 0.01
+ igcmod = 1
+ binunit = 2
+ lpe0 = 6.44e-8
+ lpeb = 0
+ minv = -0.33
+ lua1 = -7.3362164e-17
+ lub1 = 1.3390478e-25
+ luc1 = 1.4382206e-17
+ ndep = 1e+18
+ lwlc = 0
+ ijthdrev = 0.01
+ moin = 5.5538
+ nigc = 2.291
+ paigsd = -6.9790518e-23
+ lpdiblc2 = 0
+ pvoff = -9.4138231e-17
+ cdscb = 0
+ cdscd = 0
+ pvsat = 4.8577866e-10
+ noff = 2.2684
+ wk2we = 0.0
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ pvth0 = -1.2909097e-16
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ permod = 1
+ drout = 0.56
+ paigc = 8.520035e-19
+ voffl = 0
+ ntox = 1
+ pcit = -1.9287562e-17
+ pclm = 0.41497396
+ weta0 = -1.275677e-9
+ wetab = 1.1541057e-8
+ lpclm = 5.9549575e-9
+ lkvth0we = 3e-12
+ phin = 0.15
+ voffcv = -0.125
+ wpemod = 1
+ pkt1 = -1.7140714e-15
+ pkt2 = -7.0509572e-16
+ cgidl = 1
+ acnqsmod = 0
+ njtsswg = 6.489
+ rbdb = 50
+ pua1 = 3.2441676e-23
+ prwb = 0
+ pub1 = -5.4663004e-32
+ prwg = 0
+ puc1 = -1.3788915e-24
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ pbswd = 0.9
+ rbpb = 50
+ rbpd = 50
+ pbsws = 0.9
+ rbps = 50
+ rbodymod = 0
+ rbsb = 50
+ pvag = 2.1
+ ckappad = 0.6
+ ckappas = 0.6
+ rdsw = 200
+ pdiblc1 = 0
+ pdiblc2 = 0.0014658889
+ pdiblcb = 0
+ tpbswg = 0.001
+ pdits = 0
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ bigbacc = 0.0054401
+ ptvoff = -3.9364956e-17
+ pk2we = 0.0
+ wpdiblc2 = 1.4741467e-10
+ rshg = 14.1
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ waigsd = 1.9730654e-12
+ kvth0we = -0.00022
+ diomod = 1
+ tnoia = 0
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ pditsd = 0
+ pditsl = 0
+ vtsswgd = 1.1
+ peta0 = -1.6093622e-16
+ vtsswgs = 1.1
+ cjswgd = 1.81e-10
+ pku0we = 0.0
+ cjswgs = 1.81e-10
+ petab = -4.6421536e-16
+ wketa = -5.7187654e-8
+ tpbsw = 0.0025
+ tnom = 25
+ cjswd = 5.1e-11
+ cjsws = 5.1e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ tvfbsdoff = 0.1
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ wkvth0we = 0.0
+ mjswgd = 0.95
+ mjswgs = 0.95
+ wtvfbsdoff = 0
+ tcjswg = 0.00128
+ trnqsmod = 0
+ ltvfbsdoff = 0
+ wags = 2.5054667e-7
+ wcit = 2.9651259e-10
+ scref = 1e-6
+ voff = -0.12231559
+ pigcd = 2.572
+ acde = 0.5
+ aigsd = 0.0063632271
+ nfactor = 1
+ rgatemod = 0
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ tnjtsswg = 1
+ vsat = 151791.98
+ wint = 0
+ lvoff = -2.7499629e-9
+ vth0 = -0.33708607
+ fprout = 200
+ wkt1 = 3.6624982e-8
+ wkt2 = 1.5199615e-8
+ wmax = 2.7e-7
+ xrcrg1 = 12
+ xrcrg2 = 1
+ aigc = 0.0069354083
+ wmin = 1.08e-7
+ lvsat = -0.0028633534
+ lvth0 = -1.3212769e-9
+ ptvfbsdoff = 0
+ delta = 0.018814
+ laigc = -2.0078906e-11
+ wtvoff = 8.5517561e-10
+ wua1 = -6.7415611e-16
+ wub1 = 1.1717873e-24
+ wuc1 = 2.6781086e-17
+ rnoia = 0
+ rnoib = 0
+ a0 = 0.69140412
+ a1 = 0
+ a2 = 1
+ nigbacc = 10
+ b0 = 0
+ b1 = 0
+ at = -30917.36
+ cf = 8.17e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.06369048
+ k3 = -2.5823
+ em = 20000000.0
+ bigc = 0.0012521
+ ll = 0
+ lw = 0
+ u0 = -0.0027075803
+ w0 = 0
+ wwlc = 0
+ ua = -2.1984191e-9
+ ub = 1.2906289e-18
+ uc = -1.4486626e-10
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 6e-9
+ pketa = 2.3263506e-15
+ ngate = 1.7e+20
+ ngcon = 1
+ capmod = 2
+ wpclm = 8.9861524e-8
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ wku0we = 1.5e-11
+ xtid = 3
+ xtis = 3
+ gbmin = 1e-12
+ nigbinv = 2.171
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigc = 0.15259
+ jswgd = 3.69e-13
+ mobmod = 0
+ jswgs = 3.69e-13
+ )

.model pch_ff_1 pmos (
+ level = 54
+ ppclm = 0
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ bigbacc = 0.0054401
+ wpdiblc2 = 0
+ tnom = 25
+ kvth0we = -0.00022
+ tvfbsdoff = 0.1
+ dmcgt = 0
+ toxe = 2.6300000000000002e-9
+ toxm = 2.67e-9
+ tcjsw = 9.34e-5
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ toxref = 3e-9
+ bigsd = 0.0003327
+ wkvth0we = 0.0
+ wvoff = 0
+ trnqsmod = 0
+ voff = -0.11110337
+ acde = 0.5
+ wvsat = 0
+ wvfbsdoff = 0
+ wvth0 = 2.7e-9
+ lvfbsdoff = 0
+ vsat = 120000
+ wint = 0
+ vth0 = -0.36413527
+ ltvoff = 0
+ wmax = 0.00090001
+ aigc = 0.0068307507
+ wmin = 8.9974e-6
+ a0 = 2.531
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 72000
+ cf = 8.741900000000001e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.00077592763
+ k3 = -2.5823
+ em = 20000000.0
+ lketa = 0
+ ll = 0
+ lw = 0
+ u0 = 0.009505
+ w0 = 0
+ rgatemod = 0
+ ua = 1.297e-10
+ ub = 1.182572e-18
+ uc = 2.014e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 2.33e-9
+ ww = 0
+ xpart = 1
+ xw = 8.600000000000001e-9
+ nfactor = 1
+ tnjtsswg = 1
+ lku0we = 1.8e-11
+ bigc = 0.0012521
+ egidl = 0.001
+ wwlc = 0
+ epsrox = 3.9
+ cdsc = 0
+ rdsmod = 0
+ cgbo = 0
+ cgdl = 3.2212350000000004e-11
+ cgdo = 2.8335740000000002e-11
+ xtid = 3
+ xtis = 3
+ igbmod = 1
+ cgsl = 3.2212350000000004e-11
+ cgso = 2.8335740000000002e-11
+ cigc = 0.15259
+ nigbacc = 10
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ pbswgd = 0.8
+ pbswgs = 0.8
+ igcmod = 1
+ nigbinv = 2.171
+ pvoff = -2.5e-17
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ cdscb = 0
+ cdscd = 0
+ pvsat = 0
+ wk2we = 0.0
+ pvth0 = 1.5e-16
+ drout = 0.56
+ k2we = 5e-5
+ dsub = 0.5
+ dtox = 3.91e-10
+ voffl = 0
+ fnoimod = 1
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ eigbinv = 1.1
+ weta0 = 2.8e-10
+ permod = 1
+ lpclm = 0
+ eta0 = 0.1672
+ etab = -0.23
+ ijthsfwd = 0.01
+ cgidl = 1
+ voffcv = -0.125
+ wpemod = 1
+ ijthsrev = 0.01
+ pbswd = 0.9
+ pbsws = 0.9
+ cigbacc = 0.245
+ tnoimod = 0
+ pdits = 0
+ cigsd = 0.013281
+ cigbinv = 0.006
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ ppdiblc2 = 0
+ tpbswg = 0.001
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ version = 4.5
+ tempmod = 0
+ tnoia = 0
+ peta0 = 2e-17
+ ptvoff = 0
+ aigbacc = 0.012071
+ tpbsw = 0.0025
+ pkvth0we = 0.0
+ pvfbsdoff = 0
+ keta = -0.042350111
+ cjswd = 4.743e-11
+ cjsws = 4.743e-11
+ diomod = 1
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ pditsd = 0
+ pditsl = 0
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ cjswgd = 1.6832999999999998e-10
+ pku0we = 0.0
+ cjswgs = 1.6832999999999998e-10
+ lcit = -2e-11
+ aigbinv = 0.009974
+ vfbsdoff = 0.01
+ wtvfbsdoff = 0
+ kt1l = 0
+ lint = 6.5375218e-9
+ ltvfbsdoff = 0
+ mjswgd = 0.95
+ mjswgs = 0.95
+ lkt1 = 6e-10
+ paramchk = 1
+ lmax = 2.001e-5
+ lmin = 9.00077e-6
+ tcjswg = 0.00128
+ scref = 1e-6
+ lpe0 = 6.44e-8
+ lpeb = 0
+ pigcd = 2.572
+ aigsd = 0.0063636
+ minv = -0.33
+ lvoff = 0
+ poxedge = 1
+ ndep = 1e+18
+ lwlc = 0
+ ijthdfwd = 0.01
+ lvsat = -0.00028
+ moin = 5.5538
+ lvth0 = 3e-10
+ binunit = 2
+ ptvfbsdoff = 0
+ nigc = 2.291
+ delta = 0.018814
+ rnoia = 0
+ rnoib = 0
+ fprout = 200
+ noff = 2.2684
+ ags = 0.8379228
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ ijthdrev = 0.01
+ ngate = 1.7e+20
+ cjd = 0.0012517799999999999
+ cit = 5e-6
+ cjs = 0.0012517799999999999
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 1.0572421799999999e-8
+ ngcon = 1
+ k3b = 2.1176
+ wpclm = 0
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ lpdiblc2 = 0
+ ntox = 2.958
+ wtvoff = 0
+ pcit = 1e-18
+ pclm = 1.484
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ la0 = 0
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = -0.0008
+ kt1 = -0.17107633
+ lk2 = -4e-10
+ kt2 = -0.04747
+ jtsswgd = 1.75e-7
+ phin = 0.15
+ llc = 0
+ jtsswgs = 1.75e-7
+ lln = 1
+ lu0 = -1.2e-11
+ mjd = 0.335
+ mjs = 0.335
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 0
+ capmod = 2
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ pk2 = 0
+ pkt1 = 5e-17
+ pu0 = 0
+ prt = 0
+ wku0we = 1.5e-11
+ pud = 0
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 1.1969344e-9
+ ub1 = -1.3666143e-18
+ uc1 = 6.873e-11
+ mobmod = 0
+ tpb = 0.0016
+ wa0 = 0
+ lkvth0we = 3e-12
+ ute = -1
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 0
+ wlc = 0
+ wln = 1
+ rbdb = 50
+ prwb = 0
+ wu0 = 0
+ prwg = 0
+ xgl = -8.2e-9
+ xgw = 0
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ rdsw = 200
+ tvoff = 0.0026155642
+ acnqsmod = 0
+ njtsswg = 6.489
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ xtsswgd = 0.32
+ rbodymod = 0
+ xtsswgs = 0.32
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.0026729629
+ ku0we = -0.0007
+ pdiblcb = 0
+ beta0 = 13.32
+ rshg = 14.1
+ leta0 = 6e-10
+ )

.model pch_ff_2 pmos (
+ level = 54
+ aigbinv = 0.009974
+ eta0 = 0.1672
+ tnoia = 0
+ etab = -0.23
+ ijthdfwd = 0.01
+ peta0 = 2e-17
+ toxref = 3e-9
+ pvfbsdoff = 0
+ tpbsw = 0.0025
+ cjswd = 4.743e-11
+ cjsws = 4.743e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ ijthdrev = 0.01
+ lpdiblc2 = 7.1311563e-9
+ poxedge = 1
+ ltvoff = -4.7585658e-10
+ binunit = 2
+ scref = 1e-6
+ pigcd = 2.572
+ aigsd = 0.0063636
+ lku0we = 1.8e-11
+ epsrox = 3.9
+ lkvth0we = 3e-12
+ lvoff = -8.0044387e-9
+ lvsat = -0.00028
+ rdsmod = 0
+ lvth0 = -4.8267694e-9
+ ags = 0.80385259
+ igbmod = 1
+ delta = 0.018814
+ laigc = -4.8397409e-11
+ cjd = 0.0012517799999999999
+ cit = 5e-6
+ cjs = 0.0012517799999999999
+ clc = 1e-7
+ cle = 0.6
+ acnqsmod = 0
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 1.0572421799999999e-8
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ k3b = 2.1176
+ rnoia = 0
+ rnoib = 0
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ keta = -0.040853613
+ pbswgd = 0.8
+ pbswgs = 0.8
+ rbodymod = 0
+ a0 = 2.5747309
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 72000
+ lags = 3.062912e-7
+ ngate = 1.7e+20
+ cf = 8.741900000000001e-11
+ igcmod = 1
+ la0 = -3.9314047e-7
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.0012551498
+ k3 = -2.5823
+ em = 20000000.0
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = -0.0008
+ ll = 0
+ lw = 0
+ kt1 = -0.16652617
+ kt2 = -0.046491549
+ lk2 = 3.9082075e-9
+ u0 = 0.0095048901
+ ngcon = 1
+ w0 = 0
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ ua = 1.4083134e-10
+ ub = 1.1675774e-18
+ uc = 1.8373185e-11
+ ud = 0
+ llc = 0
+ wpclm = 0
+ lln = 1
+ lcit = -2e-11
+ wl = 0
+ wr = 1
+ lu0 = -1.1012209880000001e-11
+ xj = 1.1e-7
+ xl = 2.33e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ mjd = 0.335
+ mjs = 0.335
+ lua = -1.0007073e-16
+ lub = 1.3480174e-25
+ luc = 1.5883665e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ kt1l = 0
+ njs = 1.02
+ pa0 = 0
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ pk2 = 0
+ gbmin = 1e-12
+ pu0 = 0
+ jswgd = 3.69e-13
+ prt = 0
+ jswgs = 3.69e-13
+ pud = 0
+ lint = 6.5375218e-9
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 1.1817684e-9
+ ub1 = -1.3634053e-18
+ uc1 = 6.7786161e-11
+ tpb = 0.0016
+ lkt1 = -4.0306013000000005e-8
+ lkt2 = -8.7962711e-9
+ wa0 = 0
+ lmax = 9.00077e-6
+ ute = -1
+ lmin = 9.0075e-7
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 0
+ wlc = 0
+ wln = 1
+ wu0 = 0
+ xgl = -8.2e-9
+ xgw = 0
+ njtsswg = 6.489
+ lpe0 = 6.44e-8
+ wud = 0
+ wpdiblc2 = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ lpeb = 0
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ minv = -0.33
+ lua1 = 1.3634229e-16
+ lub1 = -2.8849398e-26
+ luc1 = 8.4851172e-18
+ permod = 1
+ ckappad = 0.6
+ ckappas = 0.6
+ ndep = 1e+18
+ pdiblc1 = 0
+ pdiblc2 = 0.0018797309
+ pdiblcb = 0
+ lwlc = 0
+ moin = 5.5538
+ nigc = 2.291
+ tvoff = 0.002668496
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ wkvth0we = 0.0
+ voffcv = -0.125
+ wpemod = 1
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ bigbacc = 0.0054401
+ trnqsmod = 0
+ ku0we = -0.0007
+ beta0 = 13.32
+ kvth0we = -0.00022
+ ntox = 2.958
+ pcit = 1e-18
+ pclm = 1.484
+ leta0 = 6e-10
+ lintnoi = -5e-9
+ ppclm = 0
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ phin = 0.15
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ pkt1 = 5e-17
+ rgatemod = 0
+ tpbswg = 0.001
+ tnjtsswg = 1
+ tvfbsdoff = 0.1
+ dmcgt = 0
+ rbdb = 50
+ tcjsw = 9.34e-5
+ prwb = 0
+ prwg = 0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ ptvoff = 0
+ wtvfbsdoff = 0
+ rdsw = 200
+ bigsd = 0.0003327
+ diomod = 1
+ ltvfbsdoff = 0
+ pditsd = 0
+ pditsl = 0
+ nfactor = 1
+ wvoff = 0
+ cjswgd = 1.6832999999999998e-10
+ pku0we = 0.0
+ cjswgs = 1.6832999999999998e-10
+ wvfbsdoff = 0
+ wvsat = 0
+ lvfbsdoff = 0
+ wvth0 = 2.7e-9
+ rshg = 14.1
+ mjswgd = 0.95
+ mjswgs = 0.95
+ tcjswg = 0.00128
+ lketa = -1.3453518e-8
+ ptvfbsdoff = 0
+ nigbacc = 10
+ xpart = 1
+ tnom = 25
+ egidl = 0.001
+ toxe = 2.6300000000000002e-9
+ toxm = 2.67e-9
+ ijthsfwd = 0.01
+ nigbinv = 2.171
+ fprout = 200
+ xrcrg1 = 12
+ xrcrg2 = 1
+ ijthsrev = 0.01
+ fnoimod = 1
+ voff = -0.110213
+ wtvoff = 0
+ acde = 0.5
+ eigbinv = 1.1
+ pvoff = -2.5e-17
+ vsat = 120000
+ wint = 0
+ vth0 = -0.363565
+ cdscb = 0
+ cdscd = 0
+ wmax = 0.00090001
+ pvsat = 0
+ aigc = 0.0068361342
+ wmin = 8.9974e-6
+ wk2we = 0.0
+ capmod = 2
+ pvth0 = 1.5e-16
+ drout = 0.56
+ wku0we = 1.5e-11
+ ppdiblc2 = 0
+ mobmod = 0
+ voffl = 0
+ bigc = 0.0012521
+ weta0 = 2.8e-10
+ cigbacc = 0.245
+ wwlc = 0
+ lpclm = 0
+ cdsc = 0
+ tnoimod = 0
+ cgbo = 0
+ cgidl = 1
+ cgdl = 3.2212350000000004e-11
+ cgdo = 2.8335740000000002e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.2212350000000004e-11
+ cgso = 2.8335740000000002e-11
+ cigc = 0.15259
+ pkvth0we = 0.0
+ cigbinv = 0.006
+ pbswd = 0.9
+ pbsws = 0.9
+ vfbsdoff = 0.01
+ version = 4.5
+ tempmod = 0
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ pdits = 0
+ cigsd = 0.013281
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ dvt0w = 0
+ paramchk = 1
+ dvt1w = 0
+ dvt2w = 0
+ aigbacc = 0.012071
+ k2we = 5e-5
+ dsub = 0.5
+ dtox = 3.91e-10
+ pk2we = 0.0
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ )

.model pch_ff_3 pmos (
+ level = 54
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ nigbacc = 10
+ ijthsrev = 0.01
+ wvoff = 0
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ wvsat = 0
+ ntox = 2.958
+ wvth0 = 2.7e-9
+ pcit = 1e-18
+ pclm = 1.484
+ ltvoff = -2.3123852e-10
+ nigbinv = 2.171
+ phin = 0.15
+ lketa = -1.5940244e-8
+ pkt1 = 5e-17
+ ppdiblc2 = 0
+ xpart = 1
+ lku0we = 1.8e-11
+ epsrox = 3.9
+ egidl = 0.001
+ rbdb = 50
+ fnoimod = 1
+ prwb = 0
+ prwg = 0
+ rdsmod = 0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ eigbinv = 1.1
+ igbmod = 1
+ rdsw = 200
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ pbswgd = 0.8
+ pbswgs = 0.8
+ pkvth0we = 0.0
+ igcmod = 1
+ vfbsdoff = 0.01
+ rshg = 14.1
+ cigbacc = 0.245
+ pvoff = -2.5e-17
+ cdscb = 0
+ cdscd = 0
+ pvsat = 0
+ tnoimod = 0
+ wk2we = 0.0
+ pvth0 = 1.5e-16
+ paramchk = 1
+ drout = 0.56
+ cigbinv = 0.006
+ voffl = 0
+ permod = 1
+ tnom = 25
+ weta0 = 2.8e-10
+ toxe = 2.6300000000000002e-9
+ toxm = 2.67e-9
+ a0 = 2.8917556
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ lpclm = 0
+ at = 72000
+ cf = 8.741900000000001e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = 0.0040664684
+ k3 = -2.5823
+ em = 20000000.0
+ ijthdfwd = 0.01
+ version = 4.5
+ ll = 0
+ lw = 0
+ u0 = 0.009736756
+ w0 = 0
+ ua = 1.1413788e-10
+ ub = 1.1978347e-18
+ uc = 4.3035111e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 2.33e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ tempmod = 0
+ cgidl = 1
+ voffcv = -0.125
+ wpemod = 1
+ aigbacc = 0.012071
+ ijthdrev = 0.01
+ pbswd = 0.9
+ pbsws = 0.9
+ voff = -0.10886793
+ lpdiblc2 = 1.7469722e-9
+ acde = 0.5
+ vsat = 120000
+ aigbinv = 0.009974
+ wint = 0
+ vth0 = -0.36618963000000004
+ pdits = 0
+ cigsd = 0.013281
+ wmax = 0.00090001
+ aigc = 0.00683106
+ wmin = 8.9974e-6
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ wtvfbsdoff = 0
+ tpbswg = 0.001
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ ltvfbsdoff = 0
+ lkvth0we = 3e-12
+ bigc = 0.0012521
+ wwlc = 0
+ tnoia = 0
+ ptvoff = 0
+ poxedge = 1
+ cdsc = 0
+ peta0 = 2e-17
+ cgbo = 0
+ cgdl = 3.2212350000000004e-11
+ cgdo = 2.8335740000000002e-11
+ xtid = 3
+ xtis = 3
+ acnqsmod = 0
+ pvfbsdoff = 0
+ cgsl = 3.2212350000000004e-11
+ cgso = 2.8335740000000002e-11
+ cigc = 0.15259
+ binunit = 2
+ diomod = 1
+ tpbsw = 0.0025
+ cjswd = 4.743e-11
+ cjsws = 4.743e-11
+ mjswd = 0.01
+ pditsd = 0
+ mjsws = 0.01
+ pditsl = 0
+ rbodymod = 0
+ agidl = 3.2166e-9
+ cjswgd = 1.6832999999999998e-10
+ pku0we = 0.0
+ cjswgs = 1.6832999999999998e-10
+ ptvfbsdoff = 0
+ dmcg = 3.1e-8
+ mjswgd = 0.95
+ dmci = 3.1e-8
+ dmdg = 0
+ mjswgs = 0.95
+ tcjswg = 0.00128
+ k2we = 5e-5
+ jtsswgd = 1.75e-7
+ scref = 1e-6
+ jtsswgs = 1.75e-7
+ wpdiblc2 = 0
+ dsub = 0.5
+ pigcd = 2.572
+ dtox = 3.91e-10
+ aigsd = 0.0063635603
+ ags = 0.82774541
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ lvoff = -9.201547e-9
+ cjd = 0.0012517799999999999
+ cit = -8.7888889e-5
+ cjs = 0.0012517799999999999
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 1.0572421799999999e-8
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ eta0 = 0.1672
+ etab = -0.23
+ lvsat = -0.00028
+ lvth0 = -2.4908419000000002e-9
+ delta = 0.018814
+ laigc = -4.3881382e-11
+ la0 = -6.7529244e-7
+ fprout = 200
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = -0.0008
+ kt1 = -0.19559142
+ kt2 = -0.048919444
+ lk2 = -8.2803272e-10
+ llc = 0
+ lln = 1
+ lu0 = -2.1737244e-10
+ rnoia = 0
+ rnoib = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ mjd = 0.335
+ mjs = 0.335
+ lua = -7.6313554e-17
+ lub = 1.0787275e-25
+ luc = -6.0654489e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ wkvth0we = 0.0
+ njs = 1.02
+ pa0 = 0
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ pk2 = 0
+ njtsswg = 6.489
+ pu0 = 0
+ prt = 0
+ pud = 0
+ ngate = 1.7e+20
+ trnqsmod = 0
+ wtvoff = 0
+ ngcon = 1
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 1.2804108e-9
+ ub1 = -1.1625424e-18
+ uc1 = 4.6637333e-11
+ wpclm = 0
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ tpb = 0.0016
+ wa0 = 0
+ ute = -1
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 0
+ ckappad = 0.6
+ ckappas = 0.6
+ gbmin = 1e-12
+ wlc = 0
+ wln = 1
+ wu0 = 0
+ xgl = -8.2e-9
+ xgw = 0
+ pdiblc1 = 0
+ pdiblc2 = 0.0079293759
+ wud = 0
+ jswgd = 3.69e-13
+ wwc = 0
+ jswgs = 3.69e-13
+ wwl = 0
+ wwn = 1
+ pdiblcb = 0
+ capmod = 2
+ wku0we = 1.5e-11
+ rgatemod = 0
+ mobmod = 0
+ tnjtsswg = 1
+ bigbacc = 0.0054401
+ kvth0we = -0.00022
+ lintnoi = -5e-9
+ tvoff = 0.0023936443
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ laigsd = 3.5374533e-14
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ keta = -0.03805954
+ lags = 2.8502658e-7
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 6.2671111e-11
+ ku0we = -0.0007
+ beta0 = 13.32
+ kt1l = 0
+ leta0 = 6e-10
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ ppclm = 0
+ lint = 6.5375218e-9
+ lkt1 = -1.4437938999999999e-8
+ lkt2 = -6.6354444e-9
+ dlcig = 2.5e-9
+ lmax = 9.0075e-7
+ bgidl = 1834800000.0
+ lmin = 4.5075e-7
+ lpe0 = 6.44e-8
+ lpeb = 0
+ tvfbsdoff = 0.1
+ minv = -0.33
+ lua1 = 4.8550568e-17
+ nfactor = 1
+ lub1 = -2.0761736e-25
+ luc1 = 2.7307573e-17
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ ndep = 1e+18
+ lwlc = 0
+ ijthsfwd = 0.01
+ moin = 5.5538
+ nigc = 2.291
+ toxref = 3e-9
+ bigsd = 0.0003327
+ )

.model pch_ff_4 pmos (
+ level = 54
+ aigc = 0.0067884199
+ wmin = 8.9974e-6
+ cjd = 0.0012517799999999999
+ cit = -0.00054497817
+ cjs = 0.0012517799999999999
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 1.38228675e-8
+ scref = 1e-6
+ k3b = 2.1176
+ rgatemod = 0
+ lku0we = 1.8e-11
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ pigcd = 2.572
+ tnjtsswg = 1
+ epsrox = 3.9
+ aigsd = 0.0063636407
+ njtsswg = 6.489
+ lvoff = -3.8830249e-9
+ bigc = 0.0012521
+ la0 = -4.3379389e-8
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = -0.0008
+ rdsmod = 0
+ kt1 = -0.2000222
+ kt2 = -0.054670852
+ lk2 = 9.630220999999999e-10
+ wwlc = 0
+ llc = -1.18e-13
+ xtsswgd = 0.32
+ lln = 0.7
+ xtsswgs = 0.32
+ lu0 = -4.952545e-10
+ igbmod = 1
+ mjd = 0.335
+ mjs = 0.335
+ lua = -1.5477844e-16
+ lub = 5.0676856e-26
+ luc = -5.2541764e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ lvsat = -0.00028
+ njd = 1.02
+ njs = 1.02
+ pa0 = 0
+ lvth0 = 4.6404662e-9
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ ckappad = 0.6
+ pk2 = 0
+ ckappas = 0.6
+ cdsc = 0
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ pu0 = 0
+ pdiblc1 = 0
+ pdiblc2 = 0.013802718
+ delta = 0.018814
+ cgbo = 0
+ prt = 0
+ cgdl = 3.2212350000000004e-11
+ cgdo = 2.8335740000000002e-11
+ pud = 0
+ pdiblcb = 0
+ xtid = 3
+ xtis = 3
+ laigc = -2.5119727e-11
+ pbswgd = 0.8
+ pbswgs = 0.8
+ cgsl = 3.2212350000000004e-11
+ cgso = 2.8335740000000002e-11
+ rsh = 15.2
+ tcj = 0.000832
+ cigc = 0.15259
+ ua1 = 1.2553592e-9
+ ub1 = -1.2671808e-18
+ uc1 = 1.0455371e-10
+ rnoia = 0
+ rnoib = 0
+ tpb = 0.0016
+ wa0 = 0
+ igcmod = 1
+ ute = -1
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 0
+ wlc = 0
+ wln = 1
+ wu0 = 0
+ xgl = -8.2e-9
+ xgw = 0
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ ngate = 1.7e+20
+ ngcon = 1
+ wpclm = 0
+ bigbacc = 0.0054401
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ kvth0we = -0.00022
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ k2we = 5e-5
+ vtsswgs = 1.1
+ dsub = 0.5
+ dtox = 3.91e-10
+ permod = 1
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ eta0 = 0.1672
+ ijthsfwd = 0.01
+ etab = -0.23
+ tvoff = 0.002134918
+ voffcv = -0.125
+ wpemod = 1
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ ijthsrev = 0.01
+ wtvfbsdoff = 0
+ ku0we = -0.0007
+ beta0 = 13.32
+ nfactor = 1
+ leta0 = 6e-10
+ ltvfbsdoff = 0
+ ppclm = 0
+ a0 = 1.4555895
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 72000
+ cf = 8.741900000000001e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -4.1106394e-6
+ k3 = -2.5823
+ em = 20000000.0
+ ll = -1.18e-13
+ dlcig = 2.5e-9
+ lw = 0
+ u0 = 0.010368305999999999
+ w0 = 0
+ tpbswg = 0.001
+ ua = 2.9246716e-10
+ ub = 1.3278253e-18
+ uc = 4.119131e-11
+ ud = 0
+ bgidl = 1834800000.0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 2.33e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ ppdiblc2 = 0
+ tvfbsdoff = 0.1
+ nigbacc = 10
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ ptvoff = 0
+ ptvfbsdoff = 0
+ diomod = 1
+ nigbinv = 2.171
+ pkvth0we = 0.0
+ bigsd = 0.0003327
+ keta = -0.029364427
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.6832999999999998e-10
+ pku0we = 0.0
+ cjswgs = 1.6832999999999998e-10
+ wvoff = 0
+ lags = 5.4107004e-7
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 2.6379039e-10
+ vfbsdoff = 0.01
+ wvsat = 0
+ kt1l = 0
+ wvth0 = 2.7e-9
+ mjswgd = 0.95
+ mjswgs = 0.95
+ fnoimod = 1
+ eigbinv = 1.1
+ tcjswg = 0.00128
+ lint = 9.7879675e-9
+ lkt1 = -1.2488393e-8
+ lkt2 = -4.1048253e-9
+ paramchk = 1
+ lmax = 4.5075e-7
+ lmin = 2.1744e-7
+ lketa = -1.9766093e-8
+ lpe0 = 6.44e-8
+ xpart = 1
+ lpeb = 0
+ minv = -0.33
+ lua1 = 5.9573279e-17
+ lub1 = -1.6157647e-25
+ egidl = 0.001
+ luc1 = 1.8243668e-18
+ ndep = 1e+18
+ lwlc = 0
+ ijthdfwd = 0.01
+ moin = 5.5538
+ cigbacc = 0.245
+ fprout = 200
+ nigc = 2.291
+ xrcrg1 = 12
+ xrcrg2 = 1
+ tnoimod = 0
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ ijthdrev = 0.01
+ cigbinv = 0.006
+ wtvoff = 0
+ lpdiblc2 = -8.3729822e-10
+ ntox = 2.958
+ pcit = 1e-18
+ pclm = 1.484
+ pvoff = -2.5e-17
+ capmod = 2
+ version = 4.5
+ cdscb = 0
+ cdscd = 0
+ pvsat = 0
+ phin = 0.15
+ wku0we = 1.5e-11
+ tempmod = 0
+ wk2we = 0.0
+ pvth0 = 1.5e-16
+ drout = 0.56
+ mobmod = 0
+ pkt1 = 5e-17
+ voffl = 0
+ aigbacc = 0.012071
+ lkvth0we = 3e-12
+ weta0 = 2.8e-10
+ rbdb = 50
+ prwb = 0
+ prwg = 0
+ lpclm = 0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ rdsw = 200
+ aigbinv = 0.009974
+ cgidl = 1
+ acnqsmod = 0
+ rbodymod = 0
+ pbswd = 0.9
+ pbsws = 0.9
+ rshg = 14.1
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ pdits = 0
+ poxedge = 1
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ binunit = 2
+ wpdiblc2 = 0
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ tnom = 25
+ toxe = 2.6300000000000002e-9
+ toxm = 2.67e-9
+ tnoia = 0
+ toxref = 3e-9
+ peta0 = 2e-17
+ pvfbsdoff = 0
+ tpbsw = 0.0025
+ wkvth0we = 0.0
+ cjswd = 4.743e-11
+ cjsws = 4.743e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ trnqsmod = 0
+ voff = -0.12095548
+ acde = 0.5
+ ltvoff = -1.1739897e-10
+ vsat = 120000
+ wint = 0
+ vth0 = -0.38239713
+ wmax = 0.00090001
+ ags = 0.24582847
+ )

.model pch_ff_5 pmos (
+ level = 54
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ pbswgd = 0.8
+ pbswgs = 0.8
+ acnqsmod = 0
+ version = 4.5
+ tempmod = 0
+ igcmod = 1
+ keta = -0.12863898
+ rbodymod = 0
+ lags = 3.2185083e-8
+ aigbacc = 0.012071
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 5.594557300000001e-11
+ kt1l = 0
+ pvoff = -2.5e-17
+ cdscb = 0
+ cdscd = 0
+ lint = 9.7879675e-9
+ pvsat = 0.0
+ wk2we = 0.0
+ pvth0 = 1.5e-16
+ aigbinv = 0.009974
+ lkt1 = -4.140996599999999e-9
+ lkt2 = -5.2805906e-10
+ drout = 0.56
+ lmax = 2.1744e-7
+ lmin = 9.167e-8
+ wpdiblc2 = 0
+ lpe0 = 6.44e-8
+ permod = 1
+ lpeb = 0
+ voffl = 0
+ minv = -0.33
+ lua1 = -1.5051887e-16
+ lub1 = 1.742578e-25
+ luc1 = 7.2216103e-18
+ weta0 = 2.8e-10
+ ndep = 1e+18
+ lpclm = -1.4239795e-8
+ wtvfbsdoff = 0
+ lwlc = 0
+ moin = 5.5538
+ cgidl = 1
+ voffcv = -0.125
+ wpemod = 1
+ nigc = 2.291
+ ltvfbsdoff = 0
+ poxedge = 1
+ wkvth0we = 0.0
+ noff = 2.2684
+ binunit = 2
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ pbswd = 0.9
+ pbsws = 0.9
+ trnqsmod = 0
+ ntox = 2.958
+ pcit = 1e-18
+ pclm = 1.5514872
+ pdits = 0
+ cigsd = 0.013281
+ phin = 0.15
+ tpbswg = 0.001
+ ptvfbsdoff = 0
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ pkt1 = 5e-17
+ rgatemod = 0
+ tnjtsswg = 1
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ ptvoff = 0
+ rbdb = 50
+ prwb = 0
+ prwg = 0
+ tnoia = 0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ pvfbsdoff = 0
+ rdsw = 200
+ peta0 = 2e-17
+ diomod = 1
+ tpbsw = 0.0025
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.6832999999999998e-10
+ pku0we = 0.0
+ cjswgs = 1.6832999999999998e-10
+ cjswd = 4.743e-11
+ a0 = 1.4508547
+ a1 = 0
+ a2 = 1
+ cjsws = 4.743e-11
+ b0 = 0
+ b1 = 0
+ mjswd = 0.01
+ at = 72000
+ cf = 8.741900000000001e-11
+ mjsws = 0.01
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.013949949
+ k3 = -2.5823
+ agidl = 3.2166e-9
+ em = 20000000.0
+ ll = -1.18e-13
+ lw = 0
+ u0 = 0.0089521197
+ w0 = 0
+ ua = -3.1871506e-10
+ ub = 1.6925299e-18
+ uc = 2.1642376e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 2.33e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ ags = 2.6576055
+ njtsswg = 6.489
+ mjswgd = 0.95
+ mjswgs = 0.95
+ cjd = 0.0012517799999999999
+ cit = 0.00044006838
+ cjs = 0.0012517799999999999
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ rshg = 14.1
+ bvs = 8.2
+ dlc = 1.38228675e-8
+ xtsswgd = 0.32
+ k3b = 2.1176
+ xtsswgs = 0.32
+ tcjswg = 0.00128
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.016932267
+ pdiblcb = 0
+ la0 = -4.2380342e-8
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = -0.0008
+ kt1 = -0.23958332
+ kt2 = -0.07162235
+ lk2 = 3.9055939e-9
+ scref = 1e-6
+ llc = -1.18e-13
+ lln = 0.7
+ lu0 = -1.9643925000000002e-10
+ mjd = 0.335
+ mjs = 0.335
+ lua = -2.581899e-17
+ lub = -2.6275812e-26
+ luc = -1.1293514e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ pigcd = 2.572
+ njd = 1.02
+ njs = 1.02
+ aigsd = 0.0063636407
+ pa0 = 0
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ pk2 = 0
+ pu0 = 0
+ prt = 0
+ pud = 0
+ tnom = 25
+ lvoff = -1.3382853e-9
+ rsh = 15.2
+ toxe = 2.6300000000000002e-9
+ toxm = 2.67e-9
+ tcj = 0.000832
+ ua1 = 2.2510566e-9
+ ub1 = -2.8588123e-18
+ uc1 = 7.8974359e-11
+ bigbacc = 0.0054401
+ tpb = 0.0016
+ lvsat = -0.0004495331599999999
+ ijthsfwd = 0.01
+ wa0 = 0
+ ute = -1
+ lvth0 = 4.9692121999999995e-9
+ web = 6628.3
+ wec = -16935.0
+ fprout = 200
+ wk2 = 0
+ wlc = 0
+ wln = 1
+ wu0 = 0
+ xgl = -8.2e-9
+ xgw = 0
+ delta = 0.018814
+ wud = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ laigc = -2.0986759e-11
+ kvth0we = -0.00022
+ rnoia = 0
+ rnoib = 0
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ wtvoff = 0
+ vtsswgs = 1.1
+ ijthsrev = 0.01
+ ngate = 1.7e+20
+ wcit = 0.0
+ ngcon = 1
+ wpclm = 0
+ voff = -0.13301586
+ acde = 0.5
+ gbmin = 1e-12
+ capmod = 2
+ vsat = 120803.55
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ wint = 0
+ vth0 = -0.38395511000000004
+ wku0we = 1.5e-11
+ wmax = 0.00090001
+ aigc = 0.0067688324
+ wmin = 8.9974e-6
+ mobmod = 0
+ ppdiblc2 = 0
+ bigc = 0.0012521
+ wwlc = 0
+ nfactor = 1
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.2212350000000004e-11
+ cgdo = 2.8335740000000002e-11
+ xtid = 3
+ xtis = 3
+ tvoff = 0.0018930751
+ cgsl = 3.2212350000000004e-11
+ cgso = 2.8335740000000002e-11
+ cigc = 0.15259
+ xjbvd = 1
+ xjbvs = 1
+ pkvth0we = 0.0
+ lk2we = 0.0
+ vfbsdoff = 0.01
+ ku0we = -0.0007
+ nigbacc = 10
+ beta0 = 13.32
+ leta0 = 6e-10
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ ppclm = 0
+ paramchk = 1
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ nigbinv = 2.171
+ k2we = 5e-5
+ tvfbsdoff = 0.1
+ dsub = 0.5
+ dtox = 3.91e-10
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ eta0 = 0.1672
+ ijthdfwd = 0.01
+ etab = -0.23
+ toxref = 3e-9
+ fnoimod = 1
+ eigbinv = 1.1
+ bigsd = 0.0003327
+ ijthdrev = 0.01
+ wvfbsdoff = 0
+ wvoff = 0
+ lvfbsdoff = 0
+ ltvoff = -6.6370123e-11
+ lpdiblc2 = -1.4976331e-9
+ wvsat = 0.0
+ wvth0 = 2.7e-9
+ cigbacc = 0.245
+ lku0we = 1.8e-11
+ lketa = 1.1808374e-9
+ tnoimod = 0
+ epsrox = 3.9
+ xpart = 1
+ rdsmod = 0
+ cigbinv = 0.006
+ egidl = 0.001
+ lkvth0we = 3e-12
+ igbmod = 1
+ )

.model pch_ff_6 pmos (
+ level = 54
+ wpclm = 0
+ vfbsdoff = 0.01
+ rshg = 14.1
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ nfactor = 1
+ wtvfbsdoff = 0
+ paramchk = 1
+ permod = 1
+ ltvfbsdoff = 0
+ tnom = 25
+ toxe = 2.6300000000000002e-9
+ toxm = 2.67e-9
+ nigbacc = 10
+ ijthdfwd = 0.01
+ voffcv = -0.125
+ wpemod = 1
+ tvoff = 0.00091084129
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ nigbinv = 2.171
+ ptvfbsdoff = 0
+ ijthdrev = 0.01
+ wcit = 0.0
+ ku0we = -0.0007
+ lpdiblc2 = 0
+ voff = -0.11896044
+ beta0 = 13.32
+ acde = 0.5
+ leta0 = -5.141465e-10
+ letab = 2.0255694e-8
+ vsat = 166989.83000000002
+ wint = 0
+ vth0 = -0.32252512000000005
+ ppclm = 0
+ tpbswg = 0.001
+ wmax = 0.00090001
+ fnoimod = 1
+ aigc = 0.0067067782
+ wmin = 8.9974e-6
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ eigbinv = 1.1
+ tvfbsdoff = 0.1
+ ptvoff = 0
+ lkvth0we = 3e-12
+ bigc = 0.0012521
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ wwlc = 0
+ diomod = 1
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.2212350000000004e-11
+ cgdo = 2.8335740000000002e-11
+ xtid = 3
+ xtis = 3
+ acnqsmod = 0
+ pditsd = 0
+ pditsl = 0
+ cgsl = 3.2212350000000004e-11
+ cjswgd = 1.6832999999999998e-10
+ pku0we = 0.0
+ cgso = 2.8335740000000002e-11
+ cigbacc = 0.245
+ cjswgs = 1.6832999999999998e-10
+ cigc = 0.15259
+ bigsd = 0.0003327
+ rbodymod = 0
+ wvfbsdoff = 0
+ tnoimod = 0
+ lvfbsdoff = 0
+ wvoff = 0
+ mjswgd = 0.95
+ mjswgs = 0.95
+ wvsat = 0.0
+ cigbinv = 0.006
+ wvth0 = 2.7e-9
+ tcjswg = 0.00128
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ version = 4.5
+ lketa = 8.4925319e-9
+ k2we = 5e-5
+ tempmod = 0
+ wpdiblc2 = 0
+ xpart = 1
+ dsub = 0.5
+ dtox = 3.91e-10
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ egidl = 0.001
+ a0 = 3.4166667
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 140456.11
+ cf = 8.741900000000001e-11
+ aigbacc = 0.012071
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.010241786
+ k3 = -2.5823
+ em = 20000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.0049438888999999995
+ w0 = 0
+ ua = -1.1682959e-9
+ ub = 1.2873333e-18
+ uc = -8.7638e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 2.33e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ fprout = 200
+ eta0 = 0.17905262
+ etab = -0.44548611
+ xrcrg1 = 12
+ xrcrg2 = 1
+ aigbinv = 0.009974
+ wkvth0we = 0.0
+ wtvoff = 0
+ trnqsmod = 0
+ capmod = 2
+ pvoff = -2.5e-17
+ wku0we = 1.5e-11
+ cdscb = 0
+ cdscd = 0
+ mobmod = 0
+ pvsat = 0.0
+ wk2we = 0.0
+ pvth0 = 1.5e-16
+ drout = 0.56
+ poxedge = 1
+ rgatemod = 0
+ voffl = 0
+ tnjtsswg = 1
+ binunit = 2
+ weta0 = 2.8e-10
+ lpclm = -9.8438889e-8
+ cgidl = 1
+ keta = -0.20642296
+ pbswd = 0.9
+ pbsws = 0.9
+ lags = -2.8753242e-8
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ lcit = 8.979724e-11
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ kt1l = 0
+ pdits = 0
+ cigsd = 0.013281
+ lint = 0
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ lkt1 = -6.3119e-10
+ lkt2 = 1.5220167e-10
+ lmax = 9.167e-8
+ lmin = 5.567e-8
+ lpe0 = 6.44e-8
+ lpeb = 0
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ minv = -0.33
+ lua1 = -7.3062676e-18
+ lub1 = 1.0038041e-26
+ luc1 = 7.6176556e-18
+ ndep = 1e+18
+ toxref = 3e-9
+ njtsswg = 6.489
+ tnoia = 0
+ ijthsfwd = 0.01
+ lwlc = 0
+ pvfbsdoff = 0
+ moin = 5.5538
+ xtsswgd = 0.32
+ peta0 = 2e-17
+ xtsswgs = 0.32
+ nigc = 2.291
+ ckappad = 0.6
+ ckappas = 0.6
+ tpbsw = 0.0025
+ ags = 3.3058856
+ pdiblc1 = 0
+ pdiblc2 = 0.001
+ pdiblcb = 0
+ cjswd = 4.743e-11
+ cjd = 0.0012517799999999999
+ cjsws = 4.743e-11
+ cit = 7.994489e-5
+ cjs = 0.0012517799999999999
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ dlc = 4.0349e-9
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ k3b = 2.1176
+ ijthsrev = 0.01
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ ltvoff = 2.5959859e-11
+ la0 = -2.2716667e-7
+ ntox = 2.958
+ pcit = 1e-18
+ jsd = 1.5e-7
+ pclm = 2.4472222
+ jss = 1.5e-7
+ lat = -0.007234874400000001
+ kt1 = -0.27692169
+ kt2 = -0.078859167
+ lk2 = 3.5570266e-9
+ llc = 0
+ lln = 1
+ lu0 = 1.8033444e-10
+ mjd = 0.335
+ bigbacc = 0.0054401
+ mjs = 0.335
+ lua = 5.4041604e-17
+ lub = 1.1812662e-26
+ luc = 9.143004e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 0
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ pk2 = 0
+ phin = 0.15
+ pu0 = 0
+ lku0we = 1.8e-11
+ prt = 0
+ pub = 0.0
+ pud = 0
+ kvth0we = -0.00022
+ epsrox = 3.9
+ ppdiblc2 = 0
+ rsh = 15.2
+ scref = 1e-6
+ pkt1 = 5e-17
+ tcj = 0.000832
+ ua1 = 7.2751825e-10
+ ub1 = -1.1117937e-18
+ uc1 = 7.4761111e-11
+ tpb = 0.0016
+ pigcd = 2.572
+ lintnoi = -5e-9
+ wa0 = 0
+ aigsd = 0.0063636407
+ ute = -1
+ web = 6628.3
+ wec = -16935.0
+ bigbinv = 0.00149
+ wk2 = 0
+ rdsmod = 0
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ wlc = 0
+ wln = 1
+ wu0 = 0
+ xgl = -8.2e-9
+ xgw = 0
+ wub = 0.0
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ igbmod = 1
+ lvoff = -2.6594942e-9
+ rbdb = 50
+ prwb = 0
+ prwg = 0
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ rbpb = 50
+ rbpd = 50
+ lvsat = -0.0047910409
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ lvth0 = -8.05207e-10
+ pbswgd = 0.8
+ pbswgs = 0.8
+ rdsw = 200
+ delta = 0.018814
+ laigc = -1.5153664e-11
+ igcmod = 1
+ rnoia = 0
+ rnoib = 0
+ pkvth0we = 0.0
+ ngate = 1.7e+20
+ ngcon = 1
+ )

.model pch_ff_7 pmos (
+ level = 54
+ voffl = 0
+ dsub = 0.5
+ dtox = 3.91e-10
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ weta0 = 2.8e-10
+ ptvfbsdoff = 0
+ lpclm = -4.4240467e-8
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ eta0 = 0.18948293
+ ijthsfwd = 0.01
+ voffcv = -0.125
+ wpemod = 1
+ etab = -0.27185615
+ cgidl = 1
+ ijthsrev = 0.01
+ pbswd = 0.9
+ pbsws = 0.9
+ njtsswg = 6.489
+ tpbswg = 0.001
+ pdits = 0
+ cigsd = 0.013281
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ ppdiblc2 = 0
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.001
+ pdiblcb = 0
+ pk2we = 0.0
+ ptvoff = 0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ ags = 2.81014
+ pvfbsdoff = 0
+ tnoia = 0
+ diomod = 1
+ cjd = 0.0012517799999999999
+ cit = 0.0018532278000000005
+ cjs = 0.0012517799999999999
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 4.0349e-9
+ peta0 = 2e-17
+ k3b = 2.1176
+ pditsd = 0
+ pditsl = 0
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ bigbacc = 0.0054401
+ dwj = 0
+ cjswgd = 1.6832999999999998e-10
+ pku0we = 0.0
+ cjswgs = 1.6832999999999998e-10
+ tpbsw = 0.0025
+ pkvth0we = 0.0
+ keta = 0.048888889
+ cjswd = 4.743e-11
+ kvth0we = -0.00022
+ cjsws = 4.743e-11
+ la0 = -1.5788889e-7
+ jsd = 1.5e-7
+ mjswd = 0.01
+ jss = 1.5e-7
+ lat = 0.0034661578
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ kt1 = -0.090229195
+ kt2 = -0.087042222
+ lk2 = 3.9353879e-9
+ llc = 0
+ lln = 1
+ lu0 = -8.4628889e-11
+ mjd = 0.335
+ mjs = 0.335
+ lua = -4.5270917e-17
+ lub = -2.9222082e-26
+ luc = -2.161341e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ lintnoi = -5e-9
+ njd = 1.02
+ mjswgd = 0.95
+ njs = 1.02
+ mjswgs = 0.95
+ pa0 = 0
+ bigbinv = 0.00149
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ jswd = 3.69e-13
+ vtsswgd = 1.1
+ pk2 = 0
+ jsws = 3.69e-13
+ vtsswgs = 1.1
+ vfbsdoff = 0.01
+ lcit = -1.305310999999997e-11
+ pu0 = 0
+ tcjswg = 0.00128
+ prt = 0
+ pub = 0.0
+ pud = 0
+ kt1l = 0
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 1.0031266e-9
+ ub1 = -2.5489021e-18
+ uc1 = 1.9738889e-10
+ tpb = 0.0016
+ wa0 = 0
+ ute = -1
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 0
+ lint = 0
+ wlc = 0
+ wln = 1
+ wu0 = 0
+ xgl = -8.2e-9
+ xgw = 0
+ paramchk = 1
+ wub = 0.0
+ wud = 0
+ wwc = 0
+ lkt1 = -1.1459355e-8
+ lkt2 = 6.2681889e-10
+ wwl = 0
+ wwn = 1
+ lmax = 5.567e-8
+ lmin = 4.667e-8
+ scref = 1e-6
+ lpe0 = 6.44e-8
+ lpeb = 0
+ pigcd = 2.572
+ aigsd = 0.0063636407
+ minv = -0.33
+ lvoff = -4.1866651e-9
+ lua1 = -2.3291554e-17
+ lub1 = 9.339033e-26
+ luc1 = 5.0524444e-19
+ fprout = 200
+ ndep = 1e+18
+ lvsat = -0.0019989942799999998
+ ijthdfwd = 0.01
+ xrcrg1 = 12
+ xrcrg2 = 1
+ lwlc = 0
+ lvth0 = -1.7008558999999998e-9
+ moin = 5.5538
+ delta = 0.018814
+ laigc = -9.9932362e-12
+ nigc = 2.291
+ nfactor = 1
+ rnoia = 0
+ rnoib = 0
+ wtvoff = 0
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ ijthdrev = 0.01
+ ngate = 1.7e+20
+ ngcon = 1
+ wpclm = 0
+ lpdiblc2 = 0
+ capmod = 2
+ ntox = 2.958
+ pcit = 1e-18
+ wku0we = 1.5e-11
+ pclm = 1.5127667
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ nigbacc = 10
+ a0 = 2.2222222
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = -44044.444
+ mobmod = 0
+ cf = 8.741900000000001e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.016765256
+ k3 = -2.5823
+ em = 20000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.0095122222
+ w0 = 0
+ ua = 5.4398899e-10
+ ub = 1.9948286e-18
+ uc = 4.42645e-10
+ ud = 0
+ phin = 0.15
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 2.33e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ pkt1 = 5e-17
+ nigbinv = 2.171
+ lkvth0we = 3e-12
+ rbdb = 50
+ prwb = 0
+ prwg = 0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ rdsw = 200
+ tvoff = 0.0051729841
+ acnqsmod = 0
+ fnoimod = 1
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ eigbinv = 1.1
+ rbodymod = 0
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = -1.1191043e-9
+ rshg = 14.1
+ letab = 1.0185157e-8
+ ppclm = 0
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ tvfbsdoff = 0.1
+ cigbacc = 0.245
+ wpdiblc2 = 0
+ tnoimod = 0
+ tnom = 25
+ dmcgt = 0
+ toxref = 3e-9
+ tcjsw = 9.34e-5
+ toxe = 2.6300000000000002e-9
+ toxm = 2.67e-9
+ cigbinv = 0.006
+ bigsd = 0.0003327
+ wkvth0we = 0.0
+ version = 4.5
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ tempmod = 0
+ ltvoff = -2.2124443e-10
+ wvoff = 0
+ wcit = 0.0
+ trnqsmod = 0
+ voff = -0.092629909
+ wvsat = 0.0
+ acde = 0.5
+ wvth0 = 2.7e-9
+ aigbacc = 0.012071
+ vsat = 118851.091
+ wint = 0
+ vth0 = -0.30708289
+ lku0we = 1.8e-11
+ wmax = 0.00090001
+ aigc = 0.0066178053
+ wmin = 8.9974e-6
+ epsrox = 3.9
+ lketa = -6.3155556e-9
+ rgatemod = 0
+ xpart = 1
+ aigbinv = 0.009974
+ tnjtsswg = 1
+ rdsmod = 0
+ igbmod = 1
+ egidl = 0.001
+ bigc = 0.0012521
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ wwlc = 0
+ pbswgd = 0.8
+ pbswgs = 0.8
+ cdsc = 0
+ cgbo = 0
+ igcmod = 1
+ cgdl = 3.2212350000000004e-11
+ cgdo = 2.8335740000000002e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.2212350000000004e-11
+ cgso = 2.8335740000000002e-11
+ cigc = 0.15259
+ wtvfbsdoff = 0
+ poxedge = 1
+ binunit = 2
+ ltvfbsdoff = 0
+ pvoff = -2.5e-17
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ cdscb = 0
+ cdscd = 0
+ pvsat = 0.0
+ wk2we = 0.0
+ pvth0 = 1.5e-16
+ drout = 0.56
+ permod = 1
+ k2we = 5e-5
+ )

.model pch_ff_8 pmos (
+ level = 54
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ wkvth0we = 0.0
+ cigbacc = 0.245
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ trnqsmod = 0
+ ku0we = -0.0007
+ tnoimod = 0
+ beta0 = 13.32
+ leta0 = 2.7323128e-9
+ ntox = 2.958
+ letab = 3.9337702e-9
+ pcit = 1e-18
+ pclm = 1.0208333
+ tpbswg = 0.001
+ cigbinv = 0.006
+ ppclm = 0
+ phin = 0.15
+ dlcig = 2.5e-9
+ tvfbsdoff = 0.1
+ bgidl = 1834800000.0
+ pkt1 = 5e-17
+ rgatemod = 0
+ ptvoff = 0
+ tnjtsswg = 1
+ version = 4.5
+ tempmod = 0
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ diomod = 1
+ rbdb = 50
+ prwb = 0
+ prwg = 0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ aigbacc = 0.012071
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.6832999999999998e-10
+ pku0we = 0.0
+ cjswgs = 1.6832999999999998e-10
+ rdsw = 200
+ bigsd = 0.0003327
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ mjswgd = 0.95
+ mjswgs = 0.95
+ wvoff = 0
+ aigbinv = 0.009974
+ tcjswg = 0.00128
+ wvsat = 0.0
+ wvth0 = 2.7e-9
+ rshg = 14.1
+ lketa = 8.0381778e-9
+ xpart = 1
+ poxedge = 1
+ egidl = 0.001
+ tnom = 25
+ fprout = 200
+ toxe = 2.6300000000000002e-9
+ toxm = 2.67e-9
+ xrcrg1 = 12
+ xrcrg2 = 1
+ binunit = 2
+ ijthsfwd = 0.01
+ wtvoff = 0
+ ijthsrev = 0.01
+ wcit = 0.0
+ capmod = 2
+ voff = -0.10032114
+ wku0we = 1.5e-11
+ acde = 0.5
+ pvoff = -2.5e-17
+ mobmod = 0
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ vsat = 101742.52
+ wint = 0
+ vth0 = -0.35182997000000005
+ cdscb = 0
+ cdscd = 0
+ wkt1 = 0.0
+ pvsat = 0.0
+ wmax = 0.00090001
+ wk2we = 0.0
+ pvth0 = 1.5e-16
+ aigc = 0.0065563017
+ wmin = 8.9974e-6
+ drout = 0.56
+ ppdiblc2 = 0
+ voffl = 0
+ weta0 = 2.8e-10
+ wetab = 0
+ bigc = 0.0012521
+ wwlc = 0
+ lpclm = -2.0135733e-8
+ laigsd = -2.1777787e-18
+ cdsc = 0
+ cgidl = 1
+ njtsswg = 6.489
+ cgbo = 0
+ cgdl = 3.2212350000000004e-11
+ cgdo = 2.8335740000000002e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.2212350000000004e-11
+ cgso = 2.8335740000000002e-11
+ cigc = 0.15259
+ a0 = -0.19555556
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ xtsswgd = 0.32
+ pkvth0we = 0.0
+ xtsswgs = 0.32
+ at = 45108.9
+ cf = 8.741900000000001e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.012217534
+ k3 = -2.5823
+ em = 20000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.0050077778
+ w0 = 0
+ ua = -1.1794951e-9
+ ub = 1.3471713999999999e-18
+ uc = 5.0701667e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 2.33e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.001
+ pbswd = 0.9
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ pbsws = 0.9
+ pdiblcb = 0
+ vfbsdoff = 0.01
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ pdits = 0
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ paramchk = 1
+ bigbacc = 0.0054401
+ k2we = 5e-5
+ ags = 1.0774289
+ dsub = 0.5
+ kvth0we = -0.00022
+ dtox = 3.91e-10
+ cjd = 0.0012517799999999999
+ cit = -0.00424944667
+ pk2we = 0.0
+ cjs = 0.0012517799999999999
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ dlc = 4.0349e-9
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ k3b = 2.1176
+ toxref = 3e-9
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ pvfbsdoff = 0
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ tnoia = 0
+ ijthdfwd = 0.01
+ eta0 = 0.11088258
+ etab = -0.14427684
+ la0 = -3.9417778e-8
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = -0.0009023600000000003
+ kt1 = -0.32613297
+ kt2 = -0.08425
+ lk2 = 3.7125495e-9
+ peta0 = 2e-17
+ llc = 0
+ lln = 1
+ lu0 = 1.3608888999999998e-10
+ petab = 0
+ mjd = 0.335
+ mjs = 0.335
+ lua = 3.9179804e-17
+ lub = 2.5131622e-27
+ luc = -2.4081867e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 0
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0.0
+ pbs = 0.75
+ tpbsw = 0.0025
+ pk2 = 0
+ pu0 = 0
+ prt = 0
+ pub = 0.0
+ pud = 0
+ cjswd = 4.743e-11
+ cjsws = 4.743e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ ltvoff = -2.4936809e-11
+ agidl = 3.2166e-9
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 1.4917512e-9
+ ub1 = -1.5908843e-18
+ uc1 = 1.6325556e-10
+ ijthdrev = 0.01
+ tpb = 0.0016
+ wa0 = 0
+ ute = -1
+ wat = 0.0
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 0
+ wlc = 0
+ wln = 1
+ lpdiblc2 = 0
+ wu0 = 0
+ xgl = -8.2e-9
+ xgw = 0
+ wub = 0.0
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ lku0we = 1.8e-11
+ epsrox = 3.9
+ nfactor = 1
+ scref = 1e-6
+ rdsmod = 0
+ pigcd = 2.572
+ aigsd = 0.0063636407
+ igbmod = 1
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ wtvfbsdoff = 0
+ lvoff = -3.8097951e-9
+ lkvth0we = 3e-12
+ pbswgd = 0.8
+ pbswgs = 0.8
+ lvsat = -0.0011606774000000003
+ lvth0 = 4.91746942e-10
+ igcmod = 1
+ ltvfbsdoff = 0
+ delta = 0.018814
+ nigbacc = 10
+ laigc = -6.97956e-12
+ acnqsmod = 0
+ rnoia = 0
+ rnoib = 0
+ keta = -0.24404444
+ rbodymod = 0
+ ngate = 1.7e+20
+ lags = 8.4902844e-8
+ ngcon = 1
+ nigbinv = 2.171
+ wpclm = 0
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 2.8597836999999995e-10
+ kt1l = 0
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ ptvfbsdoff = 0
+ lint = 0
+ permod = 1
+ lkt1 = 9.993259999999988e-11
+ lkt2 = 4.9e-10
+ lmax = 4.667e-8
+ lmin = 3.6e-8
+ fnoimod = 1
+ wpdiblc2 = 0
+ lpe0 = 6.44e-8
+ lpeb = 0
+ eigbinv = 1.1
+ minv = -0.33
+ lua1 = -4.7234158e-17
+ lub1 = 4.6447457e-26
+ luc1 = 2.1777778e-18
+ voffcv = -0.125
+ wpemod = 1
+ ndep = 1e+18
+ lwlc = 0
+ moin = 5.5538
+ tvoff = 0.0011667062
+ nigc = 2.291
+ )

.model pch_ff_9 pmos (
+ level = 54
+ vtsswgs = 1.1
+ ags = 0.82538676
+ vsat = 121084.96
+ wint = 0
+ vth0 = -0.36548403
+ pdits = 0
+ cjd = 0.0012517799999999999
+ cit = 5e-6
+ cjs = 0.0012517799999999999
+ clc = 1e-7
+ cle = 0.6
+ cigsd = 0.013281
+ bvd = 8.2
+ bvs = 8.2
+ wkt1 = -1.0361455e-8
+ wkt2 = -3.8769913e-9
+ dlc = 1.0572421799999999e-8
+ wmax = 8.9974e-6
+ dvt0w = 0
+ k3b = 2.1176
+ dvt1w = 0
+ aigc = 0.0068303602
+ dvt2w = 0
+ wmin = 8.974e-7
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ ptvoff = 0
+ waigsd = 1.9139418e-12
+ la0 = 0
+ pk2we = 0.0
+ jsd = 1.5e-7
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ jss = 1.5e-7
+ lat = -0.0008
+ wua1 = -3.2799159e-16
+ kt1 = -0.16992583
+ lk2 = -4e-10
+ kt2 = -0.04703951
+ wub1 = 5.9231251e-25
+ wuc1 = -8.7396626e-17
+ llc = 0
+ lln = 1
+ lu0 = -1.2e-11
+ mjd = 0.335
+ mjs = 0.335
+ lkvth0we = 3e-12
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ diomod = 1
+ pvfbsdoff = 0
+ njd = 1.02
+ bigc = 0.0012521
+ njs = 1.02
+ wute = -7.8572347e-8
+ pa0 = 0
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ wwlc = 0
+ pk2 = 0
+ tnoia = 0
+ pu0 = 0
+ pditsd = 0
+ pditsl = 0
+ prt = 0
+ pud = 0
+ cjswgd = 1.6832999999999998e-10
+ pku0we = 0.0
+ cjswgs = 1.6832999999999998e-10
+ rsh = 15.2
+ tcj = 0.000832
+ peta0 = 2e-17
+ cdsc = 0
+ ua1 = 1.2333536e-9
+ ub1 = -1.432383e-18
+ uc1 = 7.8434267e-11
+ cgbo = 0
+ tpb = 0.0016
+ cgdl = 3.2212350000000004e-11
+ cgdo = 2.8335740000000002e-11
+ acnqsmod = 0
+ xtid = 3
+ xtis = 3
+ wketa = 2.2362589e-8
+ wa0 = 3.3745816e-7
+ ute = -0.99127556
+ web = 6628.3
+ wec = -16935.0
+ cgsl = 3.2212350000000004e-11
+ cgso = 2.8335740000000002e-11
+ wk2 = -2.287053e-9
+ tpbsw = 0.0025
+ cigc = 0.15259
+ wlc = 0
+ wln = 1
+ wu0 = -8.6631049e-11
+ xgl = -8.2e-9
+ xgw = 0
+ wua = -1.124189e-16
+ wub = -6.7100784e-26
+ wuc = -2.319496e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ cjswd = 4.743e-11
+ nfactor = 1
+ cjsws = 4.743e-11
+ mjswd = 0.01
+ mjswgd = 0.95
+ mjsws = 0.01
+ mjswgs = 0.95
+ agidl = 3.2166e-9
+ rbodymod = 0
+ tcjswg = 0.00128
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ nigbacc = 10
+ scref = 1e-6
+ k2we = 5e-5
+ wpdiblc2 = 3.6469361e-10
+ pigcd = 2.572
+ dsub = 0.5
+ aigsd = 0.0063633875
+ dtox = 3.91e-10
+ fprout = 200
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ lvoff = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ nigbinv = 2.171
+ lvsat = -0.00028
+ eta0 = 0.16744607
+ etab = -0.23671111
+ lvth0 = 3e-10
+ delta = 0.018814
+ wtvoff = -9.8925647e-11
+ rnoia = 0
+ rnoib = 0
+ wkvth0we = 0.0
+ fnoimod = 1
+ ngate = 1.7e+20
+ capmod = 2
+ trnqsmod = 0
+ eigbinv = 1.1
+ ngcon = 1
+ wpclm = -3.01194e-7
+ wku0we = 1.5e-11
+ mobmod = 0
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ rgatemod = 0
+ tnjtsswg = 1
+ cigbacc = 0.245
+ tnoimod = 0
+ tvoff = 0.0026265487
+ cigbinv = 0.006
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ keta = -0.044833188
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ version = 4.5
+ jswd = 3.69e-13
+ ku0we = -0.0007
+ jsws = 3.69e-13
+ lcit = -2e-11
+ tempmod = 0
+ beta0 = 13.32
+ leta0 = 6e-10
+ kt1l = 0
+ ppclm = 0
+ aigbacc = 0.012071
+ lint = 6.5375218e-9
+ tvfbsdoff = 0.1
+ dlcig = 2.5e-9
+ lkt1 = 6e-10
+ bgidl = 1834800000.0
+ lmax = 2.001e-5
+ lmin = 9.00077e-6
+ lpe0 = 6.44e-8
+ lpeb = 0
+ a0 = 2.4935296
+ a1 = 0
+ a2 = 1
+ toxref = 3e-9
+ b0 = 0
+ b1 = 0
+ at = 72000
+ cf = 8.741900000000001e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.00052197993
+ k3 = -2.5823
+ em = 20000000.0
+ aigbinv = 0.009974
+ minv = -0.33
+ ll = 0
+ lw = 0
+ u0 = 0.009514619299999999
+ w0 = 0
+ ua = 1.4218267e-10
+ ub = 1.1900227e-18
+ uc = 2.2715501e-11
+ ud = 0
+ dmcgt = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 2.33e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ tcjsw = 9.34e-5
+ ndep = 1e+18
+ ijthsfwd = 0.01
+ lwlc = 0
+ moin = 5.5538
+ nigc = 2.291
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ bigsd = 0.0003327
+ ltvoff = 0
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ ijthsrev = 0.01
+ wvoff = 5.5905393e-9
+ poxedge = 1
+ wvsat = -0.0097711764
+ wvth0 = 1.4846626e-8
+ ntox = 2.958
+ pcit = 1e-18
+ pclm = 1.5174437
+ binunit = 2
+ lku0we = 1.8e-11
+ wtvfbsdoff = 0
+ waigc = 3.5172206e-12
+ epsrox = 3.9
+ phin = 0.15
+ lketa = 0
+ rdsmod = 0
+ ltvfbsdoff = 0
+ ppdiblc2 = 0
+ pkt1 = 5e-17
+ xpart = 1
+ igbmod = 1
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ egidl = 0.001
+ pbswgd = 0.8
+ pbswgs = 0.8
+ rbdb = 50
+ prwb = 0
+ prwg = 0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ igcmod = 1
+ rbsb = 50
+ pvag = 2.1
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ rdsw = 200
+ ptvfbsdoff = 0
+ pkvth0we = 0.0
+ vfbsdoff = 0.01
+ rshg = 14.1
+ pvoff = -2.5e-17
+ cdscb = 0
+ cdscd = 0
+ permod = 1
+ pvsat = 0
+ wk2we = 0.0
+ pvth0 = 1.5e-16
+ paramchk = 1
+ njtsswg = 6.489
+ drout = 0.56
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ voffl = 0
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.0026324684
+ weta0 = -1.9361431e-9
+ tnom = 25
+ pdiblcb = 0
+ wetab = 6.0440267e-8
+ voffcv = -0.125
+ wpemod = 1
+ lpclm = 0
+ toxe = 2.6300000000000002e-9
+ toxm = 2.67e-9
+ ijthdfwd = 0.01
+ cgidl = 1
+ bigbacc = 0.0054401
+ wags = 1.128996e-7
+ ijthdrev = 0.01
+ pbswd = 0.9
+ pbsws = 0.9
+ kvth0we = -0.00022
+ lpdiblc2 = 0
+ voff = -0.11172412
+ tpbswg = 0.001
+ acde = 0.5
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ )

.model pch_ff_10 pmos (
+ level = 54
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ lags = 3.1017116e-7
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = -2e-11
+ nfactor = 1
+ kt1l = 0
+ paramchk = 1
+ scref = 1e-6
+ pigcd = 2.572
+ aigsd = 0.0063633879
+ lint = 6.5375218e-9
+ lkt1 = -4.1307452e-8
+ lkt2 = -8.3161855e-9
+ lmax = 9.00077e-6
+ lvoff = -7.1040424e-9
+ lmin = 9.0075e-7
+ lpe0 = 6.44e-8
+ lpeb = 0
+ lvsat = -0.00028
+ lvth0 = -4.1817634e-9
+ ijthdfwd = 0.01
+ toxref = 3e-9
+ nigbacc = 10
+ minv = -0.33
+ delta = 0.018814
+ lua1 = 2.9697696e-17
+ lub1 = 1.2607181e-25
+ luc1 = -4.744495e-18
+ laigc = -4.752933e-11
+ wtvfbsdoff = 0
+ ndep = 1e+18
+ rnoia = 0
+ rnoib = 0
+ lute = -8.6179201e-9
+ lwlc = 0
+ tvfbsdoff = 0.1
+ moin = 5.5538
+ ltvfbsdoff = 0
+ pketa = -2.2807538e-14
+ nigc = 2.291
+ ngate = 1.7e+20
+ ijthdrev = 0.01
+ nigbinv = 2.171
+ ngcon = 1
+ wpclm = -3.01194e-7
+ lpdiblc2 = 7.3300428e-9
+ ltvoff = -4.2514859e-10
+ gbmin = 1e-12
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ pags = -3.4942959e-14
+ ntox = 2.958
+ pcit = 1e-18
+ pclm = 1.5174437
+ fnoimod = 1
+ wvfbsdoff = 0
+ lku0we = 1.8e-11
+ ptvfbsdoff = 0
+ eigbinv = 1.1
+ lvfbsdoff = 0
+ epsrox = 3.9
+ phin = 0.15
+ lkvth0we = 3e-12
+ pkt1 = 9.068958600000001e-15
+ pkt2 = -4.3236504e-15
+ rdsmod = 0
+ igbmod = 1
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ tvoff = 0.0026738399
+ pbswgd = 0.8
+ acnqsmod = 0
+ pbswgs = 0.8
+ rbdb = 50
+ pua1 = 9.6044121e-22
+ prwb = 0
+ pub1 = -1.3952204e-30
+ prwg = 0
+ puc1 = 1.1914589e-22
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ pute = 7.7612988e-14
+ igcmod = 1
+ cigbacc = 0.245
+ rdsw = 200
+ rbodymod = 0
+ tnoimod = 0
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = 6e-10
+ cigbinv = 0.006
+ ppclm = 0
+ paigsd = 3.3403436e-20
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ rshg = 14.1
+ version = 4.5
+ wpdiblc2 = 5.6393415e-10
+ permod = 1
+ tempmod = 0
+ ags = 0.79088496
+ dmcgt = 0
+ cjd = 0.0012517799999999999
+ cit = 5e-6
+ cjs = 0.0012517799999999999
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ tcjsw = 9.34e-5
+ dlc = 1.0572421799999999e-8
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ aigbacc = 0.012071
+ tnom = 25
+ la0 = -3.6651331e-7
+ toxe = 2.6300000000000002e-9
+ toxm = 2.67e-9
+ jsd = 1.5e-7
+ voffcv = -0.125
+ wpemod = 1
+ jss = 1.5e-7
+ lat = -0.0008
+ kt1 = -0.16526426
+ kt2 = -0.046114462
+ lk2 = 4.1045047999999995e-9
+ llc = 0
+ lln = 1
+ bigsd = 0.0003327
+ lu0 = -1.3144212000000002e-10
+ mjd = 0.335
+ mjs = 0.335
+ lua = -1.1601528e-16
+ lub = 1.1870612e-25
+ luc = 1.7407612e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = -2.3980423e-13
+ wkvth0we = 0.0
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ pk2 = -1.7678537e-15
+ aigbinv = 0.009974
+ wvoff = 6.4925381e-9
+ pu0 = 1.0845918e-15
+ prt = 0
+ pua = 1.4359661e-22
+ pub = 1.4495718e-31
+ puc = -1.3724663e-23
+ pud = 0
+ trnqsmod = 0
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 1.2300502e-9
+ ub1 = -1.4464065e-18
+ uc1 = 7.8962019e-11
+ wvsat = -0.0097711764
+ tpb = 0.0016
+ wvth0 = 1.5492791199999998e-8
+ wa0 = 3.6413271e-7
+ ute = -0.99031694
+ wags = 1.1678647e-7
+ web = 6628.3
+ wec = -16935.0
+ wk2 = -2.0904063e-9
+ wlc = 0
+ wln = 1
+ wu0 = -2.0727529e-10
+ xgl = -8.2e-9
+ waigc = 4.3868453e-12
+ xgw = 0
+ wua = -1.2839182e-16
+ wub = -8.3225053e-26
+ wuc = -2.1668301e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ voff = -0.11093391
+ acde = 0.5
+ tpbswg = 0.001
+ lketa = -1.0921036e-8
+ vsat = 121084.96
+ wint = 0
+ xpart = 1
+ vth0 = -0.3649855
+ rgatemod = 0
+ wkt1 = -1.1364676e-8
+ wkt2 = -3.3960513e-9
+ poxedge = 1
+ wmax = 8.9974e-6
+ tnjtsswg = 1
+ aigc = 0.0068356471
+ wmin = 8.974e-7
+ egidl = 0.001
+ binunit = 2
+ ptvoff = -4.5667618e-16
+ waigsd = 1.9102262e-12
+ wua1 = -4.3482598e-16
+ wub1 = 7.4750944e-25
+ wuc1 = -1.0064978e-16
+ bigc = 0.0012521
+ wute = -8.7205605e-8
+ diomod = 1
+ wwlc = 0
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.6832999999999998e-10
+ pku0we = 0.0
+ cjswgs = 1.6832999999999998e-10
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.2212350000000004e-11
+ cgdo = 2.8335740000000002e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.2212350000000004e-11
+ cgso = 2.8335740000000002e-11
+ cigc = 0.15259
+ pvoff = -8.133969200000001e-15
+ jtsswgd = 1.75e-7
+ pvfbsdoff = 0
+ mjswgd = 0.95
+ jtsswgs = 1.75e-7
+ mjswgs = 0.95
+ cdscb = 0
+ cdscd = 0
+ tcjswg = 0.00128
+ pvsat = 0
+ wk2we = 0.0
+ pvth0 = -5.658937700000001e-15
+ drout = 0.56
+ paigc = -7.8179264e-18
+ a0 = 2.5342986
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 72000
+ cf = 8.741900000000001e-11
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.0010230372
+ k3 = -2.5823
+ em = 20000000.0
+ voffl = 0
+ ll = 0
+ lw = 0
+ u0 = 0.0095279054
+ w0 = 0
+ ua = 1.5508759e-10
+ ub = 1.1768184e-18
+ uc = 2.077917e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 2.33e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ weta0 = -1.9361431e-9
+ wetab = 6.0440267e-8
+ k2we = 5e-5
+ lpclm = 0
+ dsub = 0.5
+ dtox = 3.91e-10
+ ijthsfwd = 0.01
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ njtsswg = 6.489
+ cgidl = 1
+ fprout = 200
+ xrcrg1 = 12
+ xrcrg2 = 1
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ eta0 = 0.16744607
+ etab = -0.23671111
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.0018171133
+ pdiblcb = 0
+ pbswd = 0.9
+ wtvoff = -4.8127407e-11
+ pbsws = 0.9
+ ijthsrev = 0.01
+ pdits = 0
+ capmod = 2
+ cigsd = 0.013281
+ wku0we = 1.5e-11
+ bigbacc = 0.0054401
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ mobmod = 0
+ ppdiblc2 = -1.7911725e-15
+ kvth0we = -0.00022
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ tnoia = 0
+ peta0 = 2e-17
+ wketa = 2.4899578e-8
+ laigsd = -3.7090202e-15
+ tpbsw = 0.0025
+ pkvth0we = 0.0
+ cjswd = 4.743e-11
+ cjsws = 4.743e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ keta = -0.04361839
+ vfbsdoff = 0.01
+ )

.model pch_ff_11 pmos (
+ level = 54
+ egidl = 0.001
+ ltvfbsdoff = 0
+ toxref = 3e-9
+ ijthsfwd = 0.01
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ tnom = 25
+ toxe = 2.6300000000000002e-9
+ toxm = 2.67e-9
+ ijthsrev = 0.01
+ ptvfbsdoff = 0
+ ltvoff = -2.603747e-10
+ pvfbsdoff = 0
+ wags = -5.7105665e-9
+ pvoff = 6.0260933999999995e-15
+ cdscb = 0
+ cdscd = 0
+ pvsat = 0
+ wk2we = 0.0
+ voff = -0.10782222
+ njtsswg = 6.489
+ pvth0 = 3.3963831e-15
+ drout = 0.56
+ acde = 0.5
+ paigc = 1.0166993e-17
+ lku0we = 1.8e-11
+ xtsswgd = 0.32
+ vsat = 121084.96
+ xtsswgs = 0.32
+ wint = 0
+ ppdiblc2 = 8.932051e-16
+ vth0 = -0.36648038999999993
+ epsrox = 3.9
+ voffl = 0
+ wkt1 = 3.9882501e-9
+ wkt2 = -1.3862366e-8
+ ckappad = 0.6
+ wmax = 8.9974e-6
+ ckappas = 0.6
+ aigc = 0.0068328167
+ wmin = 8.974e-7
+ pdiblc1 = 0
+ pdiblc2 = 0.0082016634
+ pdiblcb = 0
+ weta0 = -1.9361431e-9
+ rdsmod = 0
+ wetab = 6.0440267e-8
+ igbmod = 1
+ lpclm = 0
+ wua1 = 1.0350058e-15
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ wub1 = -1.41997e-24
+ wuc1 = 5.1522417e-17
+ cgidl = 1
+ pbswgd = 0.8
+ bigc = 0.0012521
+ pbswgs = 0.8
+ wwlc = 0
+ bigbacc = 0.0054401
+ igcmod = 1
+ pkvth0we = 0.0
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.2212350000000004e-11
+ cgdo = 2.8335740000000002e-11
+ xtid = 3
+ xtis = 3
+ pbswd = 0.9
+ pbsws = 0.9
+ kvth0we = -0.00022
+ cgsl = 3.2212350000000004e-11
+ cgso = 2.8335740000000002e-11
+ cigc = 0.15259
+ vfbsdoff = 0.01
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ pdits = 0
+ cigsd = 0.013281
+ paigsd = -3.7089273e-20
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ paramchk = 1
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ permod = 1
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ k2we = 5e-5
+ tnoia = 0
+ dsub = 0.5
+ dtox = 3.91e-10
+ ijthdfwd = 0.01
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ peta0 = 2e-17
+ voffcv = -0.125
+ wpemod = 1
+ wketa = -2.3248862e-8
+ tpbsw = 0.0025
+ eta0 = 0.16744607
+ nfactor = 1
+ etab = -0.23671111
+ cjswd = 4.743e-11
+ cjsws = 4.743e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ ijthdrev = 0.01
+ lpdiblc2 = 1.6477933e-9
+ nigbacc = 10
+ tpbswg = 0.001
+ scref = 1e-6
+ pigcd = 2.572
+ aigsd = 0.0063633394
+ lvoff = -9.8734428e-9
+ nigbinv = 2.171
+ ptvoff = 2.6240046e-16
+ lkvth0we = 3e-12
+ waigsd = 1.9894315e-12
+ lvsat = -0.00028
+ lvth0 = -2.8513091000000003e-9
+ delta = 0.018814
+ diomod = 1
+ laigc = -4.5010295e-11
+ acnqsmod = 0
+ rnoia = 0
+ rnoib = 0
+ tvfbsdoff = 0.1
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.6832999999999998e-10
+ pku0we = 0.0
+ cjswgs = 1.6832999999999998e-10
+ fnoimod = 1
+ pketa = 2.0044574e-14
+ rbodymod = 0
+ ngate = 1.7e+20
+ eigbinv = 1.1
+ ngcon = 1
+ wpclm = -3.01194e-7
+ keta = -0.035478054
+ mjswgd = 0.95
+ mjswgs = 0.95
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ tcjswg = 0.00128
+ lags = 2.7680102e-7
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 6.2671111e-11
+ kt1l = 0
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ wpdiblc2 = -2.4522204e-9
+ lint = 6.5375218e-9
+ cigbacc = 0.245
+ lkt1 = -1.3922155e-8
+ lkt2 = -7.1896716e-9
+ lmax = 9.0075e-7
+ lmin = 4.5075e-7
+ tnoimod = 0
+ lpe0 = 6.44e-8
+ lpeb = 0
+ fprout = 200
+ minv = -0.33
+ cigbinv = 0.006
+ lua1 = 8.7159171e-17
+ lub1 = -2.6689299e-25
+ luc1 = 2.9116076e-17
+ tvoff = 0.0024887007
+ xrcrg1 = 12
+ xrcrg2 = 1
+ ndep = 1e+18
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ lwlc = 0
+ moin = 5.5538
+ wkvth0we = 0.0
+ wtvoff = -8.5607868e-10
+ nigc = 2.291
+ version = 4.5
+ a0 = 2.8862723
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ trnqsmod = 0
+ at = 72000
+ cf = 8.741900000000001e-11
+ tempmod = 0
+ ef = 1.15
+ ku0we = -0.0007
+ k1 = 0.30425
+ k2 = 0.0046668319
+ k3 = -2.5823
+ em = 20000000.0
+ ll = 0
+ lw = 0
+ beta0 = 13.32
+ u0 = 0.0095144338
+ w0 = 0
+ ua = 8.4190146e-11
+ ub = 1.1838278e-18
+ uc = 4.9200634e-11
+ ud = 0
+ leta0 = 6e-10
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 2.33e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ capmod = 2
+ ppclm = 0
+ aigbacc = 0.012071
+ wku0we = 1.5e-11
+ pags = 7.4079401e-14
+ ags = 0.8283795
+ dlcig = 2.5e-9
+ mobmod = 0
+ bgidl = 1834800000.0
+ ntox = 2.958
+ pcit = 1e-18
+ pclm = 1.5174437
+ cjd = 0.0012517799999999999
+ cit = -8.7888889e-5
+ cjs = 0.0012517799999999999
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 1.0572421799999999e-8
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ rgatemod = 0
+ tnjtsswg = 1
+ phin = 0.15
+ aigbinv = 0.009974
+ dmcgt = 0
+ la0 = -6.797699e-7
+ pkt1 = -4.5951461000000004e-15
+ jsd = 1.5e-7
+ pkt2 = 4.9913693e-15
+ tcjsw = 9.34e-5
+ jss = 1.5e-7
+ lat = -0.0008
+ kt1 = -0.19603426
+ kt2 = -0.047380208
+ lk2 = -9.594787e-10
+ llc = 0
+ lln = 1
+ lu0 = -1.1945246e-10
+ mjd = 0.335
+ mjs = 0.335
+ lua = -5.2916554e-17
+ lub = 1.1246778e-25
+ luc = -7.8874906e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 4.0323955e-14
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ pk2 = 1.1838025e-15
+ pu0 = -8.8186737e-16
+ laigsd = 3.9492818e-14
+ prt = 0
+ pua = -2.1071339e-22
+ pub = -4.1382897e-32
+ puc = 1.6409308e-23
+ pud = 0
+ rbdb = 50
+ pua1 = -3.4770908e-22
+ prwb = 0
+ pub1 = 5.3383631e-31
+ prwg = 0
+ rsh = 15.2
+ puc1 = -1.6287371e-23
+ tcj = 0.000832
+ ua1 = 1.1654868e-9
+ ub1 = -1.004873e-18
+ uc1 = 4.0916434e-11
+ bigsd = 0.0003327
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ tpb = 0.0016
+ wa0 = 4.9381936e-8
+ ute = -1
+ web = 6628.3
+ wec = -16935.0
+ wk2 = -5.406874e-9
+ rdsw = 200
+ wlc = 0
+ wln = 1
+ wu0 = 2.0022293e-9
+ xgl = -8.2e-9
+ wvoff = -9.4176445e-9
+ xgw = 0
+ wua = 2.6970929e-16
+ wub = 1.2614582e-25
+ wuc = -5.5526695e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ poxedge = 1
+ wvsat = -0.0097711764
+ wvth0 = 5.3182589e-9
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ binunit = 2
+ waigc = -1.5820929e-11
+ rshg = 14.1
+ lketa = -1.8165935e-8
+ xpart = 1
+ wtvfbsdoff = 0
+ )

.model pch_ff_12 pmos (
+ level = 54
+ wkvth0we = 0.0
+ pketa = 2.9922765e-15
+ ngate = 1.7e+20
+ ngcon = 1
+ cigbacc = 0.245
+ ltvoff = -1.0992228e-10
+ wpclm = -3.01194e-7
+ trnqsmod = 0
+ gbmin = 1e-12
+ tnoimod = 0
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ cigbinv = 0.006
+ lku0we = 1.8e-11
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ epsrox = 3.9
+ rgatemod = 0
+ tnjtsswg = 1
+ rdsmod = 0
+ version = 4.5
+ igbmod = 1
+ tempmod = 0
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ pbswgd = 0.8
+ pbswgs = 0.8
+ tvoff = 0.0021467634
+ aigbacc = 0.012071
+ igcmod = 1
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ ku0we = -0.0007
+ ags = 0.29253015
+ aigbinv = 0.009974
+ beta0 = 13.32
+ keta = -0.031086208
+ leta0 = 6e-10
+ cjd = 0.0012517799999999999
+ cit = -0.00056559017
+ cjs = 0.0012517799999999999
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 1.38228675e-8
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ lags = 5.1257474e-7
+ ppclm = 0
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 2.7285967e-10
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ kt1l = 0
+ la0 = -1.4357692e-8
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = -0.0008
+ kt1 = -0.19916819
+ kt2 = -0.054700402
+ lk2 = 1.025099e-9
+ permod = 1
+ llc = -1.18e-13
+ lln = 0.7
+ lu0 = -4.9276045e-10
+ mjd = 0.335
+ mjs = 0.335
+ lua = -1.6078561e-16
+ lub = 5.7693033e-26
+ luc = -4.8483261e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ lint = 9.7879675e-9
+ pa0 = -2.613694e-13
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ pk2 = -5.5906497e-16
+ lkt1 = -1.2543223999999999e-8
+ lkt2 = -3.9687861e-9
+ pu0 = -2.2461433e-17
+ lmax = 4.5075e-7
+ prt = 0
+ pua = 5.4100623e-23
+ pub = -6.3187687e-32
+ puc = -3.6550877e-24
+ pud = 0
+ dmcgt = 0
+ lmin = 2.1744e-7
+ poxedge = 1
+ tcjsw = 9.34e-5
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 1.2176874e-9
+ ub1 = -1.2376668e-18
+ lpe0 = 6.44e-8
+ uc1 = 1.0272662e-10
+ lpeb = 0
+ tpb = 0.0016
+ wa0 = 7.3504866e-7
+ ijthsfwd = 0.01
+ ute = -1
+ web = 6628.3
+ wec = -16935.0
+ wk2 = -1.4458115e-9
+ binunit = 2
+ voffcv = -0.125
+ wpemod = 1
+ wlc = 0
+ wln = 1
+ minv = -0.33
+ wu0 = 4.9034036e-11
+ xgl = -8.2e-9
+ xgw = 0
+ lua1 = 6.4190903e-17
+ lub1 = -1.6446372e-25
+ wua = -3.3214073e-16
+ wub = 1.7570216e-25
+ wuc = -9.9257962e-18
+ wud = 0
+ luc1 = 1.9195943e-18
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ ndep = 1e+18
+ bigsd = 0.0003327
+ lwlc = 0
+ moin = 5.5538
+ wvoff = 6.3544834e-9
+ nigc = 2.291
+ ijthsrev = 0.01
+ wvsat = -0.0097711764
+ wvth0 = 1.2177300389999999e-8
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ waigc = 4.9938134e-12
+ tpbswg = 0.001
+ jtsswgd = 1.75e-7
+ pags = 2.5662868e-13
+ jtsswgs = 1.75e-7
+ ntox = 2.958
+ pcit = -8.0677938e-17
+ lketa = -2.0098347e-8
+ pclm = 1.5174437
+ xpart = 1
+ ppdiblc2 = -1.9289508e-16
+ phin = 0.15
+ ptvoff = -6.733506e-17
+ egidl = 0.001
+ waigsd = 1.9051377e-12
+ pkt1 = 5.4381461e-16
+ pkt2 = -1.2251691e-15
+ diomod = 1
+ pditsd = 0
+ pditsl = 0
+ rbdb = 50
+ cjswgd = 1.6832999999999998e-10
+ pku0we = 0.0
+ pua1 = -4.1586322e-23
+ prwb = 0
+ pub1 = 2.600258e-32
+ prwg = 0
+ cjswgs = 1.6832999999999998e-10
+ puc1 = -8.5761835e-25
+ njtsswg = 6.489
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ pkvth0we = 0.0
+ rdsw = 200
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ ckappad = 0.6
+ ckappas = 0.6
+ mjswgd = 0.95
+ mjswgs = 0.95
+ pdiblc1 = 0
+ pdiblc2 = 0.01380092
+ pvfbsdoff = 0
+ pdiblcb = 0
+ vfbsdoff = 0.01
+ pvoff = -9.136429e-16
+ tcjswg = 0.00128
+ cdscb = 0
+ cdscd = 0
+ pvsat = 0
+ wk2we = 0.0
+ pvth0 = 3.7840375e-16
+ drout = 0.56
+ paramchk = 1
+ rshg = 14.1
+ paigc = 1.0085061e-18
+ bigbacc = 0.0054401
+ voffl = 0
+ weta0 = -1.9361431e-9
+ kvth0we = -0.00022
+ wetab = 6.0440267e-8
+ lpclm = 0
+ lintnoi = -5e-9
+ fprout = 200
+ ijthdfwd = 0.01
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ xrcrg1 = 12
+ xrcrg2 = 1
+ cgidl = 1
+ tnom = 25
+ toxe = 2.6300000000000002e-9
+ toxm = 2.67e-9
+ wtvoff = -1.0667978e-10
+ pbswd = 0.9
+ pbsws = 0.9
+ ijthdrev = 0.01
+ lpdiblc2 = -8.1587971e-10
+ capmod = 2
+ wags = -4.2059528e-7
+ wku0we = 1.5e-11
+ wcit = 1.8563168e-10
+ pdits = 0
+ cigsd = 0.013281
+ mobmod = 0
+ voff = -0.12166106
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ acde = 0.5
+ vsat = 121084.96
+ wint = 0
+ vth0 = -0.38344941
+ nfactor = 1
+ pk2we = 0.0
+ wkt1 = -7.6912059e-9
+ wkt2 = 2.6613072e-10
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ wmax = 8.9974e-6
+ aigc = 0.0067878654
+ wmin = 8.974e-7
+ lkvth0we = 3e-12
+ tnoia = 0
+ a0 = 1.3739719
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 72000
+ wua1 = 3.3927227e-16
+ cf = 8.741900000000001e-11
+ wub1 = -2.6580249e-25
+ wuc1 = 1.6454797e-17
+ ef = 1.15
+ k1 = 0.30425
+ k2 = 0.00015642806
+ k3 = -2.5823
+ em = 20000000.0
+ peta0 = 2e-17
+ ll = -1.18e-13
+ lw = 0
+ u0 = 0.010362861
+ w0 = 0
+ ua = 3.293471e-10
+ ub = 1.3083159e-18
+ uc = 4.2293442e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 2.33e-9
+ ww = 0
+ bigc = 0.0012521
+ xw = 8.600000000000001e-9
+ wketa = 1.5506359e-8
+ wwlc = 0
+ acnqsmod = 0
+ tpbsw = 0.0025
+ nigbacc = 10
+ cjswd = 4.743e-11
+ cjsws = 4.743e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ cdsc = 0
+ cgbo = 0
+ rbodymod = 0
+ cgdl = 3.2212350000000004e-11
+ cgdo = 2.8335740000000002e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.2212350000000004e-11
+ cgso = 2.8335740000000002e-11
+ cigc = 0.15259
+ wtvfbsdoff = 0
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ nigbinv = 2.171
+ ltvfbsdoff = 0
+ scref = 1e-6
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ pigcd = 2.572
+ wpdiblc2 = 1.6189099e-11
+ aigsd = 0.0063634291
+ fnoimod = 1
+ lvoff = -3.7843526e-9
+ eigbinv = 1.1
+ k2we = 5e-5
+ toxref = 3e-9
+ lvsat = -0.00028
+ dsub = 0.5
+ dtox = 3.91e-10
+ lvth0 = 4.6151015e-9
+ ptvfbsdoff = 0
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ delta = 0.018814
+ laigc = -2.5231709e-11
+ tvfbsdoff = 0.1
+ rnoia = 0
+ rnoib = 0
+ eta0 = 0.16744607
+ etab = -0.23671111
+ )

.model pch_ff_13 pmos (
+ level = 54
+ pags = 7.0037917e-14
+ lku0we = 1.8e-11
+ pvth0 = -6.538291000000006e-17
+ drout = 0.56
+ epsrox = 3.9
+ ntox = 2.958
+ pcit = 3.2250046e-17
+ pclm = 1.5924795
+ paigc = -7.3857349e-19
+ voffl = 0
+ rdsmod = 0
+ phin = 0.15
+ igbmod = 1
+ weta0 = -1.9361431e-9
+ wetab = 6.0440267e-8
+ lkvth0we = 3e-12
+ pkt1 = 3.3071967000000004e-16
+ pkt2 = -8.6151083e-16
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ lpclm = -1.5832542e-8
+ pbswgd = 0.8
+ pbswgs = 0.8
+ cgidl = 1
+ igcmod = 1
+ acnqsmod = 0
+ rbdb = 50
+ pua1 = -5.7774504e-23
+ prwb = 0
+ pub1 = 1.0356474e-31
+ prwg = 0
+ puc1 = 6.0450908e-24
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ rdsw = 200
+ rbodymod = 0
+ pbswd = 0.9
+ pbsws = 0.9
+ nfactor = 1
+ pdits = 0
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ permod = 1
+ rshg = 14.1
+ nigbacc = 10
+ wpdiblc2 = -2.9527442e-9
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ tnoia = 0
+ voffcv = -0.125
+ wpemod = 1
+ nigbinv = 2.171
+ peta0 = 2e-17
+ tnom = 25
+ wketa = 2.8638443e-8
+ toxe = 2.6300000000000002e-9
+ toxm = 2.67e-9
+ tpbsw = 0.0025
+ cjswd = 4.743e-11
+ cjsws = 4.743e-11
+ mjswd = 0.01
+ wkvth0we = 0.0
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ trnqsmod = 0
+ fnoimod = 1
+ eigbinv = 1.1
+ wags = 4.6372111e-7
+ tpbswg = 0.001
+ wcit = -3.4957204e-10
+ voff = -0.13366619
+ acde = 0.5
+ scref = 1e-6
+ vsat = 121978.39
+ wint = 0
+ vth0 = -0.38524102000000005
+ rgatemod = 0
+ pigcd = 2.572
+ aigsd = 0.0063634291
+ wkt1 = -6.6812774e-9
+ wkt2 = -1.4573681e-9
+ tnjtsswg = 1
+ ptvoff = -1.8786066e-17
+ wmax = 8.9974e-6
+ aigc = 0.0067673585
+ wmin = 8.974e-7
+ lvoff = -1.2512704e-9
+ waigsd = 1.9051377e-12
+ cigbacc = 0.245
+ lvsat = -0.00046849676999999995
+ diomod = 1
+ lvth0 = 4.9931296e-9
+ wua1 = 4.1599351e-16
+ wub1 = -6.3339564e-25
+ wuc1 = -1.6259465e-17
+ tnoimod = 0
+ delta = 0.018814
+ laigc = -2.090475e-11
+ pditsd = 0
+ pditsl = 0
+ tvfbsdoff = 0.1
+ bigc = 0.0012521
+ cjswgd = 1.6832999999999998e-10
+ pku0we = 0.0
+ cjswgs = 1.6832999999999998e-10
+ wwlc = 0
+ rnoia = 0
+ rnoib = 0
+ cigbinv = 0.006
+ cdsc = 0
+ pketa = 2.2140676e-16
+ ngate = 1.7e+20
+ cgbo = 0
+ cgdl = 3.2212350000000004e-11
+ cgdo = 2.8335740000000002e-11
+ xtid = 3
+ xtis = 3
+ ngcon = 1
+ mjswgd = 0.95
+ cgsl = 3.2212350000000004e-11
+ cgso = 2.8335740000000002e-11
+ mjswgs = 0.95
+ wpclm = -3.6917638e-7
+ cigc = 0.15259
+ tcjswg = 0.00128
+ version = 4.5
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ tempmod = 0
+ jswgs = 3.69e-13
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ aigbacc = 0.012071
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ k2we = 5e-5
+ fprout = 200
+ aigbinv = 0.009974
+ dsub = 0.5
+ dtox = 3.91e-10
+ xrcrg1 = 12
+ xrcrg2 = 1
+ ijthsfwd = 0.01
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ tvoff = 0.0019304691
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ ags = 2.6061153
+ wtvoff = -3.3676979e-10
+ eta0 = 0.16744607
+ etab = -0.23671111
+ cjd = 0.0012517799999999999
+ cit = 0.00047888384
+ cjs = 0.0012517799999999999
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 1.38228675e-8
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ ijthsrev = 0.01
+ ku0we = -0.0007
+ beta0 = 13.32
+ capmod = 2
+ leta0 = 6e-10
+ la0 = -4.2186937e-8
+ poxedge = 1
+ wku0we = 1.5e-11
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = -0.00051178856
+ kt1 = -0.23884145
+ kt2 = -0.071460529
+ lk2 = 3.928829499999999e-9
+ llc = -1.18e-13
+ lln = 0.7
+ lu0 = -1.9651509e-10
+ mjd = 0.335
+ ppclm = 1.4344283e-14
+ mjs = 0.335
+ lua = -2.3141614e-17
+ lub = -3.0092793e-26
+ luc = -1.1168748e-18
+ lud = 0
+ lwc = 0
+ mobmod = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = -1.7418058e-15
+ nsd = 1e+20
+ binunit = 2
+ pbd = 0.75
+ pat = -2.5956322e-9
+ pbs = 0.75
+ pk2 = -2.0925962e-16
+ dlcig = 2.5e-9
+ pu0 = 6.8306111e-19
+ bgidl = 1834800000.0
+ prt = 0
+ pua = -2.4112447e-23
+ pub = 3.4375734e-32
+ puc = -1.1236355e-25
+ pud = 0
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 2.2048659e-9
+ ub1 = -2.7884819e-18
+ ppdiblc2 = 4.3354985e-16
+ uc1 = 8.0779763e-11
+ tpb = 0.0016
+ wa0 = -4.9541389e-7
+ ute = -1
+ wat = 0.012301575
+ web = 6628.3
+ wec = -16935.0
+ wk2 = -3.1036812e-9
+ wlc = 0
+ wln = 1
+ wu0 = -6.065551e-11
+ xgl = -8.2e-9
+ xgw = 0
+ wua = 3.8537331e-17
+ wub = -2.8668372e-25
+ wuc = -2.6715958e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ wtvfbsdoff = 0
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ bigsd = 0.0003327
+ ltvfbsdoff = 0
+ pkvth0we = 0.0
+ wvoff = 5.8569161e-9
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ wvsat = -0.0105806259
+ vfbsdoff = 0.01
+ keta = -0.13181891
+ wvth0 = 1.42805795e-8
+ waigc = 1.3273811e-11
+ lags = 2.4408277e-8
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 5.2475659000000004e-11
+ a0 = 1.505864
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ kt1l = 0
+ ptvfbsdoff = 0
+ at = 70634.069
+ paramchk = 1
+ cf = 8.741900000000001e-11
+ lketa = 1.156253e-9
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.013605325
+ k3 = -2.5823
+ em = 20000000.0
+ ll = -1.18e-13
+ lw = 0
+ u0 = 0.0089588547
+ w0 = 0
+ xpart = 1
+ ua = -3.2299413e-10
+ ub = 1.7243624e-18
+ uc = 2.4608838e-11
+ ud = 0
+ njtsswg = 6.489
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 2.33e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ lint = 9.7879675e-9
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ lkt1 = -4.1721668999999995e-9
+ lkt2 = -4.3239941e-10
+ egidl = 0.001
+ lmax = 2.1744e-7
+ lmin = 9.167e-8
+ toxref = 3e-9
+ ckappad = 0.6
+ ckappas = 0.6
+ lpe0 = 6.44e-8
+ pdiblc1 = 0
+ pdiblc2 = 0.017260131
+ lpeb = 0
+ pdiblcb = 0
+ ijthdfwd = 0.01
+ minv = -0.33
+ lua1 = -1.4410376e-16
+ lub1 = 1.6275827e-25
+ luc1 = 6.550381e-18
+ ndep = 1e+18
+ lwlc = 0
+ moin = 5.5538
+ bigbacc = 0.0054401
+ nigc = 2.291
+ ltvoff = -6.4284173e-11
+ ijthdrev = 0.01
+ pvfbsdoff = 0
+ lpdiblc2 = -1.5457732e-9
+ kvth0we = -0.00022
+ pvoff = -8.086562e-16
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ cdscb = 0
+ cdscd = 0
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ pvsat = 1.7077360999999997e-10
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ wk2we = 0.0
+ )

.model pch_ff_14 pmos (
+ level = 54
+ cjd = 0.0012517799999999999
+ poxedge = 1
+ cit = 7.175354000000004e-5
+ wua1 = -1.4703955e-15
+ cjs = 0.0012517799999999999
+ clc = 1e-7
+ cle = 0.6
+ wub1 = 2.631826e-24
+ bvd = 8.2
+ wuc1 = 2.762344e-16
+ bvs = 8.2
+ igcmod = 1
+ dlc = 4.0349e-9
+ k3b = 2.1176
+ tvoff = 0.0011122833
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ bigc = 0.0012521
+ wwlc = 0
+ xjbvd = 1
+ binunit = 2
+ xjbvs = 1
+ lk2we = 0.0
+ pkvth0we = 0.0
+ la0 = -2.3326483e-7
+ jsd = 1.5e-7
+ cdsc = 0
+ jss = 1.5e-7
+ lat = -0.0073502639
+ kt1 = -0.2764195
+ kt2 = -0.075556865
+ lk2 = 3.4809157e-9
+ llc = 0
+ cgbo = 0
+ lln = 1
+ cgdl = 3.2212350000000004e-11
+ cgdo = 2.8335740000000002e-11
+ lu0 = 1.9444492e-10
+ xtid = 3
+ xtis = 3
+ mjd = 0.335
+ mjs = 0.335
+ lua = 5.4621428e-17
+ lub = 1.7088257e-26
+ luc = 1.0238844e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ cgsl = 3.2212350000000004e-11
+ njs = 1.02
+ cgso = 2.8335740000000002e-11
+ pa0 = 5.4920056e-14
+ cigc = 0.15259
+ ku0we = -0.0007
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 1.0391973e-9
+ pbs = 0.75
+ pk2 = 6.854543e-16
+ beta0 = 13.32
+ vfbsdoff = 0.01
+ pu0 = -1.2707891e-16
+ leta0 = -4.8260389999999976e-11
+ prt = 0
+ pua = -5.2218942e-24
+ pub = -4.7511951e-32
+ puc = -9.869134e-24
+ pud = 0
+ letab = 2.0996791e-8
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 8.9078668e-10
+ ub1 = -1.404024e-18
+ uc1 = 4.4088848e-11
+ ppclm = 7.4853015e-14
+ tpb = 0.0016
+ wa0 = -1.0981997e-6
+ ute = -1
+ wat = -0.026366825
+ web = 6628.3
+ wec = -16935.0
+ wk2 = -1.2621914e-8
+ wlc = 0
+ dlcig = 2.5e-9
+ permod = 1
+ wln = 1
+ wu0 = 1.2985144e-9
+ xgl = -8.2e-9
+ xgw = 0
+ bgidl = 1834800000.0
+ wua = -1.62426e-16
+ wub = 5.8446154e-25
+ wuc = 7.7079472e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ paramchk = 1
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ k2we = 5e-5
+ voffcv = -0.125
+ wpemod = 1
+ dsub = 0.5
+ dtox = 3.91e-10
+ ijthdfwd = 0.01
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ bigsd = 0.0003327
+ eta0 = 0.17434246
+ etab = -0.46008122
+ njtsswg = 6.489
+ wvoff = -4.5993296e-9
+ ijthdrev = 0.01
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ wvsat = -0.015871066
+ wvth0 = 6.483999e-9
+ lpdiblc2 = 0
+ ckappad = 0.6
+ tpbswg = 0.001
+ ckappas = 0.6
+ waigc = -2.1370578e-11
+ pdiblc1 = 0
+ pdiblc2 = 0.00081573526
+ pdiblcb = 0
+ lketa = 9.0137227e-9
+ xpart = 1
+ ptvoff = 1.200911e-16
+ waigsd = 1.9051377e-12
+ bigbacc = 0.0054401
+ egidl = 0.001
+ lkvth0we = 3e-12
+ diomod = 1
+ kvth0we = -0.00022
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.6832999999999998e-10
+ pku0we = 0.0
+ cjswgs = 1.6832999999999998e-10
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ acnqsmod = 0
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ rbodymod = 0
+ mjswgd = 0.95
+ mjswgs = 0.95
+ pvfbsdoff = 0
+ tcjswg = 0.00128
+ keta = -0.21540901
+ pvoff = 1.7423089e-16
+ cdscb = 0
+ cdscd = 0
+ lags = -3.1969346e-8
+ pvsat = 6.680730999999999e-10
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ wk2we = 0.0
+ pvth0 = 6.674869e-16
+ lcit = 9.074578e-11
+ drout = 0.56
+ kt1l = 0
+ paigc = 2.5179991e-18
+ voffl = 0
+ wpdiblc2 = 1.6594883e-9
+ lint = 0
+ lkt1 = -6.398308999999999e-10
+ lkt2 = -4.7343777e-11
+ weta0 = 4.269971e-8
+ nfactor = 1
+ lmax = 9.167e-8
+ wetab = 1.3144359e-7
+ fprout = 200
+ lmin = 5.567e-8
+ lpclm = -1.0675035e-7
+ xrcrg1 = 12
+ xrcrg2 = 1
+ lpe0 = 6.44e-8
+ lpeb = 0
+ cgidl = 1
+ minv = -0.33
+ lua1 = -2.0580314e-17
+ lub1 = 3.261922e-26
+ luc1 = 9.999327e-18
+ wtvoff = -1.8141864e-9
+ ndep = 1e+18
+ lwlc = 0
+ moin = 5.5538
+ wkvth0we = 0.0
+ nigbacc = 10
+ pbswd = 0.9
+ nigc = 2.291
+ pbsws = 0.9
+ capmod = 2
+ trnqsmod = 0
+ wku0we = 1.5e-11
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ mobmod = 0
+ pdits = 0
+ nigbinv = 2.171
+ cigsd = 0.013281
+ pags = 2.8964227e-14
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ wtvfbsdoff = 0
+ ntox = 2.958
+ pcit = -7.543103999999996e-18
+ pclm = 2.5596902
+ rgatemod = 0
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ tnjtsswg = 1
+ ltvfbsdoff = 0
+ phin = 0.15
+ pkt1 = 1.2782004099999999e-16
+ pkt2 = 1.7971063e-15
+ fnoimod = 1
+ tnoia = 0
+ eigbinv = 1.1
+ peta0 = -4.1757701999999996e-15
+ petab = -6.6743123e-15
+ wketa = 8.0928346e-8
+ tpbsw = 0.0025
+ rbdb = 50
+ pua1 = 1.1954606e-22
+ prwb = 0
+ pub1 = -2.033661e-31
+ prwg = 0
+ puc1 = -2.1449333e-23
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ cjswd = 4.743e-11
+ pvag = 2.1
+ cjsws = 4.743e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ rdsw = 200
+ ptvfbsdoff = 0
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ cigbacc = 0.245
+ tnoimod = 0
+ rshg = 14.1
+ scref = 1e-6
+ pigcd = 2.572
+ cigbinv = 0.006
+ aigsd = 0.0063634291
+ lvoff = -2.6816163e-9
+ toxref = 3e-9
+ lvsat = -0.0048652254
+ lvth0 = -8.626699e-10
+ version = 4.5
+ ijthsfwd = 0.01
+ delta = 0.018814
+ tvfbsdoff = 0.1
+ tempmod = 0
+ laigc = -1.5433256e-11
+ tnom = 25
+ toxe = 2.6300000000000002e-9
+ toxm = 2.67e-9
+ rnoia = 0
+ rnoib = 0
+ aigbacc = 0.012071
+ ltvoff = 1.2625293e-11
+ pketa = -4.6938441e-15
+ a0 = 3.5386076
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ ngate = 1.7e+20
+ at = 143383.81
+ cf = 8.741900000000001e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.0088402851
+ k3 = -2.5823
+ ijthsrev = 0.01
+ em = 20000000.0
+ ngcon = 1
+ ll = 0
+ lw = 0
+ u0 = 0.0047997056
+ wpclm = -1.0128863e-6
+ w0 = 0
+ ua = -1.1502605e-9
+ ub = 1.2224364e-18
+ uc = -9.619668e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 2.33e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ gbmin = 1e-12
+ wags = 9.0067526e-7
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ aigbinv = 0.009974
+ wcit = 7.375874999999998e-11
+ lku0we = 1.8e-11
+ wvfbsdoff = 0
+ epsrox = 3.9
+ lvfbsdoff = 0
+ voff = -0.11844975
+ acde = 0.5
+ vsat = 168752.09000000003
+ ppdiblc2 = 0
+ rdsmod = 0
+ wint = 0
+ vth0 = -0.32294523999999997
+ igbmod = 1
+ wkt1 = -4.5227706e-9
+ wkt2 = -2.9740529e-8
+ wmax = 8.9974e-6
+ aigc = 0.0067091511
+ wmin = 8.974e-7
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ pbswgd = 0.8
+ ags = 3.2058772
+ pbswgs = 0.8
+ )

.model pch_ff_15 pmos (
+ level = 54
+ keta = 0.054978601
+ fnoimod = 1
+ pdits = 0
+ eigbinv = 1.1
+ cigsd = 0.013281
+ permod = 1
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 8.916000000000024e-12
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ kt1l = 0
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ lint = 0
+ lkt1 = -1.3008111999999999e-8
+ lkt2 = 1.0752811e-9
+ lmax = 5.567e-8
+ lmin = 4.667e-8
+ voffcv = -0.125
+ wpemod = 1
+ tnoia = 0
+ lpe0 = 6.44e-8
+ lpeb = 0
+ ijthsfwd = 0.01
+ cigbacc = 0.245
+ peta0 = 5.969656900000001e-15
+ petab = -1.9628815e-15
+ minv = -0.33
+ lua1 = -1.9488641e-18
+ lub1 = 6.8003561e-26
+ wketa = -5.4843946e-8
+ luc1 = -2.115524e-18
+ tpbsw = 0.0025
+ ndep = 1e+18
+ tnoimod = 0
+ cjswd = 4.743e-11
+ lwlc = 0
+ cjsws = 4.743e-11
+ moin = 5.5538
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ nigc = 2.291
+ cigbinv = 0.006
+ ijthsrev = 0.01
+ tpbswg = 0.001
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ version = 4.5
+ tempmod = 0
+ ntox = 2.958
+ pcit = -1.96856065e-16
+ pclm = 1.3082183
+ scref = 1e-6
+ ptvoff = 9.8606268e-17
+ ppdiblc2 = 0
+ pigcd = 2.572
+ aigsd = 0.0063634291
+ waigsd = 1.9051377e-12
+ aigbacc = 0.012071
+ phin = 0.15
+ lvoff = -4.1725981e-9
+ diomod = 1
+ pkt1 = 1.3998109e-14
+ pkt2 = -4.0388508e-15
+ lvsat = -0.00230101408
+ lvth0 = -1.3915855e-9
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.6832999999999998e-10
+ pku0we = 0.0
+ cjswgs = 1.6832999999999998e-10
+ tvfbsdoff = 0.1
+ delta = 0.018814
+ aigbinv = 0.009974
+ laigc = -9.3796225e-12
+ rnoia = 0
+ rnoib = 0
+ rbdb = 50
+ pua1 = -1.9221227e-22
+ prwb = 0
+ pub1 = 2.2863324e-31
+ prwg = 0
+ puc1 = 2.3602641e-23
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ pkvth0we = 0.0
+ rbsb = 50
+ pvag = 2.1
+ mjswgd = 0.95
+ mjswgs = 0.95
+ rdsw = 200
+ pketa = 3.1809489e-15
+ ngate = 1.7e+20
+ ngcon = 1
+ tcjswg = 0.00128
+ wpclm = 1.8421624e-6
+ vfbsdoff = 0.01
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ poxedge = 1
+ paramchk = 1
+ rshg = 14.1
+ binunit = 2
+ ags = 2.6546816
+ cjd = 0.0012517799999999999
+ cit = 0.0014826020999999996
+ cjs = 0.0012517799999999999
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 4.0349e-9
+ fprout = 200
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ ijthdfwd = 0.01
+ la0 = -1.5436392e-7
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0.0035243403
+ kt1 = -0.063173267
+ kt2 = -0.094912467
+ lk2 = 3.878719299999999e-9
+ llc = 0
+ tvoff = 0.0053332949
+ lln = 1
+ lu0 = -7.3856189e-11
+ wtvoff = -1.4437583e-9
+ tnom = 25
+ mjd = 0.335
+ mjs = 0.335
+ lua = -3.3837758e-17
+ lub = -4.6371448999999997e-26
+ luc = -2.4014309e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = -3.174587e-14
+ toxe = 2.6300000000000002e-9
+ toxm = 2.67e-9
+ xjbvd = 1
+ xjbvs = 1
+ nsd = 1e+20
+ pbd = 0.75
+ pat = -5.2399134e-10
+ lk2we = 0.0
+ pbs = 0.75
+ pk2 = 5.1035691e-16
+ pu0 = -9.701894e-17
+ prt = 0
+ pua = -1.0296702e-22
+ pub = 1.544478e-31
+ puc = 2.16225e-23
+ pud = 0
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ rsh = 15.2
+ wtvfbsdoff = 0
+ tcj = 0.000832
+ ua1 = 5.6955479e-10
+ ub1 = -2.0140988e-18
+ uc1 = 2.5296559e-10
+ ijthdrev = 0.01
+ capmod = 2
+ tpb = 0.0016
+ wa0 = 3.9604044e-7
+ ute = -1
+ wat = 0.00058470362
+ ku0we = -0.0007
+ web = 6628.3
+ wec = -16935.0
+ wk2 = -9.6029938e-9
+ wku0we = 1.5e-11
+ wlc = 0
+ beta0 = 13.32
+ wln = 1
+ wu0 = 7.8023907e-10
+ xgl = -8.2e-9
+ xgw = 0
+ lpdiblc2 = 0
+ wua = 1.5228349e-15
+ wub = -2.8976024e-24
+ leta0 = -1.7797369000000001e-9
+ wuc = -4.6587973e-16
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ letab = 1.0403109e-8
+ ltvfbsdoff = 0
+ mobmod = 0
+ wags = 1.4000585e-6
+ ppclm = -9.0739811e-14
+ wcit = 3.33776483e-9
+ voff = -0.092743162
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ acde = 0.5
+ vsat = 124541.767
+ wint = 0
+ vth0 = -0.31382604000000003
+ wkt1 = -2.4366569e-7
+ wkt2 = 7.087942e-8
+ wmax = 8.9974e-6
+ aigc = 0.0066047781
+ wmin = 8.974e-7
+ njtsswg = 6.489
+ dmcgt = 0
+ lkvth0we = 3e-12
+ tcjsw = 9.34e-5
+ ptvfbsdoff = 0
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ wua1 = 3.9047481e-15
+ wub1 = -4.8164385e-24
+ wuc1 = -5.0052376e-16
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.00081573526
+ pdiblcb = 0
+ bigc = 0.0012521
+ acnqsmod = 0
+ wwlc = 0
+ bigsd = 0.0003327
+ cdsc = 0
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ wvoff = 1.0199556e-9
+ rbodymod = 0
+ cgbo = 0
+ cgdl = 3.2212350000000004e-11
+ cgdo = 2.8335740000000002e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.2212350000000004e-11
+ cgso = 2.8335740000000002e-11
+ cigc = 0.15259
+ wvsat = -0.0512507946
+ bigbacc = 0.0054401
+ wvth0 = 6.342809899999999e-8
+ waigc = 1.173226e-10
+ kvth0we = -0.00022
+ lintnoi = -5e-9
+ lketa = -6.6687589e-9
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ xpart = 1
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ wpdiblc2 = 1.6594883e-9
+ toxref = 3e-9
+ egidl = 0.001
+ k2we = 5e-5
+ dsub = 0.5
+ dtox = 3.91e-10
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ eta0 = 0.2041955
+ etab = -0.27743155
+ ltvoff = -2.3219338e-10
+ wkvth0we = 0.0
+ pvfbsdoff = 0
+ trnqsmod = 0
+ nfactor = 1
+ pvoff = -1.5168764999999998e-16
+ lku0we = 1.8e-11
+ cdscb = 0
+ cdscd = 0
+ epsrox = 3.9
+ pvsat = 2.72009693e-9
+ wk2we = 0.0
+ pvth0 = -2.6352739e-15
+ drout = 0.56
+ paigc = -5.5262052e-18
+ rdsmod = 0
+ igbmod = 1
+ rgatemod = 0
+ voffl = 0
+ tnjtsswg = 1
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ nigbacc = 10
+ weta0 = -1.3222145e-7
+ wetab = 5.0212024e-8
+ pbswgd = 0.8
+ pbswgs = 0.8
+ lpclm = -3.4164983e-8
+ a0 = 2.1782471
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = -44109.368
+ cf = 8.741900000000001e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.015698968
+ k3 = -2.5823
+ em = 20000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.0094255868
+ w0 = 0
+ igcmod = 1
+ ua = 3.7489785e-10
+ ub = 2.3165696e-18
+ uc = 4.9437493e-10
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 2.33e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ cgidl = 1
+ nigbinv = 2.171
+ pbswd = 0.9
+ pbsws = 0.9
+ )

.model pch_ff_16 pmos (
+ level = 54
+ wpdiblc2 = 1.6594883e-9
+ voffcv = -0.125
+ wpemod = 1
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ bigbacc = 0.0054401
+ tnom = 25
+ kvth0we = -0.00022
+ toxe = 2.6300000000000002e-9
+ toxm = 2.67e-9
+ bigsd = 0.0003327
+ lintnoi = -5e-9
+ wkvth0we = 0.0
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ wvoff = -9.7608128e-9
+ trnqsmod = 0
+ wvsat = 0.0192458405
+ tpbswg = 0.001
+ wvth0 = -1.04850767e-8
+ wags = 3.1454838e-6
+ waigc = -1.1150212e-11
+ wcit = -3.8116619e-9
+ voff = -0.099237323
+ acde = 0.5
+ lketa = 8.2510741e-9
+ ptvoff = -1.3565734e-16
+ xpart = 1
+ waigsd = 2.0479558e-12
+ vsat = 99605.54000000001
+ wint = 0
+ rgatemod = 0
+ vth0 = -0.35036593
+ wkt1 = 1.4686808e-7
+ wkt2 = -1.0928272e-8
+ tnjtsswg = 1
+ wmax = 8.9974e-6
+ aigc = 0.0065575398
+ wmin = 8.974e-7
+ diomod = 1
+ egidl = 0.001
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.6832999999999998e-10
+ pku0we = 0.0
+ cjswgs = 1.6832999999999998e-10
+ nfactor = 1
+ wua1 = -3.8771176e-15
+ wub1 = 5.8335837000000006e-24
+ wuc1 = 9.3089203e-17
+ bigc = 0.0012521
+ wwlc = 0
+ mjswgd = 0.95
+ mjswgs = 0.95
+ pvfbsdoff = 0
+ cdsc = 0
+ tcjswg = 0.00128
+ cgbo = 0
+ cgdl = 3.2212350000000004e-11
+ cgdo = 2.8335740000000002e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.2212350000000004e-11
+ cgso = 2.8335740000000002e-11
+ cigc = 0.15259
+ nigbacc = 10
+ pvoff = 3.7656999999999997e-16
+ cdscb = 0
+ cdscd = 0
+ pvsat = -7.342336900000001e-10
+ wk2we = 0.0
+ pvth0 = 9.864756e-16
+ drout = 0.56
+ paigc = 7.6896258e-19
+ nigbinv = 2.171
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ voffl = 0
+ dmdg = 0
+ fprout = 200
+ weta0 = -1.2697795500000002e-8
+ xrcrg1 = 12
+ xrcrg2 = 1
+ wetab = 3.974597e-8
+ wtvfbsdoff = 0
+ lpclm = -2.1829165e-8
+ k2we = 5e-5
+ dsub = 0.5
+ dtox = 3.91e-10
+ ijthsfwd = 0.01
+ wtvoff = 3.3371317e-9
+ cgidl = 1
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ fnoimod = 1
+ ltvfbsdoff = 0
+ eigbinv = 1.1
+ eta0 = 0.1123236
+ etab = -0.14869011
+ capmod = 2
+ pbswd = 0.9
+ pbsws = 0.9
+ ijthsrev = 0.01
+ wku0we = 1.5e-11
+ mobmod = 0
+ pdits = 0
+ cigsd = 0.013281
+ ptvfbsdoff = 0
+ cigbacc = 0.245
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ ppdiblc2 = 0
+ tnoimod = 0
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ laigsd = 7.7486946e-16
+ cigbinv = 0.006
+ tnoia = 0
+ peta0 = 1.1299919e-16
+ petab = -1.4500449e-15
+ wketa = 4.9202854e-8
+ version = 4.5
+ tpbsw = 0.0025
+ tempmod = 0
+ cjswd = 4.743e-11
+ pkvth0we = 0.0
+ cjsws = 4.743e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ agidl = 3.2166e-9
+ aigbacc = 0.012071
+ vfbsdoff = 0.01
+ keta = -0.24950779
+ lags = 9.4399385e-8
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 2.6904918e-10
+ aigbinv = 0.009974
+ kt1l = 0
+ paramchk = 1
+ scref = 1e-6
+ pigcd = 2.572
+ aigsd = 0.0063634133
+ toxref = 3e-9
+ lint = 0
+ lvoff = -3.8543842e-9
+ lkt1 = 6.7599286e-10
+ lkt2 = 4.9336152e-10
+ lmax = 4.667e-8
+ lmin = 3.6e-8
+ lpe0 = 6.44e-8
+ lvsat = -0.0010791554000000002
+ lpeb = 0
+ tvfbsdoff = 0.1
+ lvth0 = 3.98874294e-10
+ ijthdfwd = 0.01
+ delta = 0.018814
+ laigc = -7.0649434e-12
+ minv = -0.33
+ lua1 = -6.8231177e-17
+ lub1 = 7.9005491e-26
+ luc1 = 2.786749e-18
+ poxedge = 1
+ rnoia = 0
+ rnoib = 0
+ ndep = 1e+18
+ ltvoff = -9.8738127e-12
+ lwlc = 0
+ moin = 5.5538
+ binunit = 2
+ pketa = -1.9173443e-15
+ ngate = 1.7e+20
+ nigc = 2.291
+ ijthdrev = 0.01
+ ngcon = 1
+ wpclm = -3.2091624e-7
+ lpdiblc2 = 0
+ gbmin = 1e-12
+ lku0we = 1.8e-11
+ noff = 2.2684
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ epsrox = 3.9
+ ags = 0.72816353
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ cjd = 0.0012517799999999999
+ cit = -0.0038262097499999997
+ cjs = 0.0012517799999999999
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ pags = -8.5525843e-14
+ dlc = 4.0349e-9
+ k3b = 2.1176
+ rdsmod = 0
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ ntox = 2.958
+ pcit = 1.5346675e-16
+ pclm = 1.0564669
+ igbmod = 1
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ la0 = -3.7737017e-8
+ jsd = 1.5e-7
+ phin = 0.15
+ jss = 1.5e-7
+ lat = -0.0010396322
+ jtsswgd = 1.75e-7
+ kt1 = -0.34244081
+ kt2 = -0.083036557
+ lk2 = 3.6583258000000004e-9
+ jtsswgs = 1.75e-7
+ llc = 0
+ lln = 1
+ pbswgd = 0.8
+ pbswgs = 0.8
+ lu0 = 1.4117989e-10
+ mjd = 0.335
+ mjs = 0.335
+ lua = 2.9640356e-17
+ lub = 2.1940308999999997e-26
+ luc = -2.5002144e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ lkvth0we = 3e-12
+ njd = 1.02
+ njs = 1.02
+ pa0 = -1.5136929e-14
+ pkt1 = -5.1380439999999994e-15
+ pkt2 = -3.0273858e-17
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 1.2363197e-9
+ pbs = 0.75
+ pk2 = 4.883387e-16
+ igcmod = 1
+ pu0 = -4.5849539e-17
+ prt = 0
+ pua = 8.5912273e-23
+ pub = -1.7496088000000002e-31
+ puc = 8.2880171e-25
+ pud = 0
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 1.9222551e-9
+ ub1 = -2.2386283e-18
+ uc1 = 1.529192e-10
+ tvoff = 0.00079616085
+ tpb = 0.0016
+ wa0 = 5.7082474e-8
+ acnqsmod = 0
+ xjbvd = 1
+ ute = -1
+ wat = -0.035339966
+ xjbvs = 1
+ web = 6628.3
+ wec = -16935.0
+ rbdb = 50
+ wk2 = -9.1536426e-9
+ pua1 = 1.8909915e-22
+ prwb = 0
+ lk2we = 0.0
+ pub1 = -2.9321766999999996e-31
+ prwg = 0
+ puc1 = -5.4843946e-24
+ wlc = 0
+ wln = 1
+ wu0 = -2.6403442e-10
+ xgl = -8.2e-9
+ rbpb = 50
+ rbpd = 50
+ xgw = 0
+ rbps = 50
+ rbsb = 50
+ wua = -2.3318447e-15
+ pvag = 2.1
+ wub = 3.8250249e-24
+ wuc = -4.1518546e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ rdsw = 200
+ rbodymod = 0
+ paigsd = -6.9980875e-21
+ ku0we = -0.0007
+ beta0 = 13.32
+ njtsswg = 6.489
+ leta0 = 2.7219864e-9
+ letab = 4.094779e-9
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ ppclm = 1.5251044e-14
+ permod = 1
+ a0 = -0.20189383
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ ckappad = 0.6
+ at = 49032.992
+ cf = 8.741900000000001e-11
+ ckappas = 0.6
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.01120114
+ k3 = -2.5823
+ em = 20000000.0
+ dlcig = 2.5e-9
+ pdiblc1 = 0
+ pdiblc2 = 0.00081573526
+ ll = 0
+ lw = 0
+ bgidl = 1834800000.0
+ u0 = 0.005037095399999999
+ w0 = 0
+ pdiblcb = 0
+ ua = -9.2057386e-10
+ ub = 9.224525e-19
+ uc = 5.5311765e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 2.33e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ rshg = 14.1
+ )

.model pch_ff_17 pmos (
+ level = 54
+ tpbsw = 0.0025
+ aigbinv = 0.009974
+ eta0 = 0.191845
+ cjswd = 4.743e-11
+ cjsws = 4.743e-11
+ etab = -0.18516667
+ a0 = 2.6112
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ at = 72000
+ cf = 8.741900000000001e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.0045864754
+ k3 = -2.5823
+ em = 20000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.0094159667
+ w0 = 0
+ ua = 1.9119717e-10
+ ub = 1.0765761e-18
+ uc = -8.28048e-12
+ ud = 0
+ ijthdrev = 0.01
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 2.33e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ tpbswg = 0.001
+ lpdiblc2 = 0
+ ptvoff = 0
+ waigsd = 1.9350626e-12
+ scref = 1e-6
+ poxedge = 1
+ pigcd = 2.572
+ aigsd = 0.0063633642
+ diomod = 1
+ binunit = 2
+ lvoff = 0
+ pditsd = 0
+ lkvth0we = 3e-12
+ pditsl = 0
+ cjswgd = 1.6832999999999998e-10
+ pku0we = 0.0
+ cjswgs = 1.6832999999999998e-10
+ tvfbsdoff = 0.1
+ lvsat = -0.00028
+ lvth0 = 3e-10
+ delta = 0.018814
+ acnqsmod = 0
+ rnoia = 0
+ rnoib = 0
+ mjswgd = 0.95
+ mjswgs = 0.95
+ tcjswg = 0.00128
+ ngate = 1.7e+20
+ rbodymod = 0
+ ags = 0.98525249
+ ngcon = 1
+ wpclm = -5.08417e-8
+ cjd = 0.0012517799999999999
+ cit = 5e-6
+ cjs = 0.0012517799999999999
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ dlc = 1.0572421799999999e-8
+ k3b = 2.1176
+ dwb = 0
+ keta = -0.016063969
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ gbmin = 1e-12
+ wvfbsdoff = 0
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ lvfbsdoff = 0
+ wtvfbsdoff = 0
+ la0 = 0
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = -0.0008
+ lcit = -2e-11
+ kt1 = -0.18299632
+ lk2 = -4e-10
+ kt2 = -0.042133438
+ llc = 0
+ lln = 1
+ lu0 = -1.2e-11
+ mjd = 0.335
+ kt1l = 0
+ mjs = 0.335
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 0
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ ltvfbsdoff = 0
+ pk2 = 0
+ wpdiblc2 = -1.7580235e-10
+ fprout = 200
+ pu0 = 0
+ prt = 0
+ pud = 0
+ lint = 6.5375218e-9
+ xrcrg1 = 12
+ xrcrg2 = 1
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 1.45515e-9
+ ub1 = -1.5029257e-18
+ uc1 = -4.3667733e-11
+ lkt1 = 6e-10
+ lmax = 2.001e-5
+ tpb = 0.0016
+ wa0 = 2.308488e-7
+ lmin = 9.00077e-6
+ ute = -0.96728333
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 1.3953799e-9
+ njtsswg = 6.489
+ lpe0 = 6.44e-8
+ wlc = 0
+ wln = 1
+ wu0 = 2.7482e-12
+ xgl = -8.2e-9
+ lpeb = 0
+ xgw = 0
+ wua = -1.5682603e-16
+ wub = 3.5681818e-26
+ wuc = 4.8873989e-18
+ wud = 0
+ wtvoff = -7.2458121e-11
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ tvoff = 0.0025973351
+ minv = -0.33
+ xjbvd = 1
+ xjbvs = 1
+ ckappad = 0.6
+ ckappas = 0.6
+ lk2we = 0.0
+ ndep = 1e+18
+ pdiblc1 = 0
+ pdiblc2 = 0.0032290423
+ pdiblcb = 0
+ lwlc = 0
+ ptvfbsdoff = 0
+ capmod = 2
+ wkvth0we = 0.0
+ moin = 5.5538
+ wku0we = 1.5e-11
+ nigc = 2.291
+ trnqsmod = 0
+ mobmod = 0
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = 6e-10
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ bigbacc = 0.0054401
+ ppclm = 0
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ kvth0we = -0.00022
+ ntox = 2.958
+ pcit = 1e-18
+ pclm = 1.2411167
+ rgatemod = 0
+ lintnoi = -5e-9
+ tnjtsswg = 1
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ phin = 0.15
+ vtsswgs = 1.1
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ pkt1 = 5e-17
+ bigsd = 0.0003327
+ rbdb = 50
+ prwb = 0
+ prwg = 0
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ rdsw = 200
+ wvoff = 3.276885e-9
+ wvsat = -0.017628054
+ wvth0 = 3.7594256e-9
+ waigc = -7.2361068e-12
+ nfactor = 1
+ lketa = 0
+ rshg = 14.1
+ xpart = 1
+ toxref = 3e-9
+ egidl = 0.001
+ nigbacc = 10
+ ijthsfwd = 0.01
+ tnom = 25
+ ltvoff = 0
+ toxe = 2.6300000000000002e-9
+ toxm = 2.67e-9
+ pvfbsdoff = 0
+ nigbinv = 2.171
+ ijthsrev = 0.01
+ lku0we = 1.8e-11
+ pvoff = -2.5e-17
+ epsrox = 3.9
+ wags = -3.1938756e-8
+ cdscb = 0
+ cdscd = 0
+ pvsat = 0
+ wk2we = 0.0
+ rdsmod = 0
+ pvth0 = 1.5e-16
+ fnoimod = 1
+ drout = 0.56
+ voff = -0.10917042
+ igbmod = 1
+ acde = 0.5
+ eigbinv = 1.1
+ ppdiblc2 = 0
+ vsat = 129757.01
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ wint = 0
+ voffl = 0
+ vth0 = -0.35324647
+ wkt1 = 1.4804073e-9
+ wkt2 = -8.3218931e-9
+ pbswgd = 0.8
+ pbswgs = 0.8
+ wmax = 8.974e-7
+ aigc = 0.0068422292
+ wmin = 5.374e-7
+ weta0 = -2.404157e-8
+ wetab = 1.3741e-8
+ igcmod = 1
+ lpclm = 0
+ wua1 = -5.289391e-16
+ wub1 = 6.5622425e-25
+ wuc1 = 2.3227786e-17
+ cgidl = 1
+ bigc = 0.0012521
+ wute = -1.003093e-7
+ cigbacc = 0.245
+ wwlc = 0
+ pkvth0we = 0.0
+ cdsc = 0
+ tnoimod = 0
+ pbswd = 0.9
+ pbsws = 0.9
+ cgbo = 0
+ cgdl = 3.2212350000000004e-11
+ cgdo = 2.8335740000000002e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.2212350000000004e-11
+ cgso = 2.8335740000000002e-11
+ cigc = 0.15259
+ vfbsdoff = 0.01
+ cigbinv = 0.006
+ permod = 1
+ pdits = 0
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ paramchk = 1
+ version = 4.5
+ tempmod = 0
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ voffcv = -0.125
+ wpemod = 1
+ aigbacc = 0.012071
+ k2we = 5e-5
+ tnoia = 0
+ dsub = 0.5
+ dtox = 3.91e-10
+ ijthdfwd = 0.01
+ peta0 = 2e-17
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ wketa = -3.7023239e-9
+ )

.model pch_ff_18 pmos (
+ level = 54
+ waigc = -9.2878513e-12
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ nigbacc = 10
+ ptvoff = 6.0745993e-16
+ pags = -1.6587566e-14
+ waigsd = 1.93751e-12
+ lketa = -8.0782883e-8
+ ntox = 2.958
+ pcit = 1e-18
+ pclm = 1.2411167
+ xpart = 1
+ ppdiblc2 = 2.0750737e-15
+ diomod = 1
+ nigbinv = 2.171
+ phin = 0.15
+ egidl = 0.001
+ pditsd = 0
+ pditsl = 0
+ a0 = 2.6572474
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ cjswgd = 1.6832999999999998e-10
+ pku0we = 0.0
+ cjswgs = 1.6832999999999998e-10
+ at = 72000
+ cf = 8.741900000000001e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.0050849127
+ k3 = -2.5823
+ em = 20000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.009295758099999999
+ pkt1 = 7.5378862e-15
+ pkt2 = 7.624365e-15
+ w0 = 0
+ ua = 1.8022848e-10
+ ub = 1.0497212e-18
+ uc = -5.9216956e-12
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 2.33e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ mjswgd = 0.95
+ mjswgs = 0.95
+ rbdb = 50
+ pua1 = 3.0135942e-22
+ prwb = 0
+ pub1 = -6.7644414e-31
+ prwg = 0
+ fnoimod = 1
+ puc1 = -4.7294542e-23
+ pvfbsdoff = 0
+ wtvfbsdoff = 0
+ tcjswg = 0.00128
+ pkvth0we = 0.0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ eigbinv = 1.1
+ pute = 3.5290383e-14
+ rdsw = 200
+ ltvfbsdoff = 0
+ vfbsdoff = 0.01
+ pvoff = 7.7387382e-16
+ cdscb = 0
+ cdscd = 0
+ pvsat = 0
+ wk2we = 0.0
+ pvth0 = -1.0164923999999998e-15
+ drout = 0.56
+ paramchk = 1
+ paigc = 1.8445184e-17
+ rshg = 14.1
+ cigbacc = 0.245
+ fprout = 200
+ voffl = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ tnoimod = 0
+ ptvfbsdoff = 0
+ weta0 = -2.404157e-8
+ wetab = 1.3741e-8
+ lpclm = 0
+ wtvoff = -1.4002875e-10
+ cigbinv = 0.006
+ ijthdfwd = 0.01
+ cgidl = 1
+ tnom = 25
+ toxe = 2.6300000000000002e-9
+ toxm = 2.67e-9
+ capmod = 2
+ version = 4.5
+ wku0we = 1.5e-11
+ tempmod = 0
+ pbswd = 0.9
+ pbsws = 0.9
+ ijthdrev = 0.01
+ mobmod = 0
+ lpdiblc2 = 3.0626629e-9
+ aigbacc = 0.012071
+ wags = -3.0093643e-8
+ pdits = 0
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ voff = -0.10728654
+ acde = 0.5
+ vsat = 129757.01
+ aigbinv = 0.009974
+ wint = 0
+ vth0 = -0.35217796
+ laigsd = 5.7445099e-14
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ wkt1 = 6.4749443e-10
+ wkt2 = -9.1699871e-9
+ wmax = 8.974e-7
+ aigc = 0.0068507406
+ wmin = 5.374e-7
+ lkvth0we = 3e-12
+ tnoia = 0
+ peta0 = 2e-17
+ wua1 = -5.6246072e-16
+ wub1 = 7.3146831e-25
+ wuc1 = 2.8488581e-17
+ wketa = -8.2059163e-9
+ bigc = 0.0012521
+ wute = -1.0423482e-7
+ acnqsmod = 0
+ tpbsw = 0.0025
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ wwlc = 0
+ cjswd = 4.743e-11
+ cjsws = 4.743e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ poxedge = 1
+ cdsc = 0
+ rbodymod = 0
+ cgbo = 0
+ cgdl = 3.2212350000000004e-11
+ cgdo = 2.8335740000000002e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.2212350000000004e-11
+ cgso = 2.8335740000000002e-11
+ cigc = 0.15259
+ binunit = 2
+ toxref = 3e-9
+ scref = 1e-6
+ pigcd = 2.572
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ wpdiblc2 = -4.0662257e-10
+ aigsd = 0.0063633578
+ dmdg = 0
+ lvoff = -1.6936099e-8
+ tvfbsdoff = 0.1
+ k2we = 5e-5
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ lvsat = -0.00028
+ lvth0 = -9.3058678e-9
+ dsub = 0.5
+ dtox = 3.91e-10
+ delta = 0.018814
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ laigc = -7.651731e-11
+ ltvoff = -1.5996918e-9
+ ags = 0.95300429
+ rnoia = 0
+ rnoib = 0
+ cjd = 0.0012517799999999999
+ cit = 5e-6
+ cjs = 0.0012517799999999999
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 1.0572421799999999e-8
+ k3b = 2.1176
+ eta0 = 0.191845
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ etab = -0.18516667
+ dwj = 0
+ wkvth0we = 0.0
+ pketa = 4.0487295e-14
+ ngate = 1.7e+20
+ ngcon = 1
+ wpclm = -5.08417e-8
+ trnqsmod = 0
+ la0 = -4.1396638e-7
+ lku0we = 1.8e-11
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = -0.0008
+ kt1 = -0.17852273
+ kt2 = -0.039741464
+ lk2 = 4.0809517e-9
+ llc = 0
+ lln = 1
+ epsrox = 3.9
+ lu0 = 1.0686753e-9
+ mjd = 0.335
+ wvfbsdoff = 0
+ mjs = 0.335
+ lua = 9.8608496e-17
+ lub = 2.4142536e-25
+ luc = -2.1205472e-17
+ lud = 0
+ gbmin = 1e-12
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ lvfbsdoff = 0
+ njd = 1.02
+ njs = 1.02
+ pa0 = -1.9681175e-13
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ pk2 = -1.7465146e-15
+ njtsswg = 6.489
+ pu0 = -2.7146448e-18
+ rdsmod = 0
+ prt = 0
+ pua = -5.0852536e-23
+ pub = 3.3773548e-32
+ puc = 2.1258791e-23
+ pud = 0
+ igbmod = 1
+ xtsswgd = 0.32
+ rsh = 15.2
+ xtsswgs = 0.32
+ tcj = 0.000832
+ ua1 = 1.3709274e-9
+ ub1 = -1.4287011e-18
+ uc1 = -6.3574807e-11
+ tpb = 0.0016
+ wa0 = 2.527411e-7
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ ute = -0.97152091
+ ckappad = 0.6
+ ckappas = 0.6
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 1.5896529e-9
+ wlc = 0
+ rgatemod = 0
+ wln = 1
+ pdiblc1 = 0
+ pdiblc2 = 0.0028883679
+ wu0 = 3.0501627e-12
+ xgl = -8.2e-9
+ xgw = 0
+ pbswgd = 0.8
+ pdiblcb = 0
+ wua = -1.5116947e-16
+ pbswgs = 0.8
+ wub = 3.1925028e-26
+ wuc = 2.5226836e-18
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ tnjtsswg = 1
+ igcmod = 1
+ tvoff = 0.0027752763
+ bigbacc = 0.0054401
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ kvth0we = -0.00022
+ paigsd = -2.2002196e-20
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ ku0we = -0.0007
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ beta0 = 13.32
+ leta0 = 6e-10
+ keta = -0.0070781088
+ permod = 1
+ ppclm = 0
+ lags = 2.8991134e-7
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ dlcig = 2.5e-9
+ lcit = -2e-11
+ bgidl = 1834800000.0
+ kt1l = 0
+ voffcv = -0.125
+ wpemod = 1
+ lint = 6.5375218e-9
+ lkt1 = -3.9617527e-8
+ lkt2 = -2.1503841e-8
+ dmcgt = 0
+ lmax = 9.00077e-6
+ tcjsw = 9.34e-5
+ lmin = 9.0075e-7
+ lpe0 = 6.44e-8
+ lpeb = 0
+ ijthsfwd = 0.01
+ minv = -0.33
+ lua1 = 7.5716104e-16
+ lub1 = -6.6727951e-25
+ luc1 = 1.7896459e-16
+ nfactor = 1
+ bigsd = 0.0003327
+ ndep = 1e+18
+ lute = 3.8095772e-8
+ lwlc = 0
+ moin = 5.5538
+ wvoff = 3.1880225e-9
+ tpbswg = 0.001
+ ijthsrev = 0.01
+ nigc = 2.291
+ wvsat = -0.017628054
+ wvth0 = 3.8891800000000004e-9
+ noff = 2.2684
+ )

.model pch_ff_19 pmos (
+ level = 54
+ cjd = 0.0012517799999999999
+ cit = -8.7888889e-5
+ cjs = 0.0012517799999999999
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ lvsat = -0.00028
+ dlc = 1.0572421799999999e-8
+ k3b = 2.1176
+ lvth0 = 1.3342612e-10
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ ltvfbsdoff = 0
+ wua1 = -6.1430214e-16
+ wub1 = 1.1920544e-25
+ delta = 0.018814
+ wuc1 = -4.9561039e-17
+ laigc = -1.8208261e-11
+ mjswgd = 0.95
+ mjswgs = 0.95
+ njtsswg = 6.489
+ bigc = 0.0012521
+ wute = -1.2773023e-7
+ rnoia = 0
+ rnoib = 0
+ la0 = -9.6086602e-7
+ wwlc = 0
+ tcjswg = 0.00128
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = -0.0008
+ kt1 = -0.20738899
+ kt2 = -0.065812764
+ lk2 = -6.3080411e-10
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ llc = 0
+ lln = 1
+ lu0 = -1.5402407999999999e-9
+ mjd = 0.335
+ mjs = 0.335
+ lua = -3.205013e-16
+ lub = -3.7552526e-26
+ luc = 5.1848161e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 2.9499704e-13
+ pketa = -2.8529622e-14
+ ckappad = 0.6
+ cdsc = 0
+ ckappas = 0.6
+ ngate = 1.7e+20
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ pk2 = 8.8602334e-16
+ pdiblc1 = 0
+ pdiblc2 = -8.9657994e-6
+ cgbo = 0
+ cgdl = 3.2212350000000004e-11
+ cgdo = 2.8335740000000002e-11
+ xtid = 3
+ ngcon = 1
+ xtis = 3
+ pdiblcb = 0
+ pu0 = 4.0536683e-16
+ wpclm = -5.08417e-8
+ prt = 0
+ pua = 3.1718399e-23
+ pub = 9.4535502e-32
+ puc = -3.7711192e-23
+ pud = 0
+ cgsl = 3.2212350000000004e-11
+ cgso = 2.8335740000000002e-11
+ cigc = 0.15259
+ rsh = 15.2
+ wvfbsdoff = 0
+ tcj = 0.000832
+ ua1 = 2.985915e-9
+ ub1 = -2.7037422e-18
+ uc1 = 1.5248758e-10
+ lvfbsdoff = 0
+ gbmin = 1e-12
+ tpb = 0.0016
+ wa0 = -2.9985305e-7
+ jswgd = 3.69e-13
+ ptvfbsdoff = 0
+ jswgs = 3.69e-13
+ ute = -0.85901741
+ web = 6628.3
+ wec = -16935.0
+ wk2 = -1.3682549e-9
+ a0 = 3.2717414
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ wlc = 0
+ wln = 1
+ wu0 = -4.5546835e-10
+ at = 72000
+ cf = 8.741900000000001e-11
+ xgl = -8.2e-9
+ ef = 1.15
+ k1 = 0.30425
+ k2 = 0.00020919492
+ xgw = 0
+ k3 = -2.5823
+ em = 20000000.0
+ wua = -2.439458e-16
+ wub = -3.6346832e-26
+ wuc = 6.8781092e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ ll = 0
+ lw = 0
+ u0 = 0.012227123999999999
+ w0 = 0
+ ua = 6.5113837e-10
+ ub = 1.3631795e-18
+ uc = -8.8004429e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 2.33e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ bigbacc = 0.0054401
+ fprout = 200
+ xrcrg1 = 12
+ xrcrg2 = 1
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ kvth0we = -0.00022
+ lintnoi = -5e-9
+ wtvoff = 9.9743807e-10
+ bigbinv = 0.00149
+ k2we = 5e-5
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ dsub = 0.5
+ dtox = 3.91e-10
+ ijthsfwd = 0.01
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ tvoff = 0.00044287651
+ capmod = 2
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ wku0we = 1.5e-11
+ eta0 = 0.191845
+ etab = -0.18516667
+ mobmod = 0
+ ijthsrev = 0.01
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = 6e-10
+ ppclm = 0
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ nfactor = 1
+ laigsd = -3.6354984e-15
+ ppdiblc2 = -2.7249029e-15
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ nigbacc = 10
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ bigsd = 0.0003327
+ pkvth0we = 0.0
+ wvoff = 1.2743983e-8
+ nigbinv = 2.171
+ wvsat = -0.017628054
+ vfbsdoff = 0.01
+ wvth0 = 1.9692885800000002e-9
+ keta = -0.13767457
+ waigc = 2.7297355e-11
+ lags = 8.1183869e-8
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 6.2671111e-11
+ toxref = 3e-9
+ paramchk = 1
+ lketa = 3.5447968e-8
+ kt1l = 0
+ xpart = 1
+ fnoimod = 1
+ eigbinv = 1.1
+ lint = 6.5375218e-9
+ egidl = 0.001
+ lkt1 = -1.3926561e-8
+ lkt2 = 1.6996159e-9
+ lmax = 9.0075e-7
+ lmin = 4.5075e-7
+ lpe0 = 6.44e-8
+ lpeb = 0
+ ijthdfwd = 0.01
+ ltvoff = 4.7614406e-10
+ minv = -0.33
+ lua1 = -6.8017788e-16
+ lub1 = 4.6750711e-25
+ luc1 = -1.3330934e-17
+ pvfbsdoff = 0
+ ndep = 1e+18
+ lute = -6.2032341e-8
+ lwlc = 0
+ moin = 5.5538
+ cigbacc = 0.245
+ ijthdrev = 0.01
+ nigc = 2.291
+ lku0we = 1.8e-11
+ epsrox = 3.9
+ tnoimod = 0
+ lpdiblc2 = 5.64129e-9
+ pvoff = -7.7309313e-15
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ rdsmod = 0
+ cdscb = 0
+ cdscd = 0
+ cigbinv = 0.006
+ igbmod = 1
+ pvsat = 0
+ wk2we = 0.0
+ pvth0 = 6.9221102e-16
+ drout = 0.56
+ pags = 2.5130854e-13
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ paigc = -1.411565e-17
+ ntox = 2.958
+ pcit = 1e-18
+ pclm = 1.2411167
+ pbswgd = 0.8
+ pbswgs = 0.8
+ voffl = 0
+ version = 4.5
+ igcmod = 1
+ phin = 0.15
+ tempmod = 0
+ weta0 = -2.404157e-8
+ wetab = 1.3741e-8
+ lkvth0we = 3e-12
+ lpclm = 0
+ pkt1 = -4.5911548e-15
+ pkt2 = -3.0623252e-15
+ aigbacc = 0.012071
+ cgidl = 1
+ acnqsmod = 0
+ rbdb = 50
+ pua1 = 3.4749829e-22
+ prwb = 0
+ pub1 = -1.3153018e-31
+ prwg = 0
+ puc1 = 2.216962e-23
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ paigsd = 1.9849821e-21
+ rbsb = 50
+ pvag = 2.1
+ pute = 5.6201301e-14
+ rdsw = 200
+ rbodymod = 0
+ pbswd = 0.9
+ pbsws = 0.9
+ aigbinv = 0.009974
+ permod = 1
+ pdits = 0
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ rshg = 14.1
+ voffcv = -0.125
+ wpemod = 1
+ wpdiblc2 = 4.9866096e-9
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ poxedge = 1
+ tnoia = 0
+ binunit = 2
+ peta0 = 2e-17
+ wketa = 6.9341182e-8
+ tnom = 25
+ tpbsw = 0.0025
+ toxe = 2.6300000000000002e-9
+ toxm = 2.67e-9
+ cjswd = 4.743e-11
+ cjsws = 4.743e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ wkvth0we = 0.0
+ agidl = 3.2166e-9
+ tpbswg = 0.001
+ trnqsmod = 0
+ wags = -3.311005e-7
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ ptvoff = -4.0488554e-16
+ waigsd = 1.9105581e-12
+ voff = -0.13228318
+ acde = 0.5
+ scref = 1e-6
+ diomod = 1
+ vsat = 129757.01
+ pigcd = 2.572
+ rgatemod = 0
+ wint = 0
+ aigsd = 0.0063634264
+ vth0 = -0.36278391
+ tnjtsswg = 1
+ wkt1 = 1.4275631e-8
+ wkt2 = 2.8375299e-9
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.6832999999999998e-10
+ pku0we = 0.0
+ wmax = 8.974e-7
+ wtvfbsdoff = 0
+ cjswgs = 1.6832999999999998e-10
+ aigc = 0.0067852248
+ lvoff = 5.3109112e-9
+ wmin = 5.374e-7
+ ags = 1.1875295
+ tvfbsdoff = 0.1
+ )

.model pch_ff_20 pmos (
+ level = 54
+ cjd = 0.0012517799999999999
+ cit = -0.00041212495
+ cjs = 0.0012517799999999999
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ lvsat = -0.00028
+ dlc = 1.38228675e-8
+ k3b = 2.1176
+ lvth0 = 6.8054743e-9
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ ltvfbsdoff = 0
+ wua1 = 2.4012676e-16
+ wub1 = -6.2487918e-26
+ delta = 0.018814
+ wuc1 = -3.9943707e-17
+ laigc = -2.2400472e-11
+ mjswgd = 0.95
+ mjswgs = 0.95
+ njtsswg = 6.489
+ bigc = 0.0012521
+ rnoia = 0
+ rnoib = 0
+ la0 = -7.2511148e-8
+ wwlc = 0
+ tcjswg = 0.00128
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = -0.0008
+ kt1 = -0.20886849
+ kt2 = -0.049681978
+ lk2 = 8.117425999999999e-10
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ llc = -1.18e-13
+ lln = 0.7
+ lu0 = -4.929571499999999e-10
+ mjd = 0.335
+ mjs = 0.335
+ lua = -5.9775833e-17
+ lub = -8.2990392e-26
+ luc = -8.4878869e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = -2.0868237e-13
+ pketa = -1.8963071e-15
+ ckappad = 0.6
+ cdsc = 0
+ ckappas = 0.6
+ ngate = 1.7e+20
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ pk2 = -3.6576402e-16
+ pdiblc1 = 0
+ pdiblc2 = 0.01788848
+ cgbo = 0
+ cgdl = 3.2212350000000004e-11
+ cgdo = 2.8335740000000002e-11
+ xtid = 3
+ ngcon = 1
+ xtis = 3
+ pdiblcb = 0
+ pu0 = -2.2283222e-17
+ wpclm = -5.08417e-8
+ prt = 0
+ pua = -3.7414239e-23
+ pub = 6.4271496e-32
+ puc = -3.5764571e-25
+ pud = 0
+ cgsl = 3.2212350000000004e-11
+ cgso = 2.8335740000000002e-11
+ cigc = 0.15259
+ rsh = 15.2
+ wvfbsdoff = 0
+ tcj = 0.000832
+ ua1 = 1.3271195e-9
+ ub1 = -1.4620758e-18
+ uc1 = 1.6497662e-10
+ lvfbsdoff = 0
+ gbmin = 1e-12
+ tpb = 0.0016
+ wa0 = 8.4487289e-7
+ jswgd = 3.69e-13
+ ptvfbsdoff = 0
+ jswgs = 3.69e-13
+ ute = -1
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 1.4767164e-9
+ a0 = 1.2527531
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ wlc = 0
+ wln = 1
+ wu0 = 5.1646359e-10
+ at = 72000
+ cf = 8.741900000000001e-11
+ xgl = -8.2e-9
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.0030693202
+ xgw = 0
+ k3 = -2.5823
+ em = 20000000.0
+ wua = -8.6826164e-17
+ wub = 3.2435001e-26
+ wuc = -1.6113333e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ ll = -1.18e-13
+ lw = 0
+ u0 = 0.009846934
+ w0 = 0
+ ua = 5.8580479e-11
+ ub = 1.4664474e-18
+ uc = 4.9122952e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 2.33e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ bigbacc = 0.0054401
+ fprout = 200
+ xrcrg1 = 12
+ xrcrg2 = 1
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ kvth0we = -0.00022
+ lintnoi = -5e-9
+ wtvoff = -3.604609e-11
+ bigbinv = 0.00149
+ k2we = 5e-5
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ dsub = 0.5
+ dtox = 3.91e-10
+ ijthsfwd = 0.01
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ tvoff = 0.0020688013
+ capmod = 2
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ wku0we = 1.5e-11
+ eta0 = 0.191845
+ etab = -0.18516667
+ mobmod = 0
+ ijthsrev = 0.01
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = 6e-10
+ ppclm = 0
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ nfactor = 1
+ ppdiblc2 = 1.0915468e-15
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ nigbacc = 10
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ bigsd = 0.0003327
+ pkvth0we = 0.0
+ wvoff = -5.0330429e-9
+ nigbinv = 2.171
+ wvsat = -0.017628054
+ vfbsdoff = 0.01
+ wvth0 = 7.1926608000000005e-9
+ keta = -0.023696099
+ waigc = -1.2459534e-12
+ lags = 6.5053339e-7
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 2.0533497999999998e-10
+ toxref = 3e-9
+ paramchk = 1
+ lketa = -1.4702559e-8
+ kt1l = 0
+ xpart = 1
+ fnoimod = 1
+ eigbinv = 1.1
+ lint = 9.7879675e-9
+ egidl = 0.001
+ lkt1 = -1.3275578999999999e-8
+ lkt2 = -5.3979298e-9
+ lmax = 4.5075e-7
+ lmin = 2.1744e-7
+ lpe0 = 6.44e-8
+ lpeb = 0
+ ijthdfwd = 0.01
+ ltvoff = -2.3926284e-10
+ minv = -0.33
+ lua1 = 4.9692128e-17
+ lub1 = -7.8826099e-26
+ luc1 = -1.8826114e-17
+ pvfbsdoff = 0
+ ndep = 1e+18
+ lwlc = 0
+ moin = 5.5538
+ cigbacc = 0.245
+ ijthdrev = 0.01
+ nigc = 2.291
+ lku0we = 1.8e-11
+ epsrox = 3.9
+ tnoimod = 0
+ lpdiblc2 = -2.233586e-9
+ pvoff = 9.096021e-17
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ rdsmod = 0
+ cdscb = 0
+ cdscd = 0
+ cigbinv = 0.006
+ igbmod = 1
+ pvsat = 0
+ wk2we = 0.0
+ pvth0 = -1.6060727e-15
+ drout = 0.56
+ pags = 1.3163813e-13
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ paigc = -1.5565945e-18
+ ntox = 2.958
+ pcit = -1.9500563999999998e-17
+ pclm = 1.2411167
+ pbswgd = 0.8
+ pbswgs = 0.8
+ voffl = 0
+ version = 4.5
+ igcmod = 1
+ phin = 0.15
+ tempmod = 0
+ weta0 = -2.404157e-8
+ wetab = 1.3741e-8
+ lkvth0we = 3e-12
+ lpclm = 0
+ pkt1 = 1.2073276e-15
+ pkt2 = 6.9635068e-17
+ aigbacc = 0.012071
+ cgidl = 1
+ acnqsmod = 0
+ rbdb = 50
+ pua1 = -2.8450432e-23
+ prwb = 0
+ pub1 = -5.1585101e-32
+ prwg = 0
+ puc1 = 1.7937993e-23
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ rdsw = 200
+ rbodymod = 0
+ pbswd = 0.9
+ pbsws = 0.9
+ aigbinv = 0.009974
+ permod = 1
+ pdits = 0
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ rshg = 14.1
+ voffcv = -0.125
+ wpemod = 1
+ wpdiblc2 = -3.6871397e-9
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ poxedge = 1
+ tnoia = 0
+ binunit = 2
+ peta0 = 2e-17
+ wketa = 8.8109206e-9
+ tnom = 25
+ tpbsw = 0.0025
+ toxe = 2.6300000000000002e-9
+ toxm = 2.67e-9
+ cjswd = 4.743e-11
+ cjsws = 4.743e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ wkvth0we = 0.0
+ agidl = 3.2166e-9
+ tpbswg = 0.001
+ trnqsmod = 0
+ wags = -5.9122303e-8
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ ptvoff = 4.9847489e-17
+ wcit = 4.6592191e-11
+ waigsd = 1.9150694e-12
+ voff = -0.10909205
+ acde = 0.5
+ scref = 1e-6
+ diomod = 1
+ vsat = 129757.01
+ pigcd = 2.572
+ rgatemod = 0
+ wint = 0
+ aigsd = 0.0063634182
+ vth0 = -0.37794766
+ tnjtsswg = 1
+ wkt1 = 1.0972613e-9
+ wkt2 = -4.2805615e-9
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.6832999999999998e-10
+ pku0we = 0.0
+ wmax = 8.974e-7
+ wtvfbsdoff = 0
+ cjswgs = 1.6832999999999998e-10
+ aigc = 0.0067947526
+ lvoff = -4.893186e-9
+ wmin = 5.374e-7
+ ags = -0.10644665
+ tvfbsdoff = 0.1
+ )

.model pch_ff_21 pmos (
+ level = 54
+ rbodymod = 0
+ version = 4.5
+ tempmod = 0
+ keta = -0.074839654
+ pvoff = 2.547289e-16
+ cdscb = 0
+ cdscd = 0
+ lags = 2.5597727e-7
+ pvsat = 0
+ aigbacc = 0.012071
+ wk2we = 0.0
+ pvth0 = 5.771049399999999e-16
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ drout = 0.56
+ fprout = 200
+ lcit = 1.2712816e-10
+ kt1l = 0
+ paigc = 3.3660127e-18
+ xrcrg1 = 12
+ xrcrg2 = 1
+ voffl = 0
+ wpdiblc2 = 2.1803424e-9
+ lint = 9.7879675e-9
+ weta0 = -2.404157e-8
+ wtvoff = -4.3702924e-10
+ aigbinv = 0.009974
+ wetab = 1.3741e-8
+ lkt1 = -5.564347099999999e-9
+ lkt2 = -3.8990903e-9
+ lmax = 2.1744e-7
+ lpclm = 5.4900145e-8
+ lmin = 9.167e-8
+ lpe0 = 6.44e-8
+ lpeb = 0
+ cgidl = 1
+ minv = -0.33
+ capmod = 2
+ lua1 = -2.9544713e-16
+ lub1 = 3.7855773e-25
+ luc1 = 4.6029572e-17
+ wku0we = 1.5e-11
+ a0 = 0.98313605
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ ndep = 1e+18
+ at = 41320.114
+ cf = 8.741900000000001e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.016096302
+ k3 = -2.5823
+ em = 20000000.0
+ ll = -1.18e-13
+ lwlc = 0
+ lw = 0
+ u0 = 0.008396993
+ mobmod = 0
+ w0 = 0
+ wkvth0we = 0.0
+ ua = 2.7312462e-10
+ ub = 6.1180894e-19
+ uc = 6.0007215e-11
+ ud = 0
+ moin = 5.5538
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 2.33e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ pbswd = 0.9
+ pbsws = 0.9
+ nigc = 2.291
+ trnqsmod = 0
+ poxedge = 1
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ binunit = 2
+ pdits = 0
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ pags = -1.3976359e-13
+ ntox = 2.958
+ pcit = -3.5385120000000004e-17
+ pclm = 0.98092641
+ rgatemod = 0
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ tnjtsswg = 1
+ phin = 0.15
+ pkt1 = 1.592035e-15
+ pkt2 = 2.2793112e-15
+ tnoia = 0
+ peta0 = 2e-17
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ wketa = -2.2984762e-8
+ tpbsw = 0.0025
+ rbdb = 50
+ pua1 = 7.9342593e-23
+ prwb = 0
+ pub1 = -9.194958e-32
+ prwg = 0
+ puc1 = -2.9723056e-23
+ cjswd = 4.743e-11
+ cjsws = 4.743e-11
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ mjswd = 0.01
+ rbsb = 50
+ pvag = 2.1
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ rdsw = 200
+ toxref = 3e-9
+ njtsswg = 6.489
+ ags = 1.7634876
+ scref = 1e-6
+ rshg = 14.1
+ cjd = 0.0012517799999999999
+ cit = -4.1476524e-5
+ cjs = 0.0012517799999999999
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ xtsswgd = 0.32
+ pigcd = 2.572
+ xtsswgs = 0.32
+ dlc = 1.38228675e-8
+ aigsd = 0.0063634182
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ tvfbsdoff = 0.1
+ ckappad = 0.6
+ ckappas = 0.6
+ lvoff = -2.4249846e-9
+ pdiblc1 = 0
+ pdiblc2 = 0.011594472
+ pdiblcb = 0
+ la0 = -1.5621959e-8
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0.0056734559999999995
+ lvsat = -0.00028
+ kt1 = -0.24541461
+ kt2 = -0.056785482
+ lk2 = 3.5604228000000005e-9
+ llc = -1.18e-13
+ lvth0 = 4.2839767000000005e-9
+ lln = 0.7
+ ltvoff = -2.3342435e-10
+ lu0 = -1.8701951e-10
+ mjd = 0.335
+ mjs = 0.335
+ lua = -1.0504465e-16
+ ijthsfwd = 0.01
+ lub = 9.7338322e-26
+ luc = -1.0784466e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ delta = 0.018814
+ pa0 = -2.5809676e-14
+ nsd = 1e+20
+ laigc = -2.5435198e-11
+ pbd = 0.75
+ pat = -8.1994638e-9
+ pbs = 0.75
+ pk2 = 1.2451684e-16
+ tnom = 25
+ pu0 = -7.9199366e-18
+ prt = 0
+ pua = 5.00917e-23
+ pub = -8.1076857e-32
+ puc = 8.6464743e-24
+ pud = 0
+ rnoia = 0
+ rnoib = 0
+ toxe = 2.6300000000000002e-9
+ toxm = 2.67e-9
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 2.9628506e-9
+ ub1 = -3.6297717e-18
+ uc1 = -1.423963e-10
+ bigbacc = 0.0054401
+ tpb = 0.0016
+ wa0 = -2.1822352e-8
+ pketa = 4.8125819e-15
+ ute = -1
+ wat = 0.038860018
+ ngate = 1.7e+20
+ web = 6628.3
+ wec = -16935.0
+ lku0we = 1.8e-11
+ wk2 = -8.468563e-10
+ wlc = 0
+ wln = 1
+ ijthsrev = 0.01
+ wu0 = 4.4839114e-10
+ xgl = -8.2e-9
+ ngcon = 1
+ xgw = 0
+ epsrox = 3.9
+ wua = -5.0154626e-16
+ wub = 7.2128975e-25
+ wuc = -5.8786887e-17
+ wud = 0
+ wpclm = 1.8489068e-7
+ wwc = 0
+ kvth0we = -0.00022
+ wwl = 0
+ wwn = 1
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ gbmin = 1e-12
+ lintnoi = -5e-9
+ rdsmod = 0
+ jswgd = 3.69e-13
+ bigbinv = 0.00149
+ jswgs = 3.69e-13
+ wags = 1.2271418e-6
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ igbmod = 1
+ wcit = 1.2187445e-10
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ voff = -0.12078969
+ acde = 0.5
+ pbswgd = 0.8
+ pbswgs = 0.8
+ ppdiblc2 = -1.4649193e-16
+ vsat = 129757.01
+ wint = 0
+ vth0 = -0.36599742999999996
+ igcmod = 1
+ wkt1 = -7.259963e-10
+ wkt2 = -1.475296e-8
+ wmax = 8.974e-7
+ aigc = 0.0068091352
+ wmin = 5.374e-7
+ wua1 = -2.7074066e-16
+ wub1 = 1.2881293e-25
+ wuc1 = 1.8593804e-16
+ tvoff = 0.0020411307
+ bigc = 0.0012521
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ wwlc = 0
+ pkvth0we = 0.0
+ nfactor = 1
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.2212350000000004e-11
+ cgdo = 2.8335740000000002e-11
+ xtid = 3
+ xtis = 3
+ permod = 1
+ ku0we = -0.0007
+ cgsl = 3.2212350000000004e-11
+ cgso = 2.8335740000000002e-11
+ cigc = 0.15259
+ beta0 = 13.32
+ vfbsdoff = 0.01
+ leta0 = 6e-10
+ ppclm = -4.9739531e-14
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ nigbacc = 10
+ paramchk = 1
+ voffcv = -0.125
+ wpemod = 1
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ nigbinv = 2.171
+ k2we = 5e-5
+ dsub = 0.5
+ ijthdfwd = 0.01
+ dtox = 3.91e-10
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ bigsd = 0.0003327
+ eta0 = 0.191845
+ tpbswg = 0.001
+ etab = -0.18516667
+ wvoff = -5.8091978e-9
+ fnoimod = 1
+ ijthdrev = 0.01
+ eigbinv = 1.1
+ wvsat = -0.017628054
+ wvth0 = -3.1541528999999996e-9
+ lpdiblc2 = -9.0555048e-10
+ wtvfbsdoff = 0
+ ptvoff = 1.3445493e-16
+ waigc = -2.4575845e-11
+ waigsd = 1.9150694e-12
+ ltvfbsdoff = 0
+ lketa = -3.9112692e-9
+ diomod = 1
+ xpart = 1
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.6832999999999998e-10
+ pku0we = 0.0
+ cjswgs = 1.6832999999999998e-10
+ cigbacc = 0.245
+ egidl = 0.001
+ lkvth0we = 3e-12
+ tnoimod = 0
+ mjswgd = 0.95
+ mjswgs = 0.95
+ cigbinv = 0.006
+ tcjswg = 0.00128
+ pvfbsdoff = 0
+ ptvfbsdoff = 0
+ acnqsmod = 0
+ )

.model pch_ff_22 pmos (
+ level = 54
+ xrcrg1 = 12
+ xrcrg2 = 1
+ paramchk = 1
+ rshg = 14.1
+ nfactor = 1
+ wtvoff = 2.0697628e-9
+ ijthdfwd = 0.01
+ capmod = 2
+ tvoff = -0.0031746364
+ tnom = 25
+ wku0we = 1.5e-11
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ toxe = 2.6300000000000002e-9
+ toxm = 2.67e-9
+ mobmod = 0
+ nigbacc = 10
+ ijthdrev = 0.01
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = -9.451894999999999e-9
+ lpdiblc2 = 0
+ letab = 1.4778454e-8
+ nigbinv = 2.171
+ wags = -2.597049e-7
+ ppclm = 2.5985382e-14
+ wcit = 2.8161348999999996e-10
+ dlcig = 2.5e-9
+ laigsd = 2.2969081e-18
+ bgidl = 1834800000.0
+ voff = -0.11952627
+ acde = 0.5
+ vsat = 238954.38
+ wint = 0
+ vth0 = -0.3217255
+ a0 = 2.9368155
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ wkt1 = -1.289882e-8
+ wkt2 = 2.7006409e-8
+ at = 192293.99
+ cf = 8.741900000000001e-11
+ wmax = 8.974e-7
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.02088367
+ k3 = -2.5823
+ em = 20000000.0
+ fnoimod = 1
+ aigc = 0.0066428307
+ wmin = 5.374e-7
+ ll = 0
+ lw = 0
+ u0 = 0.0079935417
+ dmcgt = 0
+ w0 = 0
+ ua = -1.5734149e-9
+ ub = 3.8310868000000005e-18
+ uc = -1.3540772e-10
+ ud = 0
+ tcjsw = 9.34e-5
+ wl = 0
+ lkvth0we = 3e-12
+ wr = 1
+ xj = 1.1e-7
+ eigbinv = 1.1
+ xl = 2.33e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ wua1 = 6.2697239e-16
+ wub1 = -9.8389336e-25
+ wuc1 = -5.3295995e-16
+ bigc = 0.0012521
+ acnqsmod = 0
+ bigsd = 0.0003327
+ wwlc = 0
+ wvoff = -3.6240027e-9
+ cdsc = 0
+ rbodymod = 0
+ cgbo = 0
+ cgdl = 3.2212350000000004e-11
+ cgdo = 2.8335740000000002e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.2212350000000004e-11
+ cgso = 2.8335740000000002e-11
+ cigbacc = 0.245
+ wvsat = -0.079474309
+ cigc = 0.15259
+ wvth0 = 5.378886400000001e-9
+ waigc = 3.8715701e-11
+ tnoimod = 0
+ toxref = 3e-9
+ lketa = 1.7736502e-8
+ cigbinv = 0.006
+ xpart = 1
+ wpdiblc2 = 6.2191766e-10
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ egidl = 0.001
+ version = 4.5
+ ltvoff = 2.5685776e-10
+ k2we = 5e-5
+ tempmod = 0
+ dsub = 0.5
+ dtox = 3.91e-10
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ pvfbsdoff = 0
+ aigbacc = 0.012071
+ eta0 = 0.29878005
+ etab = -0.34238426
+ wkvth0we = 0.0
+ lku0we = 1.8e-11
+ epsrox = 3.9
+ trnqsmod = 0
+ rdsmod = 0
+ aigbinv = 0.009974
+ pvoff = 4.9320558e-17
+ igbmod = 1
+ cdscb = 0
+ cdscd = 0
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ pvsat = 5.8135478e-9
+ wk2we = 0.0
+ pvth0 = -2.2500085000000005e-16
+ drout = 0.56
+ pbswgd = 0.8
+ pbswgs = 0.8
+ paigc = -2.5833927e-18
+ igcmod = 1
+ voffl = 0
+ rgatemod = 0
+ tnjtsswg = 1
+ weta0 = -7.0040749e-8
+ wetab = 2.4810139e-8
+ lpclm = -5.2812564e-8
+ poxedge = 1
+ cgidl = 1
+ binunit = 2
+ paigsd = -2.080997e-24
+ pbswd = 0.9
+ pbsws = 0.9
+ permod = 1
+ keta = -0.30513509
+ pdits = 0
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ jtsswgd = 1.75e-7
+ lcit = 1.3805001e-10
+ jtsswgs = 1.75e-7
+ voffcv = -0.125
+ wpemod = 1
+ kt1l = 0
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ lint = 0
+ lkt1 = -3.5189262e-9
+ lkt2 = 3.753071e-9
+ lmax = 9.167e-8
+ lmin = 5.567e-8
+ tnoia = 0
+ lpe0 = 6.44e-8
+ lpeb = 0
+ ijthsfwd = 0.01
+ peta0 = 4.3439229e-15
+ petab = -1.0404991e-15
+ wketa = 1.6222018e-7
+ minv = -0.33
+ wtvfbsdoff = 0
+ lua1 = 1.1693458e-16
+ lub1 = -2.0580342e-25
+ luc1 = -5.5456179e-17
+ tpbsw = 0.0025
+ tpbswg = 0.001
+ ndep = 1e+18
+ cjswd = 4.743e-11
+ njtsswg = 6.489
+ cjsws = 4.743e-11
+ mjswd = 0.01
+ lwlc = 0
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ moin = 5.5538
+ ltvfbsdoff = 0
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ ijthsrev = 0.01
+ nigc = 2.291
+ ckappad = 0.6
+ ckappas = 0.6
+ ags = 4.48665
+ pdiblc1 = 0
+ pdiblc2 = 0.0019609567
+ ptvoff = -1.0118352e-16
+ pdiblcb = 0
+ cjd = 0.0012517799999999999
+ cit = -0.00015766541000000002
+ waigsd = 1.9150916e-12
+ cjs = 0.0012517799999999999
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ noff = 2.2684
+ bvs = 8.2
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ dlc = 4.0349e-9
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ diomod = 1
+ scref = 1e-6
+ ntox = 2.958
+ pcit = -5.04005987e-17
+ pclm = 2.1268063
+ la0 = -1.9926782e-7
+ pditsd = 0
+ pditsl = 0
+ ppdiblc2 = 0
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = -0.0085180887
+ cjswgd = 1.6832999999999998e-10
+ pku0we = 0.0
+ pigcd = 2.572
+ kt1 = -0.26717441
+ cjswgs = 1.6832999999999998e-10
+ kt2 = -0.13819145
+ lk2 = 4.0104354e-9
+ aigsd = 0.0063634181
+ bigbacc = 0.0054401
+ llc = 0
+ ptvfbsdoff = 0
+ lln = 1
+ lu0 = -1.4909508e-10
+ mjd = 0.335
+ mjs = 0.335
+ lua = 6.8530064e-17
+ lub = -2.0527384e-25
+ luc = 7.5845372e-18
+ lud = 0
+ tvfbsdoff = 0.1
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 2.4118768e-14
+ phin = 0.15
+ lvoff = -2.5437461e-9
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 2.0972465e-9
+ pbs = 0.75
+ pk2 = 2.0570947e-16
+ pu0 = 1.8416833e-16
+ kvth0we = -0.00022
+ prt = 0
+ pua = -1.7823119e-23
+ pub = 1.5394810000000002e-31
+ puc = -7.4643321e-24
+ pud = 0
+ pkt1 = 2.7362803e-15
+ pkt2 = -1.6460695e-15
+ lvsat = -0.010544556
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = -1.4241889e-9
+ ub1 = 2.5868363e-18
+ mjswgd = 0.95
+ lvth0 = 1.224120899999999e-10
+ uc1 = 9.3723935e-10
+ mjswgs = 0.95
+ lintnoi = -5e-9
+ tpb = 0.0016
+ wa0 = -5.5297601e-7
+ delta = 0.018814
+ bigbinv = 0.00149
+ ute = -1
+ vtsswgd = 1.1
+ wat = -0.070679454
+ laigc = -9.8025804e-12
+ vtsswgs = 1.1
+ tcjswg = 0.00128
+ web = 6628.3
+ wec = -16935.0
+ wk2 = -1.7106076e-9
+ wlc = 0
+ wln = 1
+ wu0 = -1.5951011e-9
+ xgl = -8.2e-9
+ xgw = 0
+ wua = 2.2095182e-16
+ wub = -1.7789759e-24
+ wuc = 1.1260467e-16
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ rnoia = 0
+ rnoib = 0
+ rbdb = 50
+ pua1 = -5.0424332e-24
+ prwb = 0
+ pub1 = 1.2644812e-32
+ prwg = 0
+ puc1 = 3.7853356e-23
+ pkvth0we = 0.0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ pketa = -1.2596682e-14
+ ngate = 1.7e+20
+ rdsw = 200
+ ngcon = 1
+ wvfbsdoff = 0
+ wpclm = -6.2069351e-7
+ lvfbsdoff = 0
+ vfbsdoff = 0.01
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ fprout = 200
+ )

.model pch_ff_23 pmos (
+ level = 54
+ ijthsfwd = 0.01
+ dtox = 3.91e-10
+ cgidl = 1
+ wku0we = 1.5e-11
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ mobmod = 0
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ eta0 = 7.956713e-6
+ etab = -0.26192508
+ pbswd = 0.9
+ pbsws = 0.9
+ ijthsrev = 0.01
+ pdits = 0
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ ppdiblc2 = 0
+ njtsswg = 6.489
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ tnoia = 0
+ ckappad = 0.6
+ ckappas = 0.6
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ pdiblc1 = 0
+ pdiblc2 = 0.0019609567
+ pdiblcb = 0
+ peta0 = -2.7792439000000003e-15
+ petab = -1.6989745e-15
+ wketa = -4.2902456e-7
+ tpbsw = 0.0025
+ cjswd = 4.743e-11
+ cjsws = 4.743e-11
+ pkvth0we = 0.0
+ ags = 4.48665
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ cjd = 0.0012517799999999999
+ cit = 0.006990067
+ cjs = 0.0012517799999999999
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 4.0349e-9
+ bigbacc = 0.0054401
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ vfbsdoff = 0.01
+ a0 = 5.6551822
+ a1 = 0
+ a2 = 1
+ keta = 0.46798148
+ b0 = 0
+ b1 = 0
+ kvth0we = -0.00022
+ at = -40561.437
+ cf = 8.741900000000001e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.018874979
+ k3 = -2.5823
+ em = 20000000.0
+ la0 = -3.569331e-7
+ toxref = 3e-9
+ ll = 0
+ jsd = 1.5e-7
+ lw = 0
+ jss = 1.5e-7
+ lat = 0.0049875263
+ u0 = 0.0069984758999999995
+ w0 = 0
+ kt1 = -0.46532049
+ kt2 = 0.0072316444
+ lk2 = 3.8939313e-9
+ ua = 5.3944309e-9
+ ub = -9.4033093e-18
+ uc = 1.0922891e-10
+ ud = 0
+ llc = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 2.33e-9
+ ww = 0
+ lln = 1
+ xw = 8.600000000000001e-9
+ lu0 = -9.138127e-11
+ mjd = 0.335
+ lintnoi = -5e-9
+ mjs = 0.335
+ lua = -3.3560499e-16
+ lub = 5.623213400000001e-25
+ luc = -6.604387e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ bigbinv = 0.00149
+ njs = 1.02
+ pa0 = 1.517818e-13
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ nsd = 1e+20
+ lcit = -2.7651581e-10
+ pbd = 0.75
+ pat = -1.8496379e-9
+ pbs = 0.75
+ pk2 = 4.9657487e-16
+ paramchk = 1
+ pu0 = -8.1141216e-17
+ scref = 1e-6
+ kt1l = 0
+ prt = 0
+ pua = 1.7043409e-22
+ pub = -3.9702784e-31
+ puc = 5.8491101e-24
+ pud = 0
+ pigcd = 2.572
+ rsh = 15.2
+ aigsd = 0.0063634182
+ tcj = 0.000832
+ ua1 = 9.464156e-9
+ tvfbsdoff = 0.1
+ ub1 = -1.352433e-17
+ uc1 = -1.5339544e-9
+ tpb = 0.0016
+ wa0 = -2.7540628e-6
+ lint = 0
+ ute = -1
+ wat = -0.002629722
+ lvoff = -5.520199e-9
+ web = 6628.3
+ wec = -16935.0
+ wk2 = -6.7255282e-9
+ wlc = 0
+ wln = 1
+ lkt1 = 7.9735466e-9
+ lkt2 = -4.6814687e-9
+ wu0 = 2.9792015e-9
+ xgl = -8.2e-9
+ xgw = 0
+ ltvoff = -2.6406105e-10
+ wua = -3.0248621e-15
+ wub = 7.7206094e-24
+ wuc = -1.1693744e-16
+ wud = 0
+ lmax = 5.567e-8
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ lmin = 4.667e-8
+ lvsat = 0.008578704199999999
+ lpe0 = 6.44e-8
+ lvth0 = -5.4835768e-9
+ lpeb = 0
+ ijthdfwd = 0.01
+ delta = 0.018814
+ laigc = -1.6050622e-11
+ minv = -0.33
+ lua1 = -5.1458943e-16
+ lub1 = 7.2864421e-25
+ luc1 = 8.7873061e-17
+ rnoia = 0
+ rnoib = 0
+ ndep = 1e+18
+ lku0we = 1.8e-11
+ lwlc = 0
+ epsrox = 3.9
+ moin = 5.5538
+ pketa = 2.1695512e-14
+ ngate = 1.7e+20
+ wvfbsdoff = 0
+ ijthdrev = 0.01
+ lvfbsdoff = 0
+ ngcon = 1
+ nigc = 2.291
+ wpclm = -1.0386396e-6
+ nfactor = 1
+ rdsmod = 0
+ igbmod = 1
+ lpdiblc2 = 0
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ noff = 2.2684
+ pscbe1 = 926400000.0
+ noia = 2.86e+42
+ pscbe2 = 1e-20
+ noib = 2.5e+24
+ noic = 31000000000.0
+ pbswgd = 0.8
+ pbswgs = 0.8
+ igcmod = 1
+ ntox = 2.958
+ pcit = 6.1746976e-17
+ pclm = 4.4879115
+ nigbacc = 10
+ phin = 0.15
+ lkvth0we = 3e-12
+ pkt1 = -5.0112736e-15
+ pkt2 = 1.1767646e-15
+ nigbinv = 2.171
+ tvoff = 0.0058067224
+ acnqsmod = 0
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ rbdb = 50
+ pua1 = 2.7224008e-22
+ prwb = 0
+ pub1 = -3.6990718e-31
+ prwg = 0
+ puc1 = -5.7927018e-23
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ permod = 1
+ rbodymod = 0
+ rdsw = 200
+ ku0we = -0.0007
+ beta0 = 13.32
+ fnoimod = 1
+ leta0 = 7.8768866e-9
+ letab = 1.0111821e-8
+ eigbinv = 1.1
+ ppclm = 5.0226256e-14
+ voffcv = -0.125
+ wpemod = 1
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ rshg = 14.1
+ wtvfbsdoff = 0
+ wpdiblc2 = 6.2191766e-10
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ ltvfbsdoff = 0
+ cigbacc = 0.245
+ tnoimod = 0
+ tnom = 25
+ tpbswg = 0.001
+ bigsd = 0.0003327
+ toxe = 2.6300000000000002e-9
+ toxm = 2.67e-9
+ cigbinv = 0.006
+ wkvth0we = 0.0
+ wvoff = -2.1208799e-8
+ trnqsmod = 0
+ wvsat = 0.14380976
+ ptvoff = 1.2747838e-16
+ ptvfbsdoff = 0
+ wvth0 = -1.6984308000000004e-8
+ waigsd = 1.9150557e-12
+ version = 4.5
+ waigc = -1.4751759e-11
+ wags = -2.597049e-7
+ tempmod = 0
+ wcit = -1.6519588900000002e-9
+ diomod = 1
+ voff = -0.068208113
+ lketa = -2.7104259e-8
+ acde = 0.5
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.6832999999999998e-10
+ pku0we = 0.0
+ cjswgs = 1.6832999999999998e-10
+ aigbacc = 0.012071
+ xpart = 1
+ rgatemod = 0
+ vsat = -90756.867
+ wint = 0
+ vth0 = -0.2250704
+ tnjtsswg = 1
+ wkt1 = 1.206797e-7
+ wkt2 = -2.1663145e-8
+ egidl = 0.001
+ wmax = 8.974e-7
+ aigc = 0.0067505556
+ wmin = 5.374e-7
+ mjswgd = 0.95
+ mjswgs = 0.95
+ aigbinv = 0.009974
+ tcjswg = 0.00128
+ pvfbsdoff = 0
+ wua1 = -4.1537606e-15
+ wub1 = 5.6118307e-24
+ wuc1 = 1.1184258e-15
+ bigc = 0.0012521
+ wwlc = 0
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.2212350000000004e-11
+ cgdo = 2.8335740000000002e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.2212350000000004e-11
+ cgso = 2.8335740000000002e-11
+ cigc = 0.15259
+ pvoff = 1.0692388e-15
+ poxedge = 1
+ cdscb = 0
+ cdscd = 0
+ fprout = 200
+ pvsat = -7.136935500000001e-9
+ wk2we = 0.0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ pvth0 = 1.0720697000000001e-15
+ drout = 0.56
+ binunit = 2
+ paigc = 5.1772001e-19
+ voffl = 0
+ dmcg = 3.1e-8
+ wtvoff = -1.8726837e-9
+ dmci = 3.1e-8
+ dmdg = 0
+ weta0 = 5.2772471e-8
+ wetab = 3.6163164e-8
+ lpclm = -1.8975667e-7
+ k2we = 5e-5
+ capmod = 2
+ dsub = 0.5
+ )

.model pch_ff_24 pmos (
+ level = 54
+ beta0 = 13.32
+ leta0 = 3.24810824e-9
+ letab = 2.8639817e-9
+ cigbacc = 0.245
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ ppclm = -6.983762e-15
+ laigsd = -1.7489044e-14
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ tnoimod = 0
+ ntox = 2.958
+ pcit = -1.0672974999999996e-16
+ pclm = 0.55996802
+ rgatemod = 0
+ cigbinv = 0.006
+ tnjtsswg = 1
+ phin = 0.15
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ pkt1 = 4.802240900000001e-15
+ pkt2 = -6.3201272e-16
+ version = 4.5
+ tempmod = 0
+ bigsd = 0.0003327
+ rbdb = 50
+ pua1 = -2.7866327e-22
+ prwb = 0
+ pub1 = 3.5479518e-31
+ prwg = 0
+ puc1 = 2.5974765e-23
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ aigbacc = 0.012071
+ wvoff = -2.6959456e-8
+ rdsw = 200
+ wvsat = -0.002403996999999998
+ wvth0 = -2.4175461e-9
+ toxref = 3e-9
+ waigc = -9.7737582e-11
+ aigbinv = 0.009974
+ lketa = 1.4220453e-8
+ rshg = 14.1
+ xpart = 1
+ egidl = 0.001
+ ltvoff = -2.5344658e-10
+ pvfbsdoff = 0
+ ijthsfwd = 0.01
+ poxedge = 1
+ a0 = -2.5402778
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ tnom = 25
+ at = 196072.83
+ cf = 8.741900000000001e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.022656115
+ k3 = -2.5823
+ em = 20000000.0
+ lku0we = 1.8e-11
+ ll = 0
+ lw = 0
+ u0 = 0.0011078574
+ w0 = 0
+ toxe = 2.6300000000000002e-9
+ toxm = 2.67e-9
+ ua = -6.0379704e-9
+ ub = 7.7384779e-18
+ uc = -2.2784413e-10
+ ud = 0
+ binunit = 2
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 2.33e-9
+ ww = 0
+ epsrox = 3.9
+ xw = 8.600000000000001e-9
+ ijthsrev = 0.01
+ rdsmod = 0
+ igbmod = 1
+ pvoff = 1.351021e-15
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ wags = -2.597049e-7
+ cdscb = 0
+ cdscd = 0
+ pbswgd = 0.8
+ pbswgs = 0.8
+ pvsat = 2.7544300000000016e-11
+ wcit = 1.7862688999999995e-9
+ wk2we = 0.0
+ pvth0 = 3.5829728e-16
+ drout = 0.56
+ igcmod = 1
+ voff = -0.080254273
+ paigc = 4.5840253e-18
+ acde = 0.5
+ ppdiblc2 = 0
+ voffl = 0
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ vsat = 123501.56
+ wint = 0
+ vth0 = -0.35927062000000004
+ wkt1 = -7.959638e-8
+ wkt2 = 1.5250678e-8
+ wmax = 8.974e-7
+ weta0 = 3.474872000000002e-9
+ aigc = 0.0066531108
+ wetab = 8.325777e-9
+ wmin = 5.374e-7
+ lpclm = 2.7125638e-9
+ cgidl = 1
+ paigsd = 9.5490179e-21
+ wua1 = 7.089165e-15
+ wub1 = -9.1780167e-24
+ wuc1 = -5.9385548e-16
+ bigc = 0.0012521
+ wwlc = 0
+ pkvth0we = 0.0
+ permod = 1
+ cdsc = 0
+ pbswd = 0.9
+ pbsws = 0.9
+ njtsswg = 6.489
+ cgbo = 0
+ cgdl = 3.2212350000000004e-11
+ cgdo = 2.8335740000000002e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.2212350000000004e-11
+ cgso = 2.8335740000000002e-11
+ wtvfbsdoff = 0
+ cigc = 0.15259
+ vfbsdoff = 0.01
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ ckappad = 0.6
+ ckappas = 0.6
+ pdits = 0
+ voffcv = -0.125
+ wpemod = 1
+ pdiblc1 = 0
+ pdiblc2 = 0.0019609567
+ cigsd = 0.013281
+ ltvfbsdoff = 0
+ pdiblcb = 0
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ paramchk = 1
+ pk2we = 0.0
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ bigbacc = 0.0054401
+ tnoia = 0
+ k2we = 5e-5
+ ags = 4.48665
+ ijthdfwd = 0.01
+ dsub = 0.5
+ dtox = 3.91e-10
+ kvth0we = -0.00022
+ peta0 = -3.636599599999999e-16
+ ptvfbsdoff = 0
+ petab = -3.349425e-16
+ cjd = 0.0012517799999999999
+ cit = -0.010005025
+ cjs = 0.0012517799999999999
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dvt0 = 3.48
+ tpbswg = 0.001
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ wketa = 1.6324308e-7
+ dlc = 4.0349e-9
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ tpbsw = 0.0025
+ dwg = 0
+ lintnoi = -5e-9
+ dwj = 0
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ cjswd = 4.743e-11
+ cjsws = 4.743e-11
+ mjswd = 0.01
+ eta0 = 0.09447294
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ etab = -0.11400999
+ la0 = 4.4644444e-8
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = -0.0066075577
+ kt1 = -0.09248022000000003
+ kt2 = -0.11193164
+ lk2 = 4.0792069999999995e-9
+ ijthdrev = 0.01
+ llc = 0
+ lln = 1
+ lu0 = 1.9725904e-10
+ mjd = 0.335
+ ptvoff = 8.5019581e-17
+ mjs = 0.335
+ lua = 2.2458267e-16
+ lub = -2.7762652e-25
+ luc = 9.9121919e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = -8.9774533e-14
+ waigsd = 1.7201778e-12
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 6.2808619e-9
+ pbs = 0.75
+ lpdiblc2 = 0
+ pk2 = 1.0702031e-16
+ pu0 = -9.6657248e-17
+ prt = 0
+ pua = -9.0705467e-23
+ pub = 9.644662000000001e-32
+ puc = -1.0416838e-23
+ pud = 0
+ diomod = 1
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = -1.018181e-8
+ ub1 = 1.4330462e-17
+ uc1 = 9.111363e-10
+ tpb = 0.0016
+ wa0 = 2.1756583e-6
+ ute = -1
+ wat = -0.16855824
+ pditsd = 0
+ web = 6628.3
+ wec = -16935.0
+ pditsl = 0
+ wk2 = 1.2245648e-9
+ cjswgd = 1.6832999999999998e-10
+ pku0we = 0.0
+ cjswgs = 1.6832999999999998e-10
+ wlc = 0
+ wln = 1
+ wu0 = 3.2958552e-9
+ xgl = -8.2e-9
+ xgw = 0
+ scref = 1e-6
+ wua = 2.3045166e-15
+ wub = -2.3502966999999998e-24
+ wuc = 2.150207e-16
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ tvfbsdoff = 0.1
+ pigcd = 2.572
+ aigsd = 0.0063637751
+ lvoff = -4.9299372e-9
+ mjswgd = 0.95
+ mjswgs = 0.95
+ lkvth0we = 3e-12
+ nfactor = 1
+ lvsat = -0.00191997372
+ tcjswg = 0.00128
+ lvth0 = 1.09222701e-9
+ delta = 0.018814
+ laigc = -1.1275829e-11
+ acnqsmod = 0
+ rnoia = 0
+ rnoib = 0
+ wvfbsdoff = 0
+ pketa = -7.3256019e-15
+ ngate = 1.7e+20
+ lvfbsdoff = 0
+ rbodymod = 0
+ nigbacc = 10
+ ngcon = 1
+ wpclm = 1.2891178e-7
+ gbmin = 1e-12
+ keta = -0.37538
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ fprout = 200
+ xrcrg1 = 12
+ xrcrg2 = 1
+ nigbinv = 2.171
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 5.5623864e-10
+ kt1l = 0
+ wtvoff = -1.0061777e-9
+ wpdiblc2 = 6.2191766e-10
+ lint = 0
+ lkt1 = -1.0295661e-8
+ lkt2 = 1.1575324e-9
+ lmax = 4.667e-8
+ lmin = 3.6e-8
+ capmod = 2
+ fnoimod = 1
+ lpe0 = 6.44e-8
+ lpeb = 0
+ wku0we = 1.5e-11
+ eigbinv = 1.1
+ tvoff = 0.0055901005
+ mobmod = 0
+ minv = -0.33
+ lua1 = 4.4806289e-16
+ lub1 = -6.3624048e-25
+ luc1 = -3.1936385e-17
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ ndep = 1e+18
+ wkvth0we = 0.0
+ lwlc = 0
+ moin = 5.5538
+ nigc = 2.291
+ trnqsmod = 0
+ ku0we = -0.0007
+ )

.model pch_ff_25 pmos (
+ level = 54
+ wint = 0
+ ags = 0.93810347
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ vth0 = -0.34798248
+ wkt1 = -1.5318394e-9
+ wkt2 = 2.21858e-9
+ cjd = 0.0012517799999999999
+ cit = 5e-6
+ cjs = 0.0012517799999999999
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ wmax = 5.374e-7
+ bvs = 8.2
+ aigc = 0.0068215676
+ wmin = 2.674e-7
+ dlc = 1.0572421799999999e-8
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ k3b = 2.1176
+ lkvth0we = 3e-12
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ tnoia = 0
+ peta0 = 2e-17
+ la0 = 0
+ wua1 = 1.6452204e-16
+ wub1 = -6.9710259e-26
+ wuc1 = 2.1709154e-17
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = -0.0008
+ wketa = 2.2687563e-8
+ kt1 = -0.17747938
+ lk2 = -4e-10
+ kt2 = -0.061438333
+ llc = 0
+ lln = 1
+ lu0 = -1.2e-11
+ tpbsw = 0.0025
+ acnqsmod = 0
+ mjd = 0.335
+ bigc = 0.0012521
+ mjs = 0.335
+ wute = 3.2371733e-8
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ wwlc = 0
+ pa0 = 0
+ cjswd = 4.743e-11
+ nsd = 1e+20
+ cjsws = 4.743e-11
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ pk2 = 0
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ pu0 = 0
+ prt = 0
+ pud = 0
+ rbodymod = 0
+ cdsc = 0
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 1.8507467e-10
+ ub1 = -1.7337534e-19
+ uc1 = -4.0886356e-11
+ cgbo = 0
+ cgdl = 3.2212350000000004e-11
+ cgdo = 2.8335740000000002e-11
+ xtid = 3
+ xtis = 3
+ tpb = 0.0016
+ wa0 = -1.5013787e-7
+ cgsl = 3.2212350000000004e-11
+ cgso = 2.8335740000000002e-11
+ cigc = 0.15259
+ ute = -1.2102889
+ toxref = 3e-9
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 4.440518e-10
+ wlc = 0
+ wln = 1
+ wu0 = 3.7953067e-11
+ xgl = -8.2e-9
+ xgw = 0
+ nfactor = 1
+ wua = -1.5196107e-16
+ wub = 9.0507286e-26
+ wuc = 5.3799588e-18
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ scref = 1e-6
+ tvfbsdoff = 0.1
+ pigcd = 2.572
+ aigsd = 0.0063632886
+ wpdiblc2 = -7.7579138e-11
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ ltvoff = 0
+ lvoff = 0
+ nigbacc = 10
+ lvsat = -0.00028
+ k2we = 5e-5
+ lvth0 = 3e-10
+ dsub = 0.5
+ dtox = 3.91e-10
+ delta = 0.018814
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ lku0we = 1.8e-11
+ rnoia = 0
+ rnoib = 0
+ epsrox = 3.9
+ nigbinv = 2.171
+ eta0 = 0.17962267
+ wvfbsdoff = 0
+ wkvth0we = 0.0
+ etab = -0.19577778
+ lvfbsdoff = 0
+ ngate = 1.7e+20
+ rdsmod = 0
+ ngcon = 1
+ igbmod = 1
+ wpclm = -1.1447315e-8
+ trnqsmod = 0
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ pbswgd = 0.8
+ pbswgs = 0.8
+ fnoimod = 1
+ eigbinv = 1.1
+ igcmod = 1
+ a0 = 3.3089778
+ a1 = 0
+ a2 = 1
+ rgatemod = 0
+ b0 = 0
+ b1 = 0
+ at = 72000
+ cf = 8.741900000000001e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.0028441163
+ k3 = -2.5823
+ em = 20000000.0
+ tnjtsswg = 1
+ ll = 0
+ lw = 0
+ u0 = 0.0093514889
+ w0 = 0
+ ua = 1.8228697e-10
+ ub = 9.7616315e-19
+ uc = -9.1826044e-12
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 2.33e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ wtvfbsdoff = 0
+ cigbacc = 0.245
+ tvoff = 0.0026578776
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ permod = 1
+ ltvfbsdoff = 0
+ tnoimod = 0
+ cigbinv = 0.006
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = 6e-10
+ keta = -0.064397096
+ voffcv = -0.125
+ wpemod = 1
+ ppclm = 0
+ version = 4.5
+ dlcig = 2.5e-9
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ bgidl = 1834800000.0
+ lcit = -2e-11
+ tempmod = 0
+ ptvfbsdoff = 0
+ kt1l = 0
+ aigbacc = 0.012071
+ lint = 6.5375218e-9
+ dmcgt = 0
+ lkt1 = 6e-10
+ tcjsw = 9.34e-5
+ lmax = 2.001e-5
+ lmin = 9.00077e-6
+ lpe0 = 6.44e-8
+ lpeb = 0
+ ijthsfwd = 0.01
+ tpbswg = 0.001
+ minv = -0.33
+ aigbinv = 0.009974
+ bigsd = 0.0003327
+ ndep = 1e+18
+ lwlc = 0
+ moin = 5.5538
+ wvoff = 2.5521431e-9
+ ptvoff = 0
+ ijthsrev = 0.01
+ nigc = 2.291
+ waigsd = 1.9763167e-12
+ wvsat = 0.0034765009
+ wvth0 = 8.852853000000001e-10
+ diomod = 1
+ waigc = 4.045116e-12
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.6832999999999998e-10
+ pku0we = 0.0
+ cjswgs = 1.6832999999999998e-10
+ poxedge = 1
+ lketa = 0
+ ntox = 2.958
+ xpart = 1
+ pcit = 1e-18
+ pclm = 1.1689658
+ ppdiblc2 = 0
+ binunit = 2
+ egidl = 0.001
+ mjswgd = 0.95
+ mjswgs = 0.95
+ phin = 0.15
+ tcjswg = 0.00128
+ pkt1 = 5e-17
+ pvfbsdoff = 0
+ rbdb = 50
+ prwb = 0
+ prwg = 0
+ pkvth0we = 0.0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ jtsswgd = 1.75e-7
+ rdsw = 200
+ jtsswgs = 1.75e-7
+ vfbsdoff = 0.01
+ fprout = 200
+ pvoff = -2.5e-17
+ xrcrg1 = 12
+ xrcrg2 = 1
+ cdscb = 0
+ cdscd = 0
+ pvsat = 0
+ wk2we = 0.0
+ pvth0 = 1.5e-16
+ drout = 0.56
+ paramchk = 1
+ wtvoff = -1.0551434e-10
+ rshg = 14.1
+ voffl = 0
+ weta0 = -1.7368176e-8
+ wetab = 1.9534667e-8
+ njtsswg = 6.489
+ capmod = 2
+ lpclm = 0
+ wku0we = 1.5e-11
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ ijthdfwd = 0.01
+ cgidl = 1
+ mobmod = 0
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.0030491463
+ tnom = 25
+ pdiblcb = 0
+ toxe = 2.6300000000000002e-9
+ toxm = 2.67e-9
+ pbswd = 0.9
+ pbsws = 0.9
+ ijthdrev = 0.01
+ lpdiblc2 = 0
+ bigbacc = 0.0054401
+ wags = -6.1953916e-9
+ pdits = 0
+ cigsd = 0.013281
+ kvth0we = -0.00022
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ voff = -0.10784306
+ acde = 0.5
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ vsat = 91103.982
+ pk2we = 0.0
+ )

.model pch_ff_26 pmos (
+ level = 54
+ bigsd = 0.0003327
+ poxedge = 1
+ pkvth0we = 0.0
+ wvoff = 2.9007224e-9
+ binunit = 2
+ toxref = 3e-9
+ wvsat = 0.0034765009
+ wvth0 = 8.237108000000001e-10
+ vfbsdoff = 0.01
+ keta = -0.06875265
+ waigc = 4.3476029e-12
+ lags = 1.0877241e-7
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = -2e-11
+ lketa = 3.9156432e-8
+ paramchk = 1
+ kt1l = 0
+ xpart = 1
+ ltvoff = -4.4286369e-10
+ egidl = 0.001
+ lint = 6.5375218e-9
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ lkt1 = -3.4253729e-8
+ lkt2 = -1.4641311e-8
+ lmax = 9.00077e-6
+ pvfbsdoff = 0
+ lmin = 9.0075e-7
+ lpe0 = 6.44e-8
+ ijthdfwd = 0.01
+ lpeb = 0
+ lku0we = 1.8e-11
+ minv = -0.33
+ epsrox = 3.9
+ lua1 = 1.4818924e-15
+ lub1 = -2.0711788e-24
+ luc1 = 2.2491171e-16
+ ndep = 1e+18
+ lute = 1.330224e-7
+ rdsmod = 0
+ lwlc = 0
+ moin = 5.5538
+ igbmod = 1
+ ijthdrev = 0.01
+ nigc = 2.291
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ lpdiblc2 = 8.2033961e-9
+ njtsswg = 6.489
+ pbswgd = 0.8
+ pvoff = -3.1587282e-15
+ pbswgs = 0.8
+ noff = 2.2684
+ cdscb = 0
+ cdscd = 0
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ igcmod = 1
+ pvsat = 0
+ wk2we = 0.0
+ pvth0 = 7.0355474e-16
+ drout = 0.56
+ ckappad = 0.6
+ ckappas = 0.6
+ pags = 8.2314292e-14
+ wtvfbsdoff = 0
+ pdiblc1 = 0
+ pdiblc2 = 0.002136644
+ paigc = -2.7193569e-18
+ pdiblcb = 0
+ ntox = 2.958
+ pcit = 1e-18
+ pclm = 1.1689658
+ voffl = 0
+ ltvfbsdoff = 0
+ weta0 = -1.7368176e-8
+ phin = 0.15
+ wetab = 1.9534667e-8
+ lkvth0we = 3e-12
+ lpclm = 0
+ paigsd = -4.5957918e-20
+ pkt1 = 4.609252599999999e-15
+ pkt2 = 3.8774237e-15
+ bigbacc = 0.0054401
+ cgidl = 1
+ permod = 1
+ acnqsmod = 0
+ kvth0we = -0.00022
+ rbdb = 50
+ pua1 = -9.4343892e-23
+ prwb = 0
+ pub1 = 9.0084871e-32
+ prwg = 0
+ puc1 = -7.238167e-23
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ lintnoi = -5e-9
+ pute = -1.6539558e-14
+ bigbinv = 0.00149
+ rbodymod = 0
+ pbswd = 0.9
+ pbsws = 0.9
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ rdsw = 200
+ ptvfbsdoff = 0
+ a0 = 3.4253346
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 72000
+ cf = 8.741900000000001e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.0024652651
+ k3 = -2.5823
+ em = 20000000.0
+ ll = 0
+ voffcv = -0.125
+ lw = 0
+ wpemod = 1
+ u0 = 0.009235427499999999
+ w0 = 0
+ ua = 1.8429003e-10
+ ub = 9.3982253e-19
+ uc = -1.1498405e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 2.33e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ pdits = 0
+ cigsd = 0.013281
+ ags = 0.9260042
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ cjd = 0.0012517799999999999
+ cit = 5e-6
+ cjs = 0.0012517799999999999
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 1.0572421799999999e-8
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ rshg = 14.1
+ wpdiblc2 = 3.818702e-12
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ la0 = -1.0460478e-6
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = -0.0008
+ kt1 = -0.17360244
+ kt2 = -0.059809712
+ lk2 = -3.8058721e-9
+ llc = 0
+ lln = 1
+ lu0 = 1.0313917e-9
+ mjd = 0.335
+ mjs = 0.335
+ lua = -1.8007487e-17
+ lub = 3.2670219e-25
+ luc = 2.0819042e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ tnoia = 0
+ njd = 1.02
+ njs = 1.02
+ pa0 = 1.483047e-13
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ tpbswg = 0.001
+ pk2 = 2.5596912e-15
+ pu0 = 1.7642195e-17
+ nfactor = 1
+ peta0 = 2e-17
+ prt = 0
+ pua = 1.2819791e-23
+ pub = -1.2787603e-32
+ puc = -1.6865938e-24
+ pud = 0
+ wketa = 2.5468383e-8
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 2.0236805e-11
+ ub1 = 5.7011626e-20
+ uc1 = -6.5904343e-11
+ tnom = 25
+ tpbsw = 0.0025
+ tpb = 0.0016
+ wa0 = -1.666345e-7
+ toxe = 2.6300000000000002e-9
+ toxm = 2.67e-9
+ ute = -1.2250856
+ cjswd = 4.743e-11
+ cjsws = 4.743e-11
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 1.5932531e-10
+ mjswd = 0.01
+ wlc = 0
+ mjsws = 0.01
+ wln = 1
+ agidl = 3.2166e-9
+ wu0 = 3.5990642e-11
+ wkvth0we = 0.0
+ xgl = -8.2e-9
+ xgw = 0
+ wua = -1.5338707e-16
+ wub = 9.1929712e-26
+ wuc = 5.5675666e-18
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ ptvoff = -2.4168192e-17
+ waigsd = 1.9814288e-12
+ trnqsmod = 0
+ nigbacc = 10
+ diomod = 1
+ wags = -1.5351598e-8
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.6832999999999998e-10
+ pku0we = 0.0
+ cjswgs = 1.6832999999999998e-10
+ tvfbsdoff = 0.1
+ voff = -0.10676035
+ scref = 1e-6
+ acde = 0.5
+ nigbinv = 2.171
+ pigcd = 2.572
+ rgatemod = 0
+ aigsd = 0.0063632773
+ vsat = 91103.982
+ wint = 0
+ vth0 = -0.34656355000000005
+ tnjtsswg = 1
+ mjswgd = 0.95
+ mjswgs = 0.95
+ wkt1 = -2.0389865e-9
+ wkt2 = 1.7872759e-9
+ lvoff = -9.7335308e-9
+ wmax = 5.374e-7
+ aigc = 0.0068257672
+ wmin = 2.674e-7
+ tcjswg = 0.00128
+ lvsat = -0.00028
+ lvth0 = -1.2456137e-8
+ delta = 0.018814
+ laigc = -3.7754415e-11
+ wua1 = 1.7501635e-16
+ wub1 = -7.9730823e-26
+ wuc1 = 2.9760508e-17
+ fnoimod = 1
+ rnoia = 0
+ rnoib = 0
+ bigc = 0.0012521
+ eigbinv = 1.1
+ wute = 3.4211506e-8
+ wwlc = 0
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ pketa = -2.4999571e-14
+ ngate = 1.7e+20
+ cdsc = 0
+ ngcon = 1
+ cgbo = 0
+ wpclm = -1.1447315e-8
+ cgdl = 3.2212350000000004e-11
+ cgdo = 2.8335740000000002e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.2212350000000004e-11
+ cgso = 2.8335740000000002e-11
+ fprout = 200
+ cigc = 0.15259
+ gbmin = 1e-12
+ xrcrg1 = 12
+ xrcrg2 = 1
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ cigbacc = 0.245
+ wtvoff = -1.02826e-10
+ tnoimod = 0
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ capmod = 2
+ cigbinv = 0.006
+ wku0we = 1.5e-11
+ k2we = 5e-5
+ mobmod = 0
+ ijthsfwd = 0.01
+ dsub = 0.5
+ dtox = 3.91e-10
+ tvoff = 0.0027071394
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ xjbvd = 1
+ xjbvs = 1
+ version = 4.5
+ lk2we = 0.0
+ tempmod = 0
+ eta0 = 0.17962267
+ etab = -0.19577778
+ ijthsrev = 0.01
+ ku0we = -0.0007
+ aigbacc = 0.012071
+ beta0 = 13.32
+ leta0 = 6e-10
+ laigsd = 1.0132005e-13
+ ppclm = 0
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ aigbinv = 0.009974
+ ppdiblc2 = -7.3176658e-16
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ )

.model pch_ff_27 pmos (
+ level = 54
+ tvfbsdoff = 0.1
+ fnoimod = 1
+ scref = 1e-6
+ eigbinv = 1.1
+ rshg = 14.1
+ ltvoff = -3.7535707e-10
+ pigcd = 2.572
+ aigsd = 0.0063633912
+ lvoff = -1.1639377e-8
+ lvsat = -0.00028
+ lvth0 = 1.3506701e-9
+ ijthsfwd = 0.01
+ lku0we = 1.8e-11
+ delta = 0.018814
+ laigc = -5.5983746e-11
+ epsrox = 3.9
+ tnom = 25
+ rnoia = 0
+ rnoib = 0
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ cigbacc = 0.245
+ toxe = 2.6300000000000002e-9
+ toxm = 2.67e-9
+ rdsmod = 0
+ igbmod = 1
+ pketa = 5.6398736e-15
+ ngate = 1.7e+20
+ wtvfbsdoff = 0
+ ijthsrev = 0.01
+ ngcon = 1
+ tnoimod = 0
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ wpclm = -1.1447315e-8
+ pbswgd = 0.8
+ pbswgs = 0.8
+ gbmin = 1e-12
+ cigbinv = 0.006
+ jswgd = 3.69e-13
+ ltvfbsdoff = 0
+ jswgs = 3.69e-13
+ igcmod = 1
+ wags = 3.4820603e-7
+ voff = -0.10461895
+ acde = 0.5
+ version = 4.5
+ ppdiblc2 = 9.4893758e-16
+ vsat = 91103.982
+ tempmod = 0
+ wint = 0
+ vth0 = -0.36207681999999997
+ wkt1 = 1.4552168e-8
+ wkt2 = 6.9668931e-9
+ wmax = 5.374e-7
+ aigc = 0.0068462496
+ wmin = 2.674e-7
+ aigbacc = 0.012071
+ ptvfbsdoff = 0
+ tvoff = 0.0026312893
+ wua1 = 1.777316e-16
+ wub1 = 1.5048515e-26
+ wuc1 = -3.1929257e-17
+ permod = 1
+ xjbvd = 1
+ xjbvs = 1
+ bigc = 0.0012521
+ wute = 6.965504e-8
+ lk2we = 0.0
+ wwlc = 0
+ pkvth0we = 0.0
+ aigbinv = 0.009974
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.2212350000000004e-11
+ cgdo = 2.8335740000000002e-11
+ xtid = 3
+ xtis = 3
+ ku0we = -0.0007
+ beta0 = 13.32
+ cgsl = 3.2212350000000004e-11
+ cgso = 2.8335740000000002e-11
+ voffcv = -0.125
+ wpemod = 1
+ cigc = 0.15259
+ vfbsdoff = 0.01
+ leta0 = 6e-10
+ ppclm = 0
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ paramchk = 1
+ poxedge = 1
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ binunit = 2
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ tpbswg = 0.001
+ k2we = 5e-5
+ ijthdfwd = 0.01
+ dsub = 0.5
+ dtox = 3.91e-10
+ a0 = 2.4559917
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 72000
+ cf = 8.741900000000001e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.0065510297
+ k3 = -2.5823
+ em = 20000000.0
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ ll = 0
+ lw = 0
+ u0 = 0.010769968
+ w0 = 0
+ ua = 2.2475737e-10
+ ub = 1.3971204e-18
+ uc = 8.9671176e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 2.33e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ bigsd = 0.0003327
+ ptvoff = 6.0034078e-17
+ eta0 = 0.17962267
+ etab = -0.19577778
+ waigsd = 1.9297907e-12
+ wvoff = -2.3606869e-9
+ ijthdrev = 0.01
+ wvsat = 0.0034765009
+ diomod = 1
+ wvth0 = 1.5832152000000002e-9
+ lpdiblc2 = -1.0873556e-9
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ waigc = -6.0221967e-12
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.6832999999999998e-10
+ pku0we = 0.0
+ cjswgs = 1.6832999999999998e-10
+ lketa = -2.7133526e-8
+ xpart = 1
+ mjswgd = 0.95
+ mjswgs = 0.95
+ egidl = 0.001
+ tcjswg = 0.00128
+ pvfbsdoff = 0
+ lkvth0we = 3e-12
+ njtsswg = 6.489
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ acnqsmod = 0
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.012575691
+ pdiblcb = 0
+ rbodymod = 0
+ fprout = 200
+ xrcrg1 = 12
+ xrcrg2 = 1
+ pvoff = 1.5239261e-15
+ keta = 0.0057304489
+ cdscb = 0
+ cdscd = 0
+ pvsat = 0
+ bigbacc = 0.0054401
+ lags = 9.833094e-7
+ wk2we = 0.0
+ pvth0 = 2.7595820000000008e-17
+ wtvoff = -1.9743529e-10
+ drout = 0.56
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 6.2671111e-11
+ paigc = 6.5097646e-18
+ kt1l = 0
+ kvth0we = -0.00022
+ voffl = 0
+ wpdiblc2 = -1.8846129e-9
+ lintnoi = -5e-9
+ capmod = 2
+ lint = 6.5375218e-9
+ bigbinv = 0.00149
+ weta0 = -1.7368176e-8
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ wetab = 1.9534667e-8
+ wku0we = 1.5e-11
+ lkt1 = -3.7329349e-9
+ lkt2 = -2.567581e-9
+ lpclm = 0
+ lmax = 9.0075e-7
+ lmin = 4.5075e-7
+ mobmod = 0
+ lpe0 = 6.44e-8
+ lpeb = 0
+ cgidl = 1
+ minv = -0.33
+ lua1 = 1.3348283e-16
+ lub1 = 2.1611253e-25
+ luc1 = 5.928335e-17
+ ndep = 1e+18
+ lute = 1.2896693e-7
+ wkvth0we = 0.0
+ lwlc = 0
+ moin = 5.5538
+ pbswd = 0.9
+ pbsws = 0.9
+ ags = -0.056621626
+ nigc = 2.291
+ trnqsmod = 0
+ cjd = 0.0012517799999999999
+ cit = -8.7888889e-5
+ cjs = 0.0012517799999999999
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 1.0572421799999999e-8
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ pdits = 0
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ cigsd = 0.013281
+ nfactor = 1
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ la0 = -1.8333262e-7
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = -0.0008
+ pags = -2.41252e-13
+ kt1 = -0.20789546
+ kt2 = -0.0733757
+ lk2 = -1.6954158000000002e-10
+ llc = 0
+ lln = 1
+ lu0 = -3.3434965000000003e-10
+ mjd = 0.335
+ mjs = 0.335
+ lua = -5.402342e-17
+ lub = -8.029291e-26
+ luc = -6.9221885e-17
+ lud = 0
+ ntox = 2.958
+ lwc = 0
+ lwl = 0
+ pcit = 1e-18
+ lwn = 1
+ pclm = 1.1689658
+ njd = 1.02
+ njs = 1.02
+ pa0 = -1.295362e-13
+ rgatemod = 0
+ nsd = 1e+20
+ pbd = 0.75
+ pk2we = 0.0
+ pat = 0
+ pbs = 0.75
+ pk2 = 6.34174e-16
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ tnjtsswg = 1
+ pu0 = -2.5304972e-16
+ prt = 0
+ pua = -1.1377853e-22
+ pub = 1.1787175e-31
+ puc = 2.8393052e-23
+ pud = 0
+ phin = 0.15
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 1.5353037e-9
+ ub1 = -2.5129786e-18
+ uc1 = 1.2019494e-10
+ tpb = 0.0016
+ tnoia = 0
+ wa0 = 1.4554629e-7
+ pkt1 = -1.0156873999999999e-14
+ pkt2 = -7.3243565e-16
+ ute = -1.2205289
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 2.3228278e-9
+ nigbacc = 10
+ wlc = 0
+ wln = 1
+ wu0 = 3.4013886e-10
+ xgl = -8.2e-9
+ xgw = 0
+ peta0 = 2e-17
+ wua = -1.1141771e-17
+ wub = -5.4878553e-26
+ wuc = -2.8229789e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ wketa = -8.9579586e-9
+ tpbsw = 0.0025
+ cjswd = 4.743e-11
+ cjsws = 4.743e-11
+ rbdb = 50
+ pua1 = -9.6760461e-23
+ prwb = 0
+ pub1 = 5.7312604e-33
+ prwg = 0
+ puc1 = -1.747778e-23
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ nigbinv = 2.171
+ pute = -4.8084303e-14
+ rdsw = 200
+ toxref = 3e-9
+ )

.model pch_ff_28 pmos (
+ level = 54
+ wtvfbsdoff = 0
+ lku0we = 1.8e-11
+ k2we = 5e-5
+ epsrox = 3.9
+ dsub = 0.5
+ dtox = 3.91e-10
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ ltvfbsdoff = 0
+ bigbacc = 0.0054401
+ rdsmod = 0
+ igbmod = 1
+ wkvth0we = 0.0
+ eta0 = 0.17962267
+ etab = -0.19577778
+ kvth0we = -0.00022
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ trnqsmod = 0
+ pbswgd = 0.8
+ lintnoi = -5e-9
+ pbswgs = 0.8
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ pvoff = -2.5154209e-16
+ igcmod = 1
+ cdscb = 0
+ cdscd = 0
+ pvsat = 0
+ wk2we = 0.0
+ pvth0 = -5.467691400000001e-16
+ ptvfbsdoff = 0
+ drout = 0.56
+ paigc = -3.9499473e-18
+ voffl = 0
+ rgatemod = 0
+ tnjtsswg = 1
+ weta0 = -1.7368176e-8
+ wetab = 1.9534667e-8
+ lpclm = 0
+ cgidl = 1
+ permod = 1
+ ags = -1.2539967
+ nfactor = 1
+ cjd = 0.0012517799999999999
+ cit = -0.00036538451
+ cjs = 0.0012517799999999999
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 1.38228675e-8
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ pbswd = 0.9
+ pbsws = 0.9
+ voffcv = -0.125
+ wpemod = 1
+ la0 = -4.7253353e-7
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = -0.0008
+ kt1 = -0.16257215
+ kt2 = -0.066291072
+ lk2 = 5.244707700000001e-10
+ llc = -1.18e-13
+ lln = 0.7
+ lu0 = -5.5490454e-10
+ keta = -0.0061234738
+ mjd = 0.335
+ mjs = 0.335
+ lua = -1.0290148e-16
+ lub = -5.3060964e-27
+ luc = -4.0794824e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pdits = 0
+ pa0 = 9.7298482e-15
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ cigsd = 0.013281
+ pk2 = -2.0891363e-16
+ nigbacc = 10
+ lags = 1.5101544e-6
+ pu0 = 1.1540053e-17
+ dvt0w = 0
+ dvt1w = 0
+ prt = 0
+ dvt2w = 0
+ pua = -1.3867635e-23
+ pub = 2.1855871e-32
+ puc = -2.7646346e-24
+ pud = 0
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 1.8476918e-10
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 1.7313241e-9
+ ub1 = -1.3316629e-18
+ uc1 = 2.2670111e-10
+ kt1l = 0
+ tpb = 0.0016
+ wa0 = -1.7096745e-7
+ ute = -0.86054925
+ web = 6628.3
+ wec = -16935.0
+ pk2we = 0.0
+ wk2 = 4.238936e-9
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ wlc = 0
+ wln = 1
+ wu0 = -2.6120153e-10
+ xgl = -8.2e-9
+ xgw = 0
+ wua = -2.3821198e-16
+ wub = 1.6333936e-25
+ wuc = 4.2583136e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ nigbinv = 2.171
+ lint = 9.7879675e-9
+ tpbswg = 0.001
+ lkt1 = -2.3675192e-8
+ lkt2 = -5.6848171e-9
+ lmax = 4.5075e-7
+ tnoia = 0
+ lmin = 2.1744e-7
+ lpe0 = 6.44e-8
+ ijthsfwd = 0.01
+ lpeb = 0
+ peta0 = 2e-17
+ wketa = -7.8373297e-10
+ minv = -0.33
+ tpbsw = 0.0025
+ lua1 = 4.723388e-17
+ lub1 = -3.0366637e-25
+ luc1 = 1.2420632e-17
+ ptvoff = 5.0195791e-17
+ cjswd = 4.743e-11
+ cjsws = 4.743e-11
+ ndep = 1e+18
+ fnoimod = 1
+ mjswd = 0.01
+ lute = -2.9424109e-8
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ waigsd = 1.9297907e-12
+ lwlc = 0
+ eigbinv = 1.1
+ moin = 5.5538
+ ijthsrev = 0.01
+ nigc = 2.291
+ diomod = 1
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.6832999999999998e-10
+ pku0we = 0.0
+ cjswgs = 1.6832999999999998e-10
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ tvfbsdoff = 0.1
+ pags = -3.3771496e-13
+ scref = 1e-6
+ a0 = 3.1132665
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 72000
+ cf = 8.741900000000001e-11
+ ntox = 2.958
+ mjswgd = 0.95
+ ef = 1.15
+ mjswgs = 0.95
+ k1 = 0.30425
+ k2 = -0.0081283305
+ k3 = -2.5823
+ pcit = -8.2716403e-18
+ em = 20000000.0
+ ppdiblc2 = -3.8737293e-16
+ pclm = 1.1689658
+ pigcd = 2.572
+ cigbacc = 0.245
+ ll = -1.18e-13
+ aigsd = 0.0063633912
+ lw = 0
+ u0 = 0.01127123
+ w0 = 0
+ ua = 3.3584387e-10
+ ub = 1.2266958e-18
+ uc = -5.8379738e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 2.33e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ tcjswg = 0.00128
+ lvoff = -4.2658924e-9
+ phin = 0.15
+ tnoimod = 0
+ lvsat = -0.00028
+ pkt1 = 6.8855166e-15
+ pkt2 = 2.2627554e-16
+ lvth0 = 4.8653579e-9
+ cigbinv = 0.006
+ delta = 0.018814
+ laigc = -1.8017042e-11
+ wvfbsdoff = 0
+ rnoia = 0
+ rnoib = 0
+ lvfbsdoff = 0
+ rbdb = 50
+ pua1 = -2.7108228e-23
+ pkvth0we = 0.0
+ prwb = 0
+ pub1 = 7.1177686e-32
+ prwg = 0
+ puc1 = 8.7727027e-25
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ pketa = 2.0432143e-15
+ version = 4.5
+ ngate = 1.7e+20
+ pute = 1.6065563e-14
+ fprout = 200
+ rdsw = 200
+ ngcon = 1
+ tempmod = 0
+ wpclm = -1.1447315e-8
+ xrcrg1 = 12
+ xrcrg2 = 1
+ vfbsdoff = 0.01
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ aigbacc = 0.012071
+ wtvoff = -1.7507555e-10
+ paramchk = 1
+ rshg = 14.1
+ capmod = 2
+ aigbinv = 0.009974
+ wku0we = 1.5e-11
+ mobmod = 0
+ ijthdfwd = 0.01
+ tvoff = 0.002323434
+ tnom = 25
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ toxe = 2.6300000000000002e-9
+ toxm = 2.67e-9
+ poxedge = 1
+ ijthdrev = 0.01
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = 6e-10
+ lpdiblc2 = 4.7505822e-10
+ binunit = 2
+ ppclm = 0
+ wags = 5.6744004e-7
+ wcit = 2.107191e-11
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ voff = -0.12137687
+ acde = 0.5
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ vsat = 91103.982
+ wint = 0
+ vth0 = -0.37006475000000005
+ wkt1 = -2.4180539e-8
+ wkt2 = 4.7880041e-9
+ wmax = 5.374e-7
+ dmcgt = 0
+ aigc = 0.0067599617
+ wmin = 2.674e-7
+ tcjsw = 9.34e-5
+ lkvth0we = 3e-12
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ wua1 = 1.9431072e-17
+ wub1 = -1.3369336e-25
+ wuc1 = -7.3645279e-17
+ acnqsmod = 0
+ bigc = 0.0012521
+ bigsd = 0.0003327
+ wute = -7.6140111e-8
+ wwlc = 0
+ wvoff = 1.674468e-9
+ toxref = 3e-9
+ rbodymod = 0
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.2212350000000004e-11
+ cgdo = 2.8335740000000002e-11
+ xtid = 3
+ xtis = 3
+ wvsat = 0.0034765009
+ cgsl = 3.2212350000000004e-11
+ cgso = 2.8335740000000002e-11
+ wvth0 = 2.8885901000000003e-9
+ cigc = 0.15259
+ waigc = 1.7749876e-11
+ njtsswg = 6.489
+ lketa = -2.19178e-8
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ ltvoff = -2.3990075e-10
+ xpart = 1
+ ckappad = 0.6
+ wpdiblc2 = 1.1524564e-9
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.0090247504
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ pdiblcb = 0
+ egidl = 0.001
+ pvfbsdoff = 0
+ )

.model pch_ff_29 pmos (
+ level = 54
+ ijthdrev = 0.01
+ ngcon = 1
+ pbswgd = 0.8
+ pbswgs = 0.8
+ wpclm = -1.2079184e-7
+ aigbinv = 0.009974
+ nigc = 2.291
+ igcmod = 1
+ lpdiblc2 = -1.1954251e-9
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ ntox = 2.958
+ pcit = -7.1298391e-18
+ pclm = 1.5407845
+ poxedge = 1
+ phin = 0.15
+ lkvth0we = 3e-12
+ pkt1 = -1.16482e-15
+ pkt2 = -1.4992738e-15
+ binunit = 2
+ permod = 1
+ tvoff = 0.00085372815
+ acnqsmod = 0
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ rbdb = 50
+ pua1 = 1.9617826e-23
+ prwb = 0
+ pub1 = -3.1346313e-32
+ prwg = 0
+ puc1 = 1.1713402e-23
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ rbodymod = 0
+ voffcv = -0.125
+ wpemod = 1
+ rdsw = 200
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = 6e-10
+ ppclm = 2.3071337e-14
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ rshg = 14.1
+ wpdiblc2 = -7.3926191e-10
+ tpbswg = 0.001
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ njtsswg = 6.489
+ ptvoff = -3.132788e-17
+ tnom = 25
+ bigsd = 0.0003327
+ waigsd = 1.9297907e-12
+ toxe = 2.6300000000000002e-9
+ toxm = 2.67e-9
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ wkvth0we = 0.0
+ wvoff = 3.1859801e-10
+ diomod = 1
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.016941733
+ trnqsmod = 0
+ pdiblcb = 0
+ wvsat = 0.0032472346
+ pditsd = 0
+ wvth0 = -2.2669424999999996e-9
+ pditsl = 0
+ cjswgd = 1.6832999999999998e-10
+ pku0we = 0.0
+ cjswgs = 1.6832999999999998e-10
+ waigc = -1.7260908e-11
+ wags = -1.0331048e-6
+ wcit = 1.566053e-11
+ lketa = 7.1935383e-9
+ voff = -0.13201276
+ mjswgd = 0.95
+ mjswgs = 0.95
+ bigbacc = 0.0054401
+ acde = 0.5
+ xpart = 1
+ rgatemod = 0
+ tcjswg = 0.00128
+ vsat = 91523.884
+ wint = 0
+ tnjtsswg = 1
+ vth0 = -0.36762236000000004
+ pvfbsdoff = 0
+ kvth0we = -0.00022
+ egidl = 0.001
+ wkt1 = 1.3972715e-8
+ wkt2 = 1.2965963e-8
+ wmax = 5.374e-7
+ aigc = 0.0067957378
+ wmin = 2.674e-7
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ wua1 = -2.0201942e-16
+ wub1 = 3.5220237e-25
+ wuc1 = -1.2500135e-16
+ bigc = 0.0012521
+ wwlc = 0
+ fprout = 200
+ cdsc = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ a0 = 1.1444157
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ cgbo = 0
+ cgdl = 3.2212350000000004e-11
+ cgdo = 2.8335740000000002e-11
+ at = 108550.2
+ xtid = 3
+ cf = 8.741900000000001e-11
+ xtis = 3
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.025395241
+ k3 = -2.5823
+ em = 20000000.0
+ ll = -1.18e-13
+ lw = 0
+ u0 = 0.0096317592
+ cgsl = 3.2212350000000004e-11
+ cgso = 2.8335740000000002e-11
+ w0 = 0
+ ua = -3.1599722e-11
+ ub = 1.4008434e-18
+ uc = -1.6299488e-10
+ ud = 0
+ cigc = 0.15259
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 2.33e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ pvoff = 3.4546471000000004e-17
+ wtvoff = 2.1129256e-10
+ cdscb = 0
+ cdscd = 0
+ pvsat = 4.83709e-11
+ wk2we = 0.0
+ pvth0 = 5.4104824e-16
+ drout = 0.56
+ paigc = 3.4373281e-18
+ nfactor = 1
+ capmod = 2
+ voffl = 0
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ wku0we = 1.5e-11
+ dmdg = 0
+ weta0 = -1.7368176e-8
+ wetab = 1.9534667e-8
+ mobmod = 0
+ ags = 5.9031333
+ lpclm = -7.8453093e-8
+ cjd = 0.0012517799999999999
+ cit = 0.00015305446
+ cjs = 0.0012517799999999999
+ clc = 1e-7
+ cle = 0.6
+ k2we = 5e-5
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 1.38228675e-8
+ ijthsfwd = 0.01
+ k3b = 2.1176
+ dsub = 0.5
+ cgidl = 1
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ dtox = 3.91e-10
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ nigbacc = 10
+ la0 = -5.7105222e-8
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = -0.0085120921
+ kt1 = -0.27233533
+ kt2 = -0.10755274
+ lk2 = 4.167788899999999e-9
+ eta0 = 0.17962267
+ llc = -1.18e-13
+ lln = 0.7
+ lu0 = -2.0897630000000002e-10
+ etab = -0.19577778
+ mjd = 0.335
+ mjs = 0.335
+ lua = -2.5370884e-17
+ lub = -4.2051244e-26
+ luc = 1.7994313e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ pbswd = 0.9
+ pbsws = 0.9
+ njd = 1.02
+ njs = 1.02
+ pa0 = -3.159814e-15
+ ijthsrev = 0.01
+ nsd = 1e+20
+ pbd = 0.75
+ pat = -4.5415452e-10
+ pbs = 0.75
+ pk2 = -2.0710507e-16
+ pu0 = 4.0684676e-18
+ prt = 0
+ pua = 6.5898257e-24
+ pub = -4.9701536e-33
+ puc = -7.066739e-24
+ pud = 0
+ nigbinv = 2.171
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 2.8369875e-9
+ ub1 = -4.0389099e-18
+ uc1 = 4.2708978e-10
+ tpb = 0.0016
+ wa0 = -1.0988104e-7
+ pdits = 0
+ ute = -1
+ wat = 0.0021523911
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 4.2303646e-9
+ cigsd = 0.013281
+ wlc = 0
+ wln = 1
+ wu0 = -2.2579117e-10
+ xgl = -8.2e-9
+ xgw = 0
+ wua = -3.3516677e-16
+ dvt0w = 0
+ wub = 2.9047692e-25
+ wuc = 6.2972257e-17
+ wud = 0
+ dvt1w = 0
+ dvt2w = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ ppdiblc2 = 1.1779633e-17
+ pk2we = 0.0
+ fnoimod = 1
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ eigbinv = 1.1
+ tnoia = 0
+ peta0 = 2e-17
+ wketa = 1.4826965e-8
+ tpbsw = 0.0025
+ cjswd = 4.743e-11
+ cjsws = 4.743e-11
+ pkvth0we = 0.0
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ toxref = 3e-9
+ cigbacc = 0.245
+ vfbsdoff = 0.01
+ tnoimod = 0
+ keta = -0.1440919
+ tvfbsdoff = 0.1
+ wtvfbsdoff = 0
+ cigbinv = 0.006
+ ltvoff = 7.0207177e-11
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 7.537856e-11
+ paramchk = 1
+ scref = 1e-6
+ kt1l = 0
+ pigcd = 2.572
+ aigsd = 0.0063633912
+ ltvfbsdoff = 0
+ version = 4.5
+ lvoff = -2.0217201e-9
+ lint = 9.7879675e-9
+ tempmod = 0
+ lkt1 = -5.151622e-10
+ lkt2 = 3.021395e-9
+ lku0we = 1.8e-11
+ lmax = 2.1744e-7
+ lvsat = -0.00036859139999999996
+ lmin = 9.167e-8
+ epsrox = 3.9
+ lvth0 = 4.3500147e-9
+ lpe0 = 6.44e-8
+ ijthdfwd = 0.01
+ lpeb = 0
+ delta = 0.018814
+ laigc = -2.5565813e-11
+ aigbacc = 0.012071
+ wvfbsdoff = 0
+ rdsmod = 0
+ lvfbsdoff = 0
+ minv = -0.33
+ rnoia = 0
+ rnoib = 0
+ lua1 = -1.8606111e-16
+ lub1 = 2.6756274e-25
+ luc1 = -2.9861377e-17
+ igbmod = 1
+ ndep = 1e+18
+ ptvfbsdoff = 0
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ lwlc = 0
+ pketa = -1.250643e-15
+ ngate = 1.7e+20
+ moin = 5.5538
+ )

.model pch_ff_30 pmos (
+ level = 54
+ ijthdrev = 0.01
+ ngcon = 1
+ pbswgd = 0.8
+ pbswgs = 0.8
+ wpclm = 4.9341412e-7
+ aigbinv = 0.009974
+ nigc = 2.291
+ igcmod = 1
+ lpdiblc2 = 0
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ ntox = 2.958
+ pcit = 6.654835000000001e-18
+ pclm = 0.08631615
+ paigsd = 8.4526218e-25
+ poxedge = 1
+ phin = 0.15
+ lkvth0we = 3e-12
+ pkt1 = -1.6624191e-15
+ pkt2 = 2.1480498e-17
+ binunit = 2
+ permod = 1
+ tvoff = 0.0012365685
+ acnqsmod = 0
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ rbdb = 50
+ pua1 = 4.1792962e-25
+ prwb = 0
+ pub1 = 6.1746384e-33
+ prwg = 0
+ puc1 = 2.9246063e-24
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ rbodymod = 0
+ voffcv = -0.125
+ wpemod = 1
+ rdsw = 200
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = -7.965883199999999e-9
+ letab = 1.7579973e-8
+ ppclm = -3.4664022e-14
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ rshg = 14.1
+ wpdiblc2 = -6.1394667e-10
+ tpbswg = 0.001
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ njtsswg = 6.489
+ ptvoff = 2.0376593e-17
+ tnom = 25
+ bigsd = 0.0003327
+ waigsd = 1.9297817e-12
+ toxe = 2.6300000000000002e-9
+ toxm = 2.67e-9
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ wkvth0we = 0.0
+ wvoff = -2.8254962e-9
+ diomod = 1
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.0042244444
+ trnqsmod = 0
+ pdiblcb = 0
+ wvsat = 0.017016245
+ pditsd = 0
+ wvth0 = -2.9016160999999997e-9
+ pditsl = 0
+ cjswgd = 1.6832999999999998e-10
+ pku0we = 0.0
+ cjswgs = 1.6832999999999998e-10
+ waigc = 7.1461687e-12
+ wags = -1.0331048e-6
+ wcit = -1.3098452e-10
+ lketa = -1.1878561e-8
+ voff = -0.12098873
+ mjswgd = 0.95
+ mjswgs = 0.95
+ bigbacc = 0.0054401
+ acde = 0.5
+ xpart = 1
+ rgatemod = 0
+ tcjswg = 0.00128
+ vsat = 62231.739
+ wint = 0
+ tnjtsswg = 1
+ vth0 = -0.30655978
+ pvfbsdoff = 0
+ kvth0we = -0.00022
+ egidl = 0.001
+ wkt1 = 1.9266322e-8
+ wkt2 = -3.2122744e-9
+ wmax = 5.374e-7
+ aigc = 0.0067006504
+ wmin = 2.674e-7
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ wua1 = 2.2347963e-18
+ wub1 = -4.6956688e-26
+ wuc1 = -3.1503526e-17
+ bigc = 0.0012521
+ wwlc = 0
+ fprout = 200
+ cdsc = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ a0 = 3.9744452
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ cgbo = 0
+ cgdl = 3.2212350000000004e-11
+ cgdo = 2.8335740000000002e-11
+ at = 69068.642
+ xtid = 3
+ cf = 8.741900000000001e-11
+ xtis = 3
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.022825095
+ k3 = -2.5823
+ em = 20000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.0037956963000000004
+ cgsl = 3.2212350000000004e-11
+ cgso = 2.8335740000000002e-11
+ w0 = 0
+ ua = -9.2439852e-11
+ ub = -1.8842125e-18
+ uc = 5.3507127e-11
+ ud = 0
+ cigc = 0.15259
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 2.33e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ pvoff = 3.3009131999999996e-16
+ wtvoff = -3.3875503e-10
+ cdscb = 0
+ cdscd = 0
+ pvsat = -1.2459161e-9
+ wk2we = 0.0
+ pvth0 = 6.0070714e-16
+ drout = 0.56
+ paigc = 1.1430629e-18
+ nfactor = 1
+ capmod = 2
+ voffl = 0
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ wku0we = 1.5e-11
+ dmdg = 0
+ weta0 = -5.4735839e-8
+ wetab = 4.6876459e-8
+ mobmod = 0
+ ags = 5.9031333
+ lpclm = 5.8266931e-8
+ cjd = 0.0012517799999999999
+ cit = 0.00059801095
+ cjs = 0.0012517799999999999
+ clc = 1e-7
+ cle = 0.6
+ k2we = 5e-5
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 4.0349e-9
+ ijthsfwd = 0.01
+ k3b = 2.1176
+ dsub = 0.5
+ cgidl = 1
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ dtox = 3.91e-10
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ nigbacc = 10
+ la0 = -3.23128e-7
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = -0.0048008257000000006
+ kt1 = -0.32608492
+ kt2 = -0.08284588
+ lk2 = 3.9261952e-9
+ eta0 = 0.27074908
+ llc = 0
+ lln = 1
+ lu0 = 3.3961361999999997e-10
+ etab = -0.38279877
+ mjd = 0.335
+ mjs = 0.335
+ lua = -1.9651912e-17
+ lub = 2.6674400999999997e-25
+ luc = -2.356876e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ pbswd = 0.9
+ pbsws = 0.9
+ njd = 1.02
+ njs = 1.02
+ pa0 = 9.1746422e-14
+ laigsd = -3.0625433e-18
+ ijthsrev = 0.01
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 6.7620954e-11
+ pbs = 0.75
+ pk2 = 2.5170462e-16
+ pu0 = -8.2666616e-17
+ prt = 0
+ pua = 3.032424e-23
+ pub = -1.03773645e-31
+ puc = -2.0363205e-24
+ pud = 0
+ nigbinv = 2.171
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = -2.7998083e-10
+ ub1 = 8.7083504e-19
+ uc1 = 1.8820988e-11
+ tpb = 0.0016
+ wa0 = -1.1195219e-6
+ pdits = 0
+ ute = -1
+ wat = -0.0033984119
+ web = 6628.3
+ wec = -16935.0
+ wk2 = -6.5058945e-10
+ cigsd = 0.013281
+ wlc = 0
+ wln = 1
+ wu0 = 6.9692249e-10
+ xgl = -8.2e-9
+ xgw = 0
+ wua = -5.8766054e-16
+ dvt0w = 0
+ wub = 1.3415779e-24
+ wuc = 9.4571662e-18
+ wud = 0
+ dvt1w = 0
+ dvt2w = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ ppdiblc2 = 0
+ pk2we = 0.0
+ fnoimod = 1
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ eigbinv = 1.1
+ tnoia = 0
+ peta0 = 3.5325603e-15
+ petab = -2.5701285e-15
+ wketa = -3.6489897e-8
+ tpbsw = 0.0025
+ cjswd = 4.743e-11
+ cjsws = 4.743e-11
+ pkvth0we = 0.0
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ toxref = 3e-9
+ cigbacc = 0.245
+ vfbsdoff = 0.01
+ tnoimod = 0
+ keta = 0.058802768
+ tvfbsdoff = 0.1
+ wtvfbsdoff = 0
+ cigbinv = 0.006
+ ltvoff = 3.4220189e-11
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 3.355326999999999e-11
+ paramchk = 1
+ scref = 1e-6
+ kt1l = 0
+ pigcd = 2.572
+ aigsd = 0.0063633912
+ ltvfbsdoff = 0
+ version = 4.5
+ lvoff = -3.0579783e-9
+ lint = 0
+ tempmod = 0
+ lkt1 = 4.537299899999999e-9
+ lkt2 = 6.989501e-10
+ lku0we = 1.8e-11
+ lmax = 9.167e-8
+ lvsat = 0.0023848703
+ lmin = 5.567e-8
+ epsrox = 3.9
+ lvth0 = -1.3898688e-9
+ lpe0 = 6.44e-8
+ ijthdfwd = 0.01
+ lpeb = 0
+ delta = 0.018814
+ laigc = -1.6627591e-11
+ aigbacc = 0.012071
+ wvfbsdoff = 0
+ rdsmod = 0
+ lvfbsdoff = 0
+ minv = -0.33
+ rnoia = 0
+ rnoib = 0
+ lua1 = 1.0693391e-16
+ lub1 = -1.9395329e-25
+ luc1 = 8.5158894e-18
+ igbmod = 1
+ ndep = 1e+18
+ ptvfbsdoff = 0
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ lwlc = 0
+ pketa = 3.573142e-15
+ ngate = 1.7e+20
+ moin = 5.5538
+ )

.model pch_ff_31 pmos (
+ level = 54
+ paigc = -3.8652128e-18
+ voff = -0.11425646
+ nigbacc = 10
+ ags = 5.9031333
+ acde = 0.5
+ ppdiblc2 = 0
+ voffl = 0
+ cjd = 0.0012517799999999999
+ cit = 0.0026900602000000003
+ cjs = 0.0012517799999999999
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ vsat = 249488.49
+ dlc = 4.0349e-9
+ wint = 0
+ k3b = 2.1176
+ vth0 = -0.31696792000000007
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ weta0 = 4.5849198e-8
+ wkt1 = -9.053012e-8
+ wkt2 = -4.5663135e-8
+ wetab = 2.1214781e-8
+ wmax = 5.374e-7
+ aigc = 0.0065523001
+ wmin = 2.674e-7
+ lpclm = -1.6067206e-7
+ permod = 1
+ nigbinv = 2.171
+ la0 = 2.2449695e-9
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = -0.00174527867
+ kt1 = -0.078489325
+ kt2 = 0.051187672
+ lk2 = 5.0231101e-9
+ llc = 0
+ lln = 1
+ cgidl = 1
+ lu0 = -6.534920299999999e-10
+ mjd = 0.335
+ mjs = 0.335
+ lua = -5.2618623e-17
+ lub = -3.591586e-25
+ luc = -2.0280652e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ wua1 = 2.8402308e-15
+ njs = 1.02
+ wub1 = -3.9062366e-24
+ wuc1 = 2.0276364e-16
+ pa0 = -4.432942e-14
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 1.8264736e-9
+ pbs = 0.75
+ pk2 = -1.1995676e-16
+ pu0 = 2.2577126e-16
+ bigc = 0.0012521
+ prt = 0
+ pua = 1.5923531e-23
+ pub = 1.06100166e-31
+ puc = 3.3504384e-24
+ pud = 0
+ wwlc = 0
+ pkvth0we = 0.0
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = -3.345352e-9
+ ub1 = 3.9080279e-18
+ uc1 = 1.4308247e-10
+ tpb = 0.0016
+ voffcv = -0.125
+ wpemod = 1
+ pbswd = 0.9
+ pbsws = 0.9
+ wa0 = 1.2266134e-6
+ cdsc = 0
+ ute = -1
+ wat = -0.033723458
+ web = 6628.3
+ wec = -16935.0
+ fnoimod = 1
+ wk2 = 5.7573654e-9
+ wlc = 0
+ cgbo = 0
+ wln = 1
+ cgdl = 3.2212350000000004e-11
+ cgdo = 2.8335740000000002e-11
+ wu0 = -4.6209719e-9
+ xtid = 3
+ xgl = -8.2e-9
+ xtis = 3
+ xgw = 0
+ wua = -3.3937245e-16
+ wub = -2.2769359e-24
+ wuc = -8.3417988e-17
+ wud = 0
+ eigbinv = 1.1
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ cgsl = 3.2212350000000004e-11
+ cgso = 2.8335740000000002e-11
+ vfbsdoff = 0.01
+ cigc = 0.15259
+ pdits = 0
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ paramchk = 1
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ tpbswg = 0.001
+ cigbacc = 0.245
+ tnoia = 0
+ k2we = 5e-5
+ tnoimod = 0
+ ijthdfwd = 0.01
+ peta0 = -2.3013718000000002e-15
+ dsub = 0.5
+ petab = -1.0817512e-15
+ dtox = 3.91e-10
+ wketa = 7.0696889e-8
+ ptvoff = -1.3332507e-17
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ tpbsw = 0.0025
+ waigsd = 1.9297962e-12
+ cigbinv = 0.006
+ cjswd = 4.743e-11
+ cjsws = 4.743e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ eta0 = 0.012687945
+ etab = -0.23454709
+ diomod = 1
+ ijthdrev = 0.01
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.6832999999999998e-10
+ pku0we = 0.0
+ version = 4.5
+ cjswgs = 1.6832999999999998e-10
+ lpdiblc2 = 0
+ tempmod = 0
+ tvfbsdoff = 0.1
+ aigbacc = 0.012071
+ mjswgd = 0.95
+ mjswgs = 0.95
+ scref = 1e-6
+ tcjswg = 0.00128
+ pigcd = 2.572
+ aigsd = 0.0063633912
+ lvoff = -3.4484499e-9
+ lkvth0we = 3e-12
+ aigbinv = 0.009974
+ lvsat = -0.0084760193
+ lvth0 = -7.862043e-10
+ delta = 0.018814
+ wvfbsdoff = 0
+ laigc = -8.0232722e-12
+ lvfbsdoff = 0
+ rnoia = 0
+ rnoib = 0
+ acnqsmod = 0
+ fprout = 200
+ pketa = -2.6436916e-15
+ ngate = 1.7e+20
+ xrcrg1 = 12
+ xrcrg2 = 1
+ rbodymod = 0
+ ngcon = 1
+ wpclm = -6.9641486e-7
+ poxedge = 1
+ gbmin = 1e-12
+ wtvoff = 2.4243635e-10
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ keta = -0.44725926
+ binunit = 2
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = -8.778605e-11
+ capmod = 2
+ kt1l = 0
+ wku0we = 1.5e-11
+ wpdiblc2 = -6.1394667e-10
+ mobmod = 0
+ lint = 0
+ lkt1 = -9.823245e-9
+ lkt2 = -7.0749959e-9
+ lmax = 5.567e-8
+ lmin = 4.667e-8
+ a0 = -1.6354335
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 16386.797
+ cf = 8.741900000000001e-11
+ lpe0 = 6.44e-8
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.041737421
+ k3 = -2.5823
+ em = 20000000.0
+ lpeb = 0
+ ll = 0
+ lw = 0
+ u0 = 0.020918207
+ w0 = 0
+ tvoff = 0.0019328761
+ ua = 4.7595173e-10
+ ub = 8.907212200000001e-18
+ uc = 4.7837975e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 2.33e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ minv = -0.33
+ xjbvd = 1
+ xjbvs = 1
+ lua1 = 2.8472544e-16
+ lub1 = -3.7011047e-25
+ lk2we = 0.0
+ luc1 = 1.3087235e-18
+ ndep = 1e+18
+ wkvth0we = 0.0
+ lwlc = 0
+ moin = 5.5538
+ ku0we = -0.0007
+ trnqsmod = 0
+ nigc = 2.291
+ beta0 = 13.32
+ leta0 = 7.0016629000000005e-9
+ letab = 8.9813755e-9
+ ppclm = 3.4346058e-14
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ njtsswg = 6.489
+ ntox = 2.958
+ pcit = -4.1299209999999995e-17
+ pclm = 3.8611263
+ rgatemod = 0
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ tnjtsswg = 1
+ dmcgt = 0
+ ckappad = 0.6
+ phin = 0.15
+ ckappas = 0.6
+ tcjsw = 9.34e-5
+ pdiblc1 = 0
+ pdiblc2 = 0.0042244444
+ pdiblcb = 0
+ pkt1 = 4.7057745e-15
+ pkt2 = 2.4836304e-15
+ bigsd = 0.0003327
+ toxref = 3e-9
+ rbdb = 50
+ pua1 = -1.6418584e-22
+ prwb = 0
+ pub1 = 2.3001287e-31
+ prwg = 0
+ puc1 = -1.0662889e-23
+ wtvfbsdoff = 0
+ bigbacc = 0.0054401
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ wvoff = 3.9335999e-9
+ rdsw = 200
+ wvsat = -0.041964219000000004
+ kvth0we = -0.00022
+ ltvfbsdoff = 0
+ wvth0 = 3.3191681000000005e-8
+ waigc = 9.3495749e-11
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ ltvoff = -6.1656569e-12
+ lketa = 1.7473037e-8
+ xpart = 1
+ rshg = 14.1
+ pvfbsdoff = 0
+ egidl = 0.001
+ ptvfbsdoff = 0
+ lku0we = 1.8e-11
+ epsrox = 3.9
+ ijthsfwd = 0.01
+ rdsmod = 0
+ igbmod = 1
+ tnom = 25
+ toxe = 2.6300000000000002e-9
+ toxm = 2.67e-9
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ nfactor = 1
+ pbswgd = 0.8
+ pbswgs = 0.8
+ ijthsrev = 0.01
+ igcmod = 1
+ pvoff = -6.1936248e-17
+ cdscb = 0
+ cdscd = 0
+ wags = -1.0331048e-6
+ pvsat = 2.1749471e-9
+ wk2we = 0.0
+ pvth0 = -1.49270254e-15
+ wcit = 6.9580393e-10
+ drout = 0.56
+ )

.model pch_ff_32 pmos (
+ level = 54
+ tvoff = 0.0050068134
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ voffcv = -0.125
+ wpemod = 1
+ njtsswg = 6.489
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = 3.3114638e-9
+ ckappad = 0.6
+ letab = 1.8240871e-9
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.0042244444
+ pdiblcb = 0
+ keta = -0.10111506
+ ppclm = 1.7398739e-15
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = -5.51337e-11
+ kt1l = 0
+ tpbswg = 0.001
+ bigbacc = 0.0054401
+ lint = 0
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ lkt1 = -7.393592e-9
+ lkt2 = 2.2261728e-10
+ lmax = 4.667e-8
+ kvth0we = -0.00022
+ lmin = 3.6e-8
+ lpe0 = 6.44e-8
+ ijthsfwd = 0.01
+ lpeb = 0
+ ptvoff = 3.2244316e-17
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ waigsd = 1.9257033e-12
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ minv = -0.33
+ bigsd = 0.0003327
+ lua1 = -1.7116539e-16
+ lub1 = 1.5979691e-25
+ luc1 = 2.2025561e-17
+ ndep = 1e+18
+ diomod = 1
+ lwlc = 0
+ wvoff = 1.094003e-8
+ moin = 5.5538
+ ijthsrev = 0.01
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.6832999999999998e-10
+ pku0we = 0.0
+ cjswgs = 1.6832999999999998e-10
+ nigc = 2.291
+ wvsat = -0.011797954000000001
+ wvth0 = -1.1236766999999998e-8
+ waigc = 1.753535e-10
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ mjswgd = 0.95
+ mjswgs = 0.95
+ lketa = 5.1197136e-10
+ tcjswg = 0.00128
+ xpart = 1
+ ntox = 2.958
+ ppdiblc2 = 0
+ pcit = 2.2708203999999996e-16
+ pclm = 0.85281474
+ pvfbsdoff = 0
+ nfactor = 1
+ egidl = 0.001
+ phin = 0.15
+ pkt1 = 3.217758e-15
+ pkt2 = -1.2154904e-16
+ fprout = 200
+ pkvth0we = 0.0
+ rbdb = 50
+ pua1 = 5.9435365e-23
+ prwb = 0
+ pub1 = -7.9841225e-32
+ prwg = 0
+ puc1 = -3.4884574e-24
+ xrcrg1 = 12
+ xrcrg2 = 1
+ nigbacc = 10
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ rdsw = 200
+ wtvoff = -6.8770288e-10
+ vfbsdoff = 0.01
+ pvoff = -4.0525133000000003e-16
+ ags = 5.9031333
+ nigbinv = 2.171
+ cdscb = 0
+ cdscd = 0
+ cjd = 0.0012517799999999999
+ cit = 0.0020236730999999997
+ cjs = 0.0012517799999999999
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ pvsat = 6.968022699999999e-10
+ dlc = 4.0349e-9
+ wk2we = 0.0
+ pvth0 = 6.842891999999999e-16
+ k3b = 2.1176
+ dwb = 0
+ drout = 0.56
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ capmod = 2
+ paramchk = 1
+ paigc = -7.8762427e-18
+ wku0we = 1.5e-11
+ rshg = 14.1
+ voffl = 0
+ la0 = -2.1218621e-7
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0.009491273
+ mobmod = 0
+ kt1 = -0.128073887
+ kt2 = -0.09774321
+ lk2 = 3.6572258000000005e-9
+ llc = 0
+ lln = 1
+ lu0 = -2.555917e-10
+ mjd = 0.335
+ mjs = 0.335
+ lua = 4.1444844e-17
+ lub = -1.9107845e-25
+ luc = -1.4956542e-17
+ lud = 0
+ lwc = 0
+ weta0 = 7.0101382e-9
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ wetab = -5.613608e-9
+ njs = 1.02
+ pa0 = 5.0455005e-14
+ fnoimod = 1
+ nsd = 1e+20
+ pbd = 0.75
+ pat = -2.5091026e-9
+ pbs = 0.75
+ pk2 = 3.3742201e-16
+ lpclm = -1.3264792e-8
+ pu0 = 1.5059926e-16
+ eigbinv = 1.1
+ prt = 0
+ pua = 9.2877876e-24
+ pub = 4.9191362e-32
+ puc = 3.1614905e-24
+ pud = 0
+ ijthdfwd = 0.01
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 5.9585425e-9
+ ub1 = -6.9064063e-18
+ uc1 = -2.7971012e-10
+ cgidl = 1
+ tpb = 0.0016
+ wa0 = -7.0776268e-7
+ ute = -1
+ wat = 0.054757684
+ web = 6628.3
+ wec = -16935.0
+ wk2 = -3.5768953e-9
+ wlc = 0
+ wln = 1
+ wu0 = -3.0868494e-9
+ tnom = 25
+ xgl = -8.2e-9
+ xgw = 0
+ wua = -2.0394912e-16
+ wub = -1.11553208e-24
+ wuc = -7.9561907e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ toxe = 2.6300000000000002e-9
+ toxm = 2.67e-9
+ laigsd = -3.6731852e-16
+ pbswd = 0.9
+ pbsws = 0.9
+ ijthdrev = 0.01
+ cigbacc = 0.245
+ lpdiblc2 = 0
+ pdits = 0
+ wags = -1.0331048e-6
+ cigsd = 0.013281
+ tnoimod = 0
+ dvt0w = 0
+ dvt1w = 0
+ wcit = -4.7813426e-9
+ dvt2w = 0
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ a0 = 2.7407131
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = -212930.58000000002
+ cf = 8.741900000000001e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.013862232
+ k3 = -2.5823
+ em = 20000000.0
+ voff = -0.14966725
+ ll = 0
+ lw = 0
+ u0 = 0.012797793
+ w0 = 0
+ cigbinv = 0.006
+ acde = 0.5
+ ua = -1.4437109e-9
+ ub = 5.4770079e-18
+ uc = 3.1168444e-10
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 2.33e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ vsat = 140706.62
+ wint = 0
+ vth0 = -0.34311832999999997
+ wkt1 = -6.016252499999999e-8
+ wkt2 = 7.5037926e-9
+ wtvfbsdoff = 0
+ wmax = 5.374e-7
+ aigc = 0.006152944
+ wmin = 2.674e-7
+ lkvth0we = 3e-12
+ tnoia = 0
+ version = 4.5
+ tempmod = 0
+ peta0 = -3.9825789e-16
+ ltvfbsdoff = 0
+ petab = 2.3283989e-16
+ wketa = 1.3494424e-8
+ wua1 = -1.7234672e-15
+ wub1 = 2.4173164e-24
+ wuc1 = 5.6346661e-17
+ tpbsw = 0.0025
+ acnqsmod = 0
+ toxref = 3e-9
+ bigc = 0.0012521
+ aigbacc = 0.012071
+ cjswd = 4.743e-11
+ cjsws = 4.743e-11
+ wwlc = 0
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ rbodymod = 0
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.2212350000000004e-11
+ cgdo = 2.8335740000000002e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.2212350000000004e-11
+ cgso = 2.8335740000000002e-11
+ cigc = 0.15259
+ aigbinv = 0.009974
+ tvfbsdoff = 0.1
+ ptvfbsdoff = 0
+ ltvoff = -1.5678858e-10
+ scref = 1e-6
+ pigcd = 2.572
+ aigsd = 0.0063633987
+ wpdiblc2 = -6.1394667e-10
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ lku0we = 1.8e-11
+ lvoff = -1.7133213e-9
+ epsrox = 3.9
+ lvsat = -0.0031457151
+ poxedge = 1
+ lvth0 = 4.951746e-10
+ k2we = 5e-5
+ wvfbsdoff = 0
+ rdsmod = 0
+ lvfbsdoff = 0
+ delta = 0.018814
+ dsub = 0.5
+ dtox = 3.91e-10
+ laigc = 1.1545174e-11
+ igbmod = 1
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ binunit = 2
+ rnoia = 0
+ rnoib = 0
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ pbswgd = 0.8
+ wkvth0we = 0.0
+ pbswgs = 0.8
+ eta0 = 0.08799813
+ pketa = 1.5922924e-16
+ etab = -0.088479977
+ ngate = 1.7e+20
+ ngcon = 1
+ igcmod = 1
+ wpclm = -3.0982532e-8
+ trnqsmod = 0
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ paigsd = 2.0055591e-22
+ rgatemod = 0
+ tnjtsswg = 1
+ permod = 1
+ )

.model pch_ff_33 pmos (
+ level = 54
+ version = 4.5
+ pdits = 0
+ cigsd = 0.013281
+ tempmod = 0
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ tpbswg = 0.001
+ rshg = 14.1
+ aigbacc = 0.012071
+ wpdiblc2 = 3.3638075e-10
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ tnoia = 0
+ ptvoff = 0
+ aigbinv = 0.009974
+ peta0 = 2e-17
+ waigsd = 1.9846811e-12
+ wketa = -1.9384664e-9
+ tpbsw = 0.0025
+ tnom = 25
+ diomod = 1
+ cjswd = 4.743e-11
+ cjsws = 4.743e-11
+ toxe = 2.6300000000000002e-9
+ toxm = 2.67e-9
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ wkvth0we = 0.0
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.6832999999999998e-10
+ pku0we = 0.0
+ cjswgs = 1.6832999999999998e-10
+ trnqsmod = 0
+ tvfbsdoff = 0.1
+ poxedge = 1
+ mjswgd = 0.95
+ wags = 5.1942014e-9
+ mjswgs = 0.95
+ tcjswg = 0.00128
+ binunit = 2
+ scref = 1e-6
+ voff = -0.10372023
+ acde = 0.5
+ pigcd = 2.572
+ aigsd = 0.0063632583
+ rgatemod = 0
+ vsat = 108525.44
+ tnjtsswg = 1
+ wint = 0
+ vth0 = -0.34287115999999995
+ lvoff = 0
+ wkt1 = -3.0503659e-9
+ wkt2 = -7.2833333e-10
+ wmax = 2.674e-7
+ aigc = 0.0068302204
+ wmin = 1.08e-7
+ lvsat = -0.00028
+ lvth0 = 3e-10
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ delta = 0.018814
+ wua1 = -5.5326541e-17
+ wub1 = -1.0689498e-25
+ wuc1 = -1.2119467e-17
+ fprout = 200
+ rnoia = 0
+ rnoib = 0
+ bigc = 0.0012521
+ wute = -7.6523556e-8
+ xrcrg1 = 12
+ xrcrg2 = 1
+ wwlc = 0
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ ngate = 1.7e+20
+ ngcon = 1
+ cdsc = 0
+ wpclm = 7.1298978e-9
+ cgbo = 0
+ cgdl = 3.2212350000000004e-11
+ wtvoff = -7.3630015e-11
+ cgdo = 2.8335740000000002e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.2212350000000004e-11
+ cgso = 2.8335740000000002e-11
+ cigc = 0.15259
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ capmod = 2
+ wku0we = 1.5e-11
+ mobmod = 0
+ njtsswg = 6.489
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ k2we = 5e-5
+ ckappad = 0.6
+ ckappas = 0.6
+ ijthsfwd = 0.01
+ pdiblc1 = 0
+ pdiblc2 = 0.0015492917
+ dsub = 0.5
+ pdiblcb = 0
+ dtox = 3.91e-10
+ tvoff = 0.0025423547
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ eta0 = 0.10792519
+ etab = -0.13555556
+ ijthsrev = 0.01
+ ku0we = -0.0007
+ bigbacc = 0.0054401
+ beta0 = 13.32
+ leta0 = 6e-10
+ wtvfbsdoff = 0
+ kvth0we = -0.00022
+ ppclm = 0
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ dlcig = 2.5e-9
+ lintnoi = -5e-9
+ bgidl = 1834800000.0
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ ltvfbsdoff = 0
+ ppdiblc2 = 0
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ toxref = 3e-9
+ bigsd = 0.0003327
+ ptvfbsdoff = 0
+ pkvth0we = 0.0
+ wvoff = 1.4142431e-9
+ a0 = 2.5876667
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 72000
+ cf = 8.741900000000001e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.015389268
+ k3 = -2.5823
+ em = 20000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.0092771852
+ w0 = 0
+ ua = -1.9215717e-10
+ ub = 1.2747184e-18
+ uc = -1.7585185e-12
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 2.33e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ wvsat = -0.0013318206
+ nfactor = 1
+ wvth0 = -5.254371999999997e-10
+ vfbsdoff = 0.01
+ waigc = 1.6569661e-12
+ keta = 0.02482765
+ ltvoff = 0
+ jswd = 3.69e-13
+ lketa = 0
+ jsws = 3.69e-13
+ paramchk = 1
+ lcit = -2e-11
+ xpart = 1
+ pvfbsdoff = 0
+ kt1l = 0
+ lku0we = 1.8e-11
+ nigbacc = 10
+ egidl = 0.001
+ epsrox = 3.9
+ lint = 6.5375218e-9
+ lkt1 = 6e-10
+ lmax = 2.001e-5
+ lmin = 9.00077e-6
+ rdsmod = 0
+ ijthdfwd = 0.01
+ lpe0 = 6.44e-8
+ igbmod = 1
+ lpeb = 0
+ nigbinv = 2.171
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ minv = -0.33
+ pbswgd = 0.8
+ pbswgs = 0.8
+ ndep = 1e+18
+ ags = 0.89683683
+ lwlc = 0
+ igcmod = 1
+ moin = 5.5538
+ ijthdrev = 0.01
+ cjd = 0.0012517799999999999
+ cit = 5e-6
+ cjs = 0.0012517799999999999
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 1.0572421799999999e-8
+ nigc = 2.291
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ lpdiblc2 = 0
+ fnoimod = 1
+ pvoff = -2.5e-17
+ eigbinv = 1.1
+ cdscb = 0
+ cdscd = 0
+ la0 = 0
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ jsd = 1.5e-7
+ pvsat = 0
+ jss = 1.5e-7
+ lat = -0.0008
+ kt1 = -0.17197747
+ lk2 = -4e-10
+ kt2 = -0.050761111
+ wk2we = 0.0
+ pvth0 = 1.5e-16
+ llc = 0
+ lln = 1
+ lu0 = -1.2e-11
+ drout = 0.56
+ mjd = 0.335
+ mjs = 0.335
+ lub = 0
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 0
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ pk2 = 0
+ pu0 = 0
+ ntox = 2.958
+ voffl = 0
+ prt = 0
+ pub = 0
+ pcit = 1e-18
+ pud = 0
+ pclm = 1.101657
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 9.8162749e-10
+ ub1 = -3.8648101e-20
+ uc1 = 8.1681111e-11
+ tpb = 0.0016
+ weta0 = 2.4203288999999997e-9
+ permod = 1
+ wa0 = 4.8944e-8
+ wetab = 2.9133333e-9
+ ute = -0.81574074
+ phin = 0.15
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 3.9065138e-9
+ lkvth0we = 3e-12
+ lpclm = 0
+ wlc = 0
+ wln = 1
+ wu0 = 5.8460889e-11
+ xgl = -8.2e-9
+ xgw = 0
+ wua = -4.8614483e-17
+ wub = 8.106039e-27
+ wuc = 3.3309111e-18
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ cigbacc = 0.245
+ pkt1 = 5e-17
+ cgidl = 1
+ tnoimod = 0
+ acnqsmod = 0
+ voffcv = -0.125
+ wpemod = 1
+ rbdb = 50
+ prwb = 0
+ prwg = 0
+ rbpb = 50
+ rbpd = 50
+ cigbinv = 0.006
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ pbswd = 0.9
+ rbodymod = 0
+ pbsws = 0.9
+ rdsw = 200
+ )

.model pch_ff_34 pmos (
+ level = 54
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ nfactor = 1
+ ptvoff = -5.393716e-17
+ k2we = 5e-5
+ waigsd = 1.9861139e-12
+ ijthdfwd = 0.01
+ dsub = 0.5
+ dtox = 3.91e-10
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ diomod = 1
+ bigsd = 0.0003327
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.6832999999999998e-10
+ pku0we = 0.0
+ cjswgs = 1.6832999999999998e-10
+ eta0 = 0.10792519
+ wvoff = 1.3100722e-9
+ etab = -0.13555556
+ ijthdrev = 0.01
+ nigbacc = 10
+ wvsat = -0.0013318206
+ wvth0 = -6.211130999999999e-10
+ lpdiblc2 = 6.2970633e-9
+ waigc = 1.4905459e-12
+ mjswgd = 0.95
+ mjswgs = 0.95
+ tcjswg = 0.00128
+ nigbinv = 2.171
+ lketa = -5.5366519e-8
+ pvfbsdoff = 0
+ xpart = 1
+ egidl = 0.001
+ lkvth0we = 3e-12
+ fnoimod = 1
+ ags = 0.84380759
+ eigbinv = 1.1
+ fprout = 200
+ cjd = 0.0012517799999999999
+ cit = 5e-6
+ cjs = 0.0012517799999999999
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ acnqsmod = 0
+ dlc = 1.0572421799999999e-8
+ xrcrg1 = 12
+ xrcrg2 = 1
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ rbodymod = 0
+ la0 = -3.9401851e-7
+ wtvoff = -6.7630331e-11
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = -0.0008
+ kt1 = -0.17107141
+ kt2 = -0.050597496
+ lk2 = 5.1319403e-9
+ llc = 0
+ lln = 1
+ lu0 = 9.8478999e-10
+ mjd = 0.335
+ mjs = 0.335
+ lua = -7.2048384e-17
+ lub = 4.3514377e-25
+ luc = 1.4270275e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = -3.1655381e-14
+ pvoff = 9.1149624e-16
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ pk2 = 9.285497e-17
+ keta = 0.030986328
+ pu0 = 3.0504276e-17
+ prt = 0
+ cdscb = 0
+ cdscd = 0
+ pua = 2.7735079e-23
+ pub = -4.2717478e-32
+ puc = 1.20866e-25
+ pud = 0
+ cigbacc = 0.245
+ capmod = 2
+ pvsat = 0
+ rsh = 15.2
+ wk2we = 0.0
+ tcj = 0.000832
+ ua1 = 8.0734953e-10
+ pvth0 = 1.01012639e-15
+ ub1 = 2.6826436e-19
+ uc1 = 8.9789043e-11
+ drout = 0.56
+ lags = 4.7673289e-7
+ wku0we = 1.5e-11
+ tpb = 0.0016
+ wa0 = 5.2465177e-8
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ ute = -0.817454
+ paigc = 1.4961177e-18
+ lcit = -2e-11
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 3.8961851e-9
+ tnoimod = 0
+ mobmod = 0
+ wlc = 0
+ wln = 1
+ wu0 = 5.5067755e-11
+ xgl = -8.2e-9
+ xgw = 0
+ kt1l = 0
+ wua = -5.1699586e-17
+ wub = 1.2857705e-26
+ wuc = 3.3174666e-18
+ wud = 0
+ voffl = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ wpdiblc2 = 3.5925269e-10
+ cigbinv = 0.006
+ weta0 = 2.4203288999999997e-9
+ wetab = 2.9133333e-9
+ lint = 6.5375218e-9
+ lpclm = 0
+ lkt1 = -7.5454893e-9
+ lkt2 = -1.4709041e-9
+ lmax = 9.00077e-6
+ lmin = 9.0075e-7
+ lpe0 = 6.44e-8
+ cgidl = 1
+ lpeb = 0
+ version = 4.5
+ tempmod = 0
+ minv = -0.33
+ wtvfbsdoff = 0
+ laigsd = -1.8524358e-14
+ lua1 = 1.5667589e-15
+ lub1 = -2.759143e-24
+ luc1 = -7.2890309e-17
+ ndep = 1e+18
+ wkvth0we = 0.0
+ lute = 1.5402209e-8
+ lwlc = 0
+ pbswd = 0.9
+ pbsws = 0.9
+ moin = 5.5538
+ aigbacc = 0.012071
+ ltvfbsdoff = 0
+ trnqsmod = 0
+ nigc = 2.291
+ pdits = 0
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ noff = 2.2684
+ cigsd = 0.013281
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ aigbinv = 0.009974
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ pags = -1.92428e-14
+ ntox = 2.958
+ pcit = 1e-18
+ rgatemod = 0
+ pclm = 1.101657
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ ptvfbsdoff = 0
+ tnjtsswg = 1
+ phin = 0.15
+ tnoia = 0
+ pkt1 = -2.7622214e-15
+ pkt2 = 2.4239149e-16
+ peta0 = 2e-17
+ toxref = 3e-9
+ wketa = -2.0595747e-9
+ poxedge = 1
+ tpbsw = 0.0025
+ cjswd = 4.743e-11
+ cjsws = 4.743e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ rbdb = 50
+ pua1 = -1.1776704e-22
+ binunit = 2
+ prwb = 0
+ pub1 = 2.7996299e-31
+ prwg = 0
+ puc1 = 9.811687e-24
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ pute = 1.5923616e-14
+ rdsw = 200
+ tvfbsdoff = 0.1
+ ltvoff = -3.3500511e-10
+ scref = 1e-6
+ pigcd = 2.572
+ rshg = 14.1
+ aigsd = 0.0063632604
+ lku0we = 1.8e-11
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ epsrox = 3.9
+ lvoff = -2.4480721e-8
+ a0 = 2.6314952
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ rdsmod = 0
+ wvfbsdoff = 0
+ at = 72000
+ cf = 8.741900000000001e-11
+ lvsat = -0.00028
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.016004612
+ k3 = -2.5823
+ em = 20000000.0
+ lvfbsdoff = 0
+ lvth0 = -1.3566904e-8
+ igbmod = 1
+ ll = 0
+ lw = 0
+ u0 = 0.0091663075
+ w0 = 0
+ ua = -1.8414289e-10
+ ub = 1.2263153e-18
+ uc = -3.3458683e-12
+ ud = 0
+ ijthsfwd = 0.01
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 2.33e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ delta = 0.018814
+ laigc = -5.3027874e-11
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ rnoia = 0
+ rnoib = 0
+ pbswgd = 0.8
+ pbswgs = 0.8
+ tnom = 25
+ toxe = 2.6300000000000002e-9
+ toxm = 2.67e-9
+ igcmod = 1
+ pketa = 1.0887638e-15
+ ngate = 1.7e+20
+ ngcon = 1
+ ijthsrev = 0.01
+ wpclm = 7.1298978e-9
+ njtsswg = 6.489
+ gbmin = 1e-12
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ wags = 7.3346686e-9
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.00084883969
+ pdiblcb = 0
+ paigsd = -1.2880862e-20
+ voff = -0.10099712
+ acde = 0.5
+ ppdiblc2 = -2.0561872e-16
+ vsat = 108525.44
+ wint = 0
+ permod = 1
+ vth0 = -0.34132868000000005
+ wkt1 = -2.7375492e-9
+ wkt2 = -7.5529568e-10
+ wmax = 2.674e-7
+ aigc = 0.0068361189
+ wmin = 1.08e-7
+ bigbacc = 0.0054401
+ tvoff = 0.0025796189
+ kvth0we = -0.00022
+ wua1 = -4.222676e-17
+ wub1 = -1.3803658e-25
+ wuc1 = -1.3210867e-17
+ xjbvd = 1
+ xjbvs = 1
+ voffcv = -0.125
+ wpemod = 1
+ lk2we = 0.0
+ lintnoi = -5e-9
+ bigc = 0.0012521
+ wute = -7.8294814e-8
+ bigbinv = 0.00149
+ pkvth0we = 0.0
+ wwlc = 0
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ cdsc = 0
+ ku0we = -0.0007
+ cgbo = 0
+ cgdl = 3.2212350000000004e-11
+ cgdo = 2.8335740000000002e-11
+ xtid = 3
+ xtis = 3
+ beta0 = 13.32
+ leta0 = 6e-10
+ vfbsdoff = 0.01
+ cgsl = 3.2212350000000004e-11
+ cgso = 2.8335740000000002e-11
+ cigc = 0.15259
+ ppclm = 0
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ paramchk = 1
+ tpbswg = 0.001
+ )

.model pch_ff_35 pmos (
+ level = 54
+ cjsws = 4.743e-11
+ cjswgd = 1.6832999999999998e-10
+ pku0we = 0.0
+ cjswgs = 1.6832999999999998e-10
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ ndep = 1e+18
+ lute = -1.0958354e-8
+ lwlc = 0
+ moin = 5.5538
+ ijthsrev = 0.01
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ tvfbsdoff = 0.1
+ nigc = 2.291
+ mjswgd = 0.95
+ mjswgs = 0.95
+ tcjswg = 0.00128
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ scref = 1e-6
+ pags = 1.1742809e-13
+ ppdiblc2 = -6.1367245e-16
+ pigcd = 2.572
+ ntox = 2.958
+ aigsd = 0.0063632396
+ pcit = 1e-18
+ pclm = 1.101657
+ lvoff = -2.4340257e-9
+ phin = 0.15
+ wvfbsdoff = 0
+ njtsswg = 6.489
+ lvfbsdoff = 0
+ lvsat = -0.00028
+ lvth0 = 2.7200595e-10
+ pkt1 = 5.797333199999999e-15
+ pkt2 = -5.7270183e-16
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ delta = 0.018814
+ fprout = 200
+ laigc = -3.3884553e-11
+ xrcrg1 = 12
+ xrcrg2 = 1
+ ckappad = 0.6
+ ckappas = 0.6
+ rnoia = 0
+ rnoib = 0
+ pdiblc1 = 0
+ pdiblc2 = 0.0027845581
+ pdiblcb = 0
+ pkvth0we = 0.0
+ rbdb = 50
+ pua1 = -9.8048843e-24
+ prwb = 0
+ pub1 = -2.3189739e-32
+ prwg = 0
+ puc1 = -4.5795492e-24
+ pketa = -3.0075994e-15
+ rbpb = 50
+ rbpd = 50
+ ngate = 1.7e+20
+ rbps = 50
+ rbsb = 50
+ wtvoff = -2.2790108e-10
+ pvag = 2.1
+ pute = -9.4649237e-15
+ ngcon = 1
+ wpclm = 7.1298978e-9
+ rdsw = 200
+ vfbsdoff = 0.01
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ bigbacc = 0.0054401
+ capmod = 2
+ wku0we = 1.5e-11
+ kvth0we = -0.00022
+ mobmod = 0
+ paramchk = 1
+ lintnoi = -5e-9
+ rshg = 14.1
+ bigbinv = 0.00149
+ wtvfbsdoff = 0
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ ltvfbsdoff = 0
+ ijthdfwd = 0.01
+ tvoff = 0.0027416725
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ tnom = 25
+ toxe = 2.6300000000000002e-9
+ toxm = 2.67e-9
+ ijthdrev = 0.01
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = 6e-10
+ lpdiblc2 = 4.574275e-9
+ ptvfbsdoff = 0
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ nfactor = 1
+ ppclm = 0
+ wags = -1.4622812e-7
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ voff = -0.12576869
+ acde = 0.5
+ vsat = 108525.44
+ wint = 0
+ vth0 = -0.35687802
+ wkt1 = -1.2355026e-8
+ wkt2 = 1.605395e-10
+ dmcgt = 0
+ wmax = 2.674e-7
+ tcjsw = 9.34e-5
+ lkvth0we = 3e-12
+ aigc = 0.0068146096
+ wmin = 1.08e-7
+ nigbacc = 10
+ toxref = 3e-9
+ wua1 = -1.6353255e-16
+ wub1 = 2.0258446e-25
+ wuc1 = 2.9590615e-18
+ acnqsmod = 0
+ bigsd = 0.0003327
+ bigc = 0.0012521
+ wute = -4.9768365e-8
+ nigbinv = 2.171
+ wwlc = 0
+ wvoff = 3.4766421e-9
+ rbodymod = 0
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.2212350000000004e-11
+ cgdo = 2.8335740000000002e-11
+ wvsat = -0.0013318206
+ xtid = 3
+ xtis = 3
+ wvth0 = 1.4834680000000002e-10
+ ltvoff = -4.7923289e-10
+ cgsl = 3.2212350000000004e-11
+ cgso = 2.8335740000000002e-11
+ cigc = 0.15259
+ waigc = 2.7104678e-12
+ fnoimod = 1
+ eigbinv = 1.1
+ pvfbsdoff = 0
+ lketa = 4.197898e-9
+ xpart = 1
+ lku0we = 1.8e-11
+ epsrox = 3.9
+ wpdiblc2 = 8.1773971e-10
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ ags = 1.7348065
+ dmdg = 0
+ egidl = 0.001
+ cjd = 0.0012517799999999999
+ rdsmod = 0
+ cit = -8.7888889e-5
+ cjs = 0.0012517799999999999
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 1.0572421799999999e-8
+ igbmod = 1
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ k2we = 5e-5
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ dsub = 0.5
+ dtox = 3.91e-10
+ pbswgd = 0.8
+ la0 = -1.044589e-6
+ cigbacc = 0.245
+ pbswgs = 0.8
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = -0.0008
+ kt1 = -0.11040563
+ kt2 = -0.048714998
+ lk2 = 2.6890726e-9
+ llc = 0
+ lln = 1
+ lu0 = -1.8292817999999999e-9
+ mjd = 0.335
+ mjs = 0.335
+ lua = -6.2776752e-16
+ lub = 4.4518935e-25
+ luc = 5.1177769e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ igcmod = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 1.0817056e-13
+ wkvth0we = 0.0
+ nsd = 1e+20
+ pbd = 0.75
+ tnoimod = 0
+ pat = 0
+ pbs = 0.75
+ pk2 = -1.5480351e-16
+ eta0 = 0.10792519
+ etab = -0.13555556
+ pu0 = 1.5955157e-16
+ prt = 0
+ pua = 4.4574845e-23
+ pub = -2.7161351e-32
+ puc = -4.8372521e-24
+ pud = 0
+ rsh = 15.2
+ trnqsmod = 0
+ tcj = 0.000832
+ ua1 = 2.771768e-9
+ ub1 = -3.1924567e-18
+ uc1 = -6.2120134e-12
+ cigbinv = 0.006
+ tpb = 0.0016
+ wa0 = -1.0464262e-7
+ ute = -0.78783539
+ pvoff = -1.01675093e-15
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 4.174453e-9
+ wlc = 0
+ wln = 1
+ wu0 = -8.9929205e-11
+ xgl = -8.2e-9
+ xgw = 0
+ wua = -7.0620672e-17
+ wub = -4.621089e-27
+ wuc = 8.8883858e-18
+ wud = 0
+ cdscb = 0
+ cdscd = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ pvsat = 0
+ a0 = 3.3624733
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ wk2we = 0.0
+ pvth0 = 3.2530712e-16
+ at = 72000
+ cf = 8.741900000000001e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.013259817
+ k3 = -2.5823
+ em = 20000000.0
+ drout = 0.56
+ version = 4.5
+ ll = 0
+ lw = 0
+ u0 = 0.012328186
+ w0 = 0
+ ua = 4.4026063e-10
+ ub = 1.2150282e-18
+ uc = -4.4814963e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 2.33e-9
+ ww = 0
+ paigc = 4.1038726e-19
+ xw = 8.600000000000001e-9
+ tempmod = 0
+ voffl = 0
+ rgatemod = 0
+ permod = 1
+ tnjtsswg = 1
+ weta0 = 2.4203288999999997e-9
+ wetab = 2.9133333e-9
+ aigbacc = 0.012071
+ lpclm = 0
+ cgidl = 1
+ voffcv = -0.125
+ wpemod = 1
+ aigbinv = 0.009974
+ pbswd = 0.9
+ pbsws = 0.9
+ keta = -0.035939983
+ pdits = 0
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ lags = -3.1625612e-7
+ tpbswg = 0.001
+ poxedge = 1
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 6.2671111e-11
+ kt1l = 0
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ binunit = 2
+ lint = 6.5375218e-9
+ ptvoff = 8.8703803e-17
+ lkt1 = -6.1538035e-8
+ lkt2 = -3.1463267e-9
+ tnoia = 0
+ lmax = 9.0075e-7
+ waigsd = 1.9716411e-12
+ lmin = 4.5075e-7
+ ijthsfwd = 0.01
+ peta0 = 2e-17
+ lpe0 = 6.44e-8
+ lpeb = 0
+ wketa = 2.5430806e-9
+ diomod = 1
+ tpbsw = 0.0025
+ minv = -0.33
+ lua1 = -1.8157361e-16
+ lub1 = 3.2089876e-25
+ luc1 = 1.2550631e-17
+ pditsd = 0
+ cjswd = 4.743e-11
+ pditsl = 0
+ )

.model pch_ff_36 pmos (
+ level = 54
+ ags = 0.79842724
+ pvfbsdoff = 0
+ wcit = 5.8162887e-11
+ lketa = -1.0850486e-8
+ cigbacc = 0.245
+ cjd = 0.0012517799999999999
+ cit = -0.00049977211
+ cjs = 0.0012517799999999999
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ voff = -0.11894985
+ xpart = 1
+ dlc = 1.38228675e-8
+ k3b = 2.1176
+ acde = 0.5
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ rgatemod = 0
+ tnjtsswg = 1
+ vsat = 108525.44
+ tnoimod = 0
+ wint = 0
+ vth0 = -0.36350625999999997
+ egidl = 0.001
+ wkt1 = 8.365112e-10
+ wkt2 = -1.4765978e-9
+ la0 = -3.2362015e-7
+ wmax = 2.674e-7
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = -0.0008
+ aigc = 0.0068096243
+ wmin = 1.08e-7
+ kt1 = -0.25321364
+ kt2 = -0.04359324
+ lk2 = -7.427309000000001e-10
+ llc = -1.18e-13
+ lln = 0.7
+ cigbinv = 0.006
+ lu0 = -4.6259608e-10
+ mjd = 0.335
+ mjs = 0.335
+ lua = -1.7021816e-16
+ lub = 1.0550853e-25
+ luc = -1.2975077e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ fprout = 200
+ njs = 1.02
+ pa0 = -3.1370244e-14
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ pk2 = 1.4083403e-16
+ xrcrg1 = 12
+ xrcrg2 = 1
+ pu0 = -1.3937081e-17
+ prt = 0
+ pua = 4.7117679e-24
+ pub = -8.7289665e-33
+ puc = -3.0945045e-25
+ pud = 0
+ wua1 = -2.3000717e-16
+ wub1 = 1.2114667e-25
+ wuc1 = -1.9684753e-17
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 2.6350858e-9
+ ub1 = -2.2549964e-18
+ uc1 = 3.1191962e-11
+ bigc = 0.0012521
+ wute = -1.1762912e-7
+ version = 4.5
+ tpb = 0.0016
+ wa0 = 2.1249557e-7
+ wwlc = 0
+ ute = -0.71022675
+ wtvoff = -1.1036076e-10
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 3.5025496e-9
+ tempmod = 0
+ wlc = 0
+ wln = 1
+ wu0 = 3.0436319e-10
+ xgl = -8.2e-9
+ xgw = 0
+ wua = 1.9977231e-17
+ wub = -4.6512873e-26
+ wuc = -1.4020724e-18
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.2212350000000004e-11
+ cgdo = 2.8335740000000002e-11
+ xtid = 3
+ xtis = 3
+ wtvfbsdoff = 0
+ aigbacc = 0.012071
+ cgsl = 3.2212350000000004e-11
+ cgso = 2.8335740000000002e-11
+ cigc = 0.15259
+ pvoff = 7.0942711e-17
+ capmod = 2
+ cdscb = 0
+ cdscd = 0
+ wku0we = 1.5e-11
+ pvsat = 0
+ wk2we = 0.0
+ pvth0 = -8.393785000000001e-17
+ ltvfbsdoff = 0
+ drout = 0.56
+ mobmod = 0
+ paigc = -1.759214e-19
+ aigbinv = 0.009974
+ voffl = 0
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ weta0 = 2.4203288999999997e-9
+ wetab = 2.9133333e-9
+ lpclm = 0
+ k2we = 5e-5
+ ijthsfwd = 0.01
+ cgidl = 1
+ dsub = 0.5
+ ptvfbsdoff = 0
+ dtox = 3.91e-10
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ poxedge = 1
+ eta0 = 0.10792519
+ pbswd = 0.9
+ etab = -0.13555556
+ pbsws = 0.9
+ ijthsrev = 0.01
+ binunit = 2
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ pdits = 0
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ ppdiblc2 = 9.2177422e-17
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ tnoia = 0
+ toxref = 3e-9
+ peta0 = 2e-17
+ wketa = -1.9938172e-9
+ tpbsw = 0.0025
+ cjswd = 4.743e-11
+ cjsws = 4.743e-11
+ pkvth0we = 0.0
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ tvfbsdoff = 0.1
+ ltvoff = -1.9203223e-10
+ vfbsdoff = 0.01
+ njtsswg = 6.489
+ keta = -0.0017391106
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ lags = 9.5750741e-8
+ lku0we = 1.8e-11
+ paramchk = 1
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ scref = 1e-6
+ ckappad = 0.6
+ ckappas = 0.6
+ lcit = 2.4389973e-10
+ pdiblc1 = 0
+ pdiblc2 = 0.016049816
+ epsrox = 3.9
+ pdiblcb = 0
+ pigcd = 2.572
+ kt1l = 0
+ aigsd = 0.0063632396
+ rdsmod = 0
+ lvoff = -5.4343156e-9
+ wvfbsdoff = 0
+ lint = 9.7879675e-9
+ igbmod = 1
+ lvfbsdoff = 0
+ lkt1 = 1.297866e-9
+ lkt2 = -5.3999005e-9
+ lvsat = -0.00028
+ lmax = 4.5075e-7
+ lvth0 = 3.1884329e-9
+ lmin = 2.1744e-7
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ ijthdfwd = 0.01
+ lpe0 = 6.44e-8
+ delta = 0.018814
+ bigbacc = 0.0054401
+ lpeb = 0
+ pbswgd = 0.8
+ laigc = -3.1691048e-11
+ pbswgs = 0.8
+ rnoia = 0
+ rnoib = 0
+ minv = -0.33
+ igcmod = 1
+ lua1 = -1.2143343e-16
+ lub1 = -9.158653e-26
+ luc1 = -3.907118e-18
+ kvth0we = -0.00022
+ ndep = 1e+18
+ lute = -4.5106156e-8
+ pketa = -1.0113644e-15
+ ngate = 1.7e+20
+ lwlc = 0
+ lintnoi = -5e-9
+ moin = 5.5538
+ ijthdrev = 0.01
+ ngcon = 1
+ bigbinv = 0.00149
+ wpclm = 7.1298978e-9
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ nigc = 2.291
+ lpdiblc2 = -1.262443e-9
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ pags = 5.2660461e-14
+ permod = 1
+ ntox = 2.958
+ pcit = -2.459167e-17
+ pclm = 1.101657
+ phin = 0.15
+ lkvth0we = 3e-12
+ pkt1 = -7.047500000000005e-18
+ pkt2 = 1.4763857e-16
+ voffcv = -0.125
+ wpemod = 1
+ tvoff = 0.0020889601
+ nfactor = 1
+ xjbvd = 1
+ acnqsmod = 0
+ xjbvs = 1
+ lk2we = 0.0
+ a0 = 1.7239078
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ rbdb = 50
+ pua1 = 1.9443948e-23
+ prwb = 0
+ pub1 = 1.2643651e-32
+ prwg = 0
+ at = 72000
+ puc1 = 5.3837292e-24
+ cf = 8.741900000000001e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.0054602636
+ k3 = -2.5823
+ em = 20000000.0
+ rbpb = 50
+ rbpd = 50
+ ll = -1.18e-13
+ lw = 0
+ rbps = 50
+ u0 = 0.009222082
+ rbsb = 50
+ pvag = 2.1
+ w0 = 0
+ rbodymod = 0
+ ua = -5.9962427e-10
+ ub = 1.98703e-18
+ uc = 1.0098696e-10
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 2.33e-9
+ ww = 0
+ pute = 2.0393808e-14
+ xw = 8.600000000000001e-9
+ rdsw = 200
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = 6e-10
+ nigbacc = 10
+ ppclm = 0
+ tpbswg = 0.001
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ rshg = 14.1
+ nigbinv = 2.171
+ wpdiblc2 = -7.8646151e-10
+ ptvoff = 3.6984079e-17
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ waigsd = 1.9716411e-12
+ diomod = 1
+ fnoimod = 1
+ pditsd = 0
+ pditsl = 0
+ bigsd = 0.0003327
+ cjswgd = 1.6832999999999998e-10
+ pku0we = 0.0
+ tnom = 25
+ cjswgs = 1.6832999999999998e-10
+ eigbinv = 1.1
+ toxe = 2.6300000000000002e-9
+ toxm = 2.67e-9
+ wkvth0we = 0.0
+ wvoff = 1.0046111e-9
+ trnqsmod = 0
+ wvsat = -0.0013318206
+ mjswgd = 0.95
+ wvth0 = 1.0784490000000002e-9
+ mjswgs = 0.95
+ tcjswg = 0.00128
+ waigc = 4.0429874e-12
+ wags = 9.7102189e-10
+ )

.model pch_ff_37 pmos (
+ level = 54
+ fprout = 200
+ lvth0 = 5.8274905e-9
+ xrcrg1 = 12
+ xrcrg2 = 1
+ delta = 0.018814
+ wtvfbsdoff = 0
+ laigc = -4.357169e-12
+ rnoia = 0
+ rnoib = 0
+ acnqsmod = 0
+ wtvoff = 1.2048366e-10
+ ltvfbsdoff = 0
+ pketa = 4.1278959e-16
+ ngate = 1.7e+20
+ rbodymod = 0
+ ngcon = 1
+ wpclm = 6.8691006e-8
+ capmod = 2
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ wku0we = 1.5e-11
+ keta = -0.058692164
+ mobmod = 0
+ nfactor = 1
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 5.2914770000000015e-12
+ ptvfbsdoff = 0
+ kt1l = 0
+ wpdiblc2 = -7.28246e-10
+ lint = 9.7879675e-9
+ lkt1 = -4.0770694e-9
+ lkt2 = -3.7791597e-9
+ lmax = 2.1744e-7
+ lmin = 9.167e-8
+ lpe0 = 6.44e-8
+ nigbacc = 10
+ lpeb = 0
+ tvoff = 0.0011827459
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ minv = -0.33
+ lua1 = -2.1218464e-16
+ lub1 = 2.7818737e-25
+ luc1 = 2.2554944e-17
+ ndep = 1e+18
+ wkvth0we = 0.0
+ lute = 1.5508066e-9
+ lwlc = 0
+ moin = 5.5538
+ nigbinv = 2.171
+ ku0we = -0.0007
+ trnqsmod = 0
+ beta0 = 13.32
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ nigc = 2.291
+ leta0 = 6e-10
+ ppclm = -1.2989269e-14
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ fnoimod = 1
+ eigbinv = 1.1
+ ntox = 2.958
+ rgatemod = 0
+ pcit = 1.2214196e-17
+ pclm = 0.85425247
+ tnjtsswg = 1
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ phin = 0.15
+ toxref = 3e-9
+ pkt1 = -1.8173360000000001e-16
+ pkt2 = 3.7767926e-16
+ bigsd = 0.0003327
+ cigbacc = 0.245
+ rbdb = 50
+ pua1 = 2.6827919e-23
+ prwb = 0
+ pub1 = -3.4278711e-32
+ prwg = 0
+ puc1 = -2.7535024e-24
+ wvoff = 8.5374562e-10
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ pute = -4.2802262e-16
+ ltvoff = -8.1627e-13
+ rdsw = 200
+ tnoimod = 0
+ wvsat = -0.00089129698
+ ags = 1.2522222
+ wvth0 = 4.9052000000000173e-11
+ cjd = 0.0012517799999999999
+ cit = 0.00063107268
+ cjs = 0.0012517799999999999
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 1.38228675e-8
+ waigc = 1.4660694e-11
+ k3b = 2.1176
+ cigbinv = 0.006
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ pvfbsdoff = 0
+ lku0we = 1.8e-11
+ lketa = 1.1666086e-9
+ epsrox = 3.9
+ la0 = 6.219346e-9
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = -0.0083443287
+ xpart = 1
+ kt1 = -0.22773883
+ kt2 = -0.051274476
+ lk2 = 3.2711471e-9
+ llc = -1.18e-13
+ lln = 0.7
+ lu0 = -1.7514862000000002e-10
+ mjd = 0.335
+ version = 4.5
+ mjs = 0.335
+ lua = 1.3101868e-17
+ lub = -8.7271368e-26
+ luc = -1.2812174e-17
+ lud = 0
+ rshg = 14.1
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = -2.0637395e-14
+ rdsmod = 0
+ nsd = 1e+20
+ pbd = 0.75
+ tempmod = 0
+ pat = -5.0045721e-10
+ pbs = 0.75
+ pk2 = 4.0368065e-17
+ egidl = 0.001
+ igbmod = 1
+ pu0 = -5.2679707e-18
+ prt = 0
+ pua = -4.0286539e-24
+ pub = 7.5106005e-33
+ puc = 1.4358513e-24
+ pud = 0
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 3.0651863e-9
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ ub1 = -4.0074881e-18
+ uc1 = -9.4220652e-11
+ tpb = 0.0016
+ aigbacc = 0.012071
+ wa0 = 1.6162969e-7
+ pbswgd = 0.8
+ pbswgs = 0.8
+ ute = -0.93134979
+ ijthsfwd = 0.01
+ wat = 0.0023718351
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 3.9786916e-9
+ wlc = 0
+ wln = 1
+ wu0 = 2.6327735e-10
+ xgl = -8.2e-9
+ xgw = 0
+ wua = 6.1401032e-17
+ wub = -1.2347765e-25
+ wuc = -9.6736445e-18
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ igcmod = 1
+ tnom = 25
+ toxe = 2.6300000000000002e-9
+ toxm = 2.67e-9
+ aigbinv = 0.009974
+ ijthsrev = 0.01
+ pvoff = 1.0277532000000001e-16
+ cdscb = 0
+ cdscd = 0
+ pvsat = -9.2948987e-11
+ wags = 2.5054667e-7
+ wk2we = 0.0
+ pvth0 = 1.3326490799999998e-16
+ drout = 0.56
+ wcit = -1.162725e-10
+ paigc = -2.4162575e-18
+ permod = 1
+ voff = -0.1339517
+ acde = 0.5
+ ppdiblc2 = 7.9894307e-17
+ voffl = 0
+ poxedge = 1
+ vsat = 106518.57
+ wint = 0
+ vth0 = -0.37601365
+ weta0 = 2.4203288999999997e-9
+ wetab = 2.9133333e-9
+ wkt1 = 1.664079e-9
+ wkt2 = -2.566838e-9
+ wmax = 2.674e-7
+ lpclm = 5.2201277e-8
+ binunit = 2
+ aigc = 0.0066800799
+ wmin = 1.08e-7
+ voffcv = -0.125
+ wpemod = 1
+ cgidl = 1
+ wua1 = -2.6500229e-16
+ wub1 = 3.4352994e-25
+ wuc1 = 1.8880326e-17
+ bigc = 0.0012521
+ wute = -1.8947457e-8
+ pkvth0we = 0.0
+ wwlc = 0
+ pbswd = 0.9
+ pbsws = 0.9
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.2212350000000004e-11
+ cgdo = 2.8335740000000002e-11
+ xtid = 3
+ xtis = 3
+ vfbsdoff = 0.01
+ cgsl = 3.2212350000000004e-11
+ cgso = 2.8335740000000002e-11
+ cigc = 0.15259
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ pdits = 0
+ tpbswg = 0.001
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ paramchk = 1
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ ptvoff = -1.1725409e-17
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ a0 = 0.16068118
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ waigsd = 1.9716411e-12
+ at = 107755.11
+ cf = 8.741900000000001e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.024483382
+ k3 = -2.5823
+ em = 20000000.0
+ ll = -1.18e-13
+ lw = 0
+ u0 = 0.0078597718
+ tnoia = 0
+ w0 = 0
+ ua = -1.4684396e-9
+ ub = 2.9006788e-18
+ uc = 1.0021491e-10
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 2.33e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ diomod = 1
+ k2we = 5e-5
+ ijthdfwd = 0.01
+ peta0 = 2e-17
+ njtsswg = 6.489
+ dsub = 0.5
+ dtox = 3.91e-10
+ wketa = -8.743362e-9
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.6832999999999998e-10
+ pku0we = 0.0
+ cjswgs = 1.6832999999999998e-10
+ tpbsw = 0.0025
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ cjswd = 4.743e-11
+ cjsws = 4.743e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.01690182
+ eta0 = 0.10792519
+ pdiblcb = 0
+ etab = -0.13555556
+ tvfbsdoff = 0.1
+ ijthdrev = 0.01
+ mjswgd = 0.95
+ mjswgs = 0.95
+ lpdiblc2 = -1.4422174e-9
+ tcjswg = 0.00128
+ bigbacc = 0.0054401
+ scref = 1e-6
+ pigcd = 2.572
+ aigsd = 0.0063632396
+ kvth0we = -0.00022
+ wvfbsdoff = 0
+ lvoff = -2.268926e-9
+ lintnoi = -5e-9
+ lvfbsdoff = 0
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ lkvth0we = 3e-12
+ lvsat = 0.00014343719
+ )

.model pch_ff_38 pmos (
+ level = 54
+ poxedge = 1
+ ptvfbsdoff = 0
+ rdsw = 200
+ capmod = 2
+ vfbsdoff = 0.01
+ wku0we = 1.5e-11
+ pvoff = -1.6873466999999998e-16
+ binunit = 2
+ cdscb = 0
+ cdscd = 0
+ mobmod = 0
+ pvsat = 1.729604e-10
+ wk2we = 0.0
+ pvth0 = 8.910713399999999e-17
+ drout = 0.56
+ paramchk = 1
+ paigc = -1.1563004e-18
+ voffl = 0
+ rshg = 14.1
+ weta0 = 1.3237501e-8
+ wetab = 4.1458967e-9
+ lpclm = -1.0127779e-7
+ ijthdfwd = 0.01
+ jtsswgd = 1.75e-7
+ cgidl = 1
+ jtsswgs = 1.75e-7
+ tnom = 25
+ toxe = 2.6300000000000002e-9
+ toxm = 2.67e-9
+ pbswd = 0.9
+ pbsws = 0.9
+ ijthdrev = 0.01
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ lpdiblc2 = -1.4113545e-11
+ pdits = 0
+ cigsd = 0.013281
+ wags = 2.5054667e-7
+ dvt0w = 0
+ dvt1w = 0
+ njtsswg = 6.489
+ dvt2w = 0
+ wcit = 4.14692744e-10
+ xtsswgd = 0.32
+ voff = -0.14478455
+ xtsswgs = 0.32
+ acde = 0.5
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ ckappad = 0.6
+ ckappas = 0.6
+ vsat = 137363.5
+ wint = 0
+ pdiblc1 = 0
+ pdiblc2 = 0.0017092259
+ vth0 = -0.31895262
+ pdiblcb = 0
+ wkt1 = -1.350742e-8
+ wkt2 = 1.8825744e-9
+ toxref = 3e-9
+ wmax = 2.674e-7
+ lkvth0we = 3e-12
+ aigc = 0.0067219883
+ wmin = 1.08e-7
+ tnoia = 0
+ peta0 = -9.968142000000002e-16
+ petab = -1.1586096e-16
+ wketa = -6.6698086e-9
+ wua1 = 1.6631395e-16
+ wub1 = -2.121384e-25
+ wuc1 = 2.5860689e-17
+ tpbsw = 0.0025
+ acnqsmod = 0
+ bigbacc = 0.0054401
+ cjswd = 4.743e-11
+ bigc = 0.0012521
+ cjsws = 4.743e-11
+ wute = -6.1363432e-8
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ wwlc = 0
+ tvfbsdoff = 0.1
+ ltvoff = 3.7319947e-11
+ rbodymod = 0
+ kvth0we = -0.00022
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.2212350000000004e-11
+ cgdo = 2.8335740000000002e-11
+ xtid = 3
+ xtis = 3
+ lintnoi = -5e-9
+ cgsl = 3.2212350000000004e-11
+ cgso = 2.8335740000000002e-11
+ bigbinv = 0.00149
+ cigc = 0.15259
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ lku0we = 1.8e-11
+ epsrox = 3.9
+ scref = 1e-6
+ pigcd = 2.572
+ aigsd = 0.0063632396
+ rdsmod = 0
+ wpdiblc2 = 8.0253658e-11
+ igbmod = 1
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ lvoff = -1.2506377e-9
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ lvsat = -0.0027559865
+ pbswgd = 0.8
+ pbswgs = 0.8
+ lvth0 = 4.6375330000000005e-10
+ k2we = 5e-5
+ delta = 0.018814
+ laigc = -8.2965642e-12
+ dsub = 0.5
+ igcmod = 1
+ dtox = 3.91e-10
+ rnoia = 0
+ rnoib = 0
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ nfactor = 1
+ wkvth0we = 0.0
+ pketa = 2.1787556e-16
+ ngate = 1.7e+20
+ eta0 = 0.024468866
+ etab = -0.22797789
+ ngcon = 1
+ wpclm = -1.6917696e-7
+ trnqsmod = 0
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ nigbacc = 10
+ permod = 1
+ rgatemod = 0
+ tnjtsswg = 1
+ nigbinv = 2.171
+ voffcv = -0.125
+ wpemod = 1
+ tvoff = 0.00077704148
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ fnoimod = 1
+ eigbinv = 1.1
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = 8.444894e-9
+ letab = 8.6876992e-9
+ tpbswg = 0.001
+ ppclm = 9.3703198e-15
+ keta = -0.049241031
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 1.9424599e-10
+ kt1l = 0
+ ptvoff = 1.952106e-17
+ cigbacc = 0.245
+ waigsd = 1.9716411e-12
+ dmcgt = 0
+ lint = 0
+ tcjsw = 9.34e-5
+ tnoimod = 0
+ lkt1 = -5.994607400000001e-9
+ lkt2 = 9.2375447e-10
+ diomod = 1
+ lmax = 9.167e-8
+ lmin = 5.567e-8
+ ijthsfwd = 0.01
+ lpe0 = 6.44e-8
+ pditsd = 0
+ pditsl = 0
+ lpeb = 0
+ cigbinv = 0.006
+ cjswgd = 1.6832999999999998e-10
+ pku0we = 0.0
+ cjswgs = 1.6832999999999998e-10
+ bigsd = 0.0003327
+ minv = -0.33
+ ags = 1.2522222
+ lua1 = 1.5814311e-16
+ lub1 = -2.3663254e-25
+ luc1 = 3.1466117e-17
+ cjd = 0.0012517799999999999
+ cit = -0.0013790818100000001
+ cjs = 0.0012517799999999999
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ ndep = 1e+18
+ bvs = 8.2
+ lute = -1.2895214e-8
+ dlc = 4.0349e-9
+ wvoff = 3.7421498e-9
+ k3b = 2.1176
+ lwlc = 0
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ version = 4.5
+ moin = 5.5538
+ mjswgd = 0.95
+ mjswgs = 0.95
+ ijthsrev = 0.01
+ tempmod = 0
+ wvsat = -0.0037201203
+ nigc = 2.291
+ tcjswg = 0.00128
+ wvth0 = 5.188060000000002e-10
+ la0 = 3.4503642e-8
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = -0.0088528059
+ kt1 = -0.20733948
+ kt2 = -0.10130548
+ lk2 = 5.147862999999999e-9
+ waigc = 1.256895e-12
+ llc = 0
+ lln = 1
+ a0 = -0.1402156
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ lu0 = 3.380914000000001e-11
+ mjd = 0.335
+ mjs = 0.335
+ lua = 1.1003971e-16
+ lub = -1.3774164e-25
+ luc = -1.072064e-17
+ at = 113164.44
+ lud = 0
+ cf = 8.741900000000001e-11
+ lwc = 0
+ pvfbsdoff = 0
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.044448444
+ k3 = -2.5823
+ lwl = 0
+ lwn = 1
+ em = 20000000.0
+ aigbacc = 0.012071
+ njd = 1.02
+ njs = 1.02
+ ll = 0
+ noff = 2.2684
+ pa0 = -6.959911e-15
+ lw = 0
+ u0 = 0.0056368169
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ w0 = 0
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 1.1859675e-9
+ ua = -2.4996932e-9
+ ub = 3.4375966e-18
+ uc = 7.7964547e-11
+ ud = 0
+ pbs = 0.75
+ pk2 = -8.547569e-17
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 2.33e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ pu0 = 1.7354186999999972e-18
+ prt = 0
+ lketa = 2.7820203e-10
+ pua = -5.4706466e-24
+ pub = 7.864388699999999e-33
+ puc = 2.7207836e-25
+ pud = 0
+ wtvfbsdoff = 0
+ xpart = 1
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = -8.7447052e-10
+ ub1 = 1.4693195e-18
+ uc1 = -1.8902037e-10
+ ppdiblc2 = 3.8953385e-18
+ ntox = 2.958
+ tpb = 0.0016
+ pcit = -3.76965667e-17
+ pclm = 2.4870084
+ wa0 = 1.612455e-8
+ ute = -0.77766872
+ wat = -0.015568853
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 5.3174549e-9
+ aigbinv = 0.009974
+ wlc = 0
+ egidl = 0.001
+ wln = 1
+ wu0 = 1.8877321000000002e-10
+ xgl = -8.2e-9
+ xgw = 0
+ wua = 7.6741379e-17
+ wub = -1.2724134000000002e-25
+ wuc = 2.7069183e-18
+ wud = 0
+ wwc = 0
+ ltvfbsdoff = 0
+ wwl = 0
+ wwn = 1
+ phin = 0.15
+ fprout = 200
+ xrcrg1 = 12
+ xrcrg2 = 1
+ pkt1 = 1.2443873e-15
+ pkt2 = -4.056551e-17
+ wtvoff = -2.1192558e-10
+ pkvth0we = 0.0
+ rbdb = 50
+ pua1 = -1.3715808e-23
+ prwb = 0
+ pub1 = 1.7954113e-32
+ prwg = 0
+ puc1 = -3.4096566e-24
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ pute = 3.5590791e-15
+ )

.model pch_ff_39 pmos (
+ level = 54
+ fnoimod = 1
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ eigbinv = 1.1
+ k2we = 5e-5
+ ijthsfwd = 0.01
+ tvoff = 0.00092289205
+ dsub = 0.5
+ dtox = 3.91e-10
+ xjbvd = 1
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ xjbvs = 1
+ lk2we = 0.0
+ eta0 = 0.19463541
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ etab = -0.16706384
+ ijthsrev = 0.01
+ cigbacc = 0.245
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = -1.4247657000000001e-9
+ letab = 5.1546845e-9
+ tnoimod = 0
+ ppclm = 7.8094068e-15
+ dlcig = 2.5e-9
+ cigbinv = 0.006
+ bgidl = 1834800000.0
+ ppdiblc2 = 0
+ toxref = 3e-9
+ version = 4.5
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ tempmod = 0
+ ags = 1.2522222
+ cjd = 0.0012517799999999999
+ cit = 0.0091909913
+ cjs = 0.0012517799999999999
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 4.0349e-9
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ aigbacc = 0.012071
+ bigsd = 0.0003327
+ pkvth0we = 0.0
+ la0 = -1.4904033e-7
+ ltvoff = 2.8860613e-11
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0.008572508999999999
+ kt1 = -0.53950997
+ kt2 = -0.12590838
+ lk2 = 3.8165993e-9
+ wvoff = 1.4341134e-10
+ llc = 0
+ lln = 1
+ lu0 = 4.0451088999999997e-10
+ mjd = 0.335
+ mjs = 0.335
+ lua = 7.9060667e-17
+ lub = -1.2409918e-26
+ luc = 5.5424848e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = -2.574678e-15
+ nsd = 1e+20
+ pbd = 0.75
+ pat = -1.0212358e-9
+ wvsat = -0.0027183660000000003
+ pbs = 0.75
+ pk2 = 2.1304022e-16
+ aigbinv = 0.009974
+ wvth0 = -6.603598e-9
+ pu0 = -6.6237547e-17
+ vfbsdoff = 0.01
+ prt = 0
+ pua = -2.0419953e-23
+ pub = 1.0397510000000001e-32
+ puc = 1.2609666e-24
+ pud = 0
+ waigc = 6.0357037e-12
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 8.3453493e-9
+ ub1 = -1.1410668e-17
+ pvfbsdoff = 0
+ uc1 = 1.6197295e-9
+ keta = -0.31465021
+ lku0we = 1.8e-11
+ tpb = 0.0016
+ wa0 = -5.9482929e-8
+ epsrox = 3.9
+ ute = -1
+ wat = 0.022486376
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 1.7062889e-10
+ wlc = 0
+ wln = 1
+ wu0 = 1.3607208999999997e-9
+ xgl = -8.2e-9
+ xgw = 0
+ wua = 3.3448805e-16
+ wub = -1.7091596e-25
+ wuc = -1.434288e-17
+ wud = 0
+ lketa = 1.5671934e-8
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ paramchk = 1
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = -4.1881614e-10
+ xpart = 1
+ rdsmod = 0
+ kt1l = 0
+ igbmod = 1
+ egidl = 0.001
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ lint = 0
+ poxedge = 1
+ pbswgd = 0.8
+ pbswgs = 0.8
+ lkt1 = 1.3271281e-8
+ lkt2 = 2.350723e-9
+ lmax = 5.567e-8
+ lmin = 4.667e-8
+ ijthdfwd = 0.01
+ igcmod = 1
+ binunit = 2
+ lpe0 = 6.44e-8
+ lpeb = 0
+ minv = -0.33
+ lua1 = -3.7660644e-16
+ lub1 = 5.1040674e-25
+ luc1 = -7.3441373e-17
+ ndep = 1e+18
+ lwlc = 0
+ ijthdrev = 0.01
+ moin = 5.5538
+ nigc = 2.291
+ lpdiblc2 = 0
+ pvoff = 3.9992158e-17
+ cdscb = 0
+ cdscd = 0
+ pvsat = 1.14858808e-10
+ noff = 2.2684
+ wk2we = 0.0
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ pvth0 = 5.02207603e-16
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ permod = 1
+ drout = 0.56
+ paigc = -1.4334713e-18
+ voffl = 0
+ ntox = 2.958
+ pcit = 5.0064882e-17
+ pclm = 1.8533357
+ weta0 = -4.3683037e-9
+ wetab = 2.5894049e-9
+ lpclm = -6.4524768e-8
+ lkvth0we = 3e-12
+ phin = 0.15
+ voffcv = -0.125
+ wpemod = 1
+ pkt1 = -1.6683146e-15
+ pkt2 = -1.1786798e-16
+ cgidl = 1
+ acnqsmod = 0
+ njtsswg = 6.489
+ rbdb = 50
+ pua1 = 1.8341764e-23
+ prwb = 0
+ pub1 = -1.3009877e-32
+ prwg = 0
+ puc1 = 9.9681375e-24
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ pbswd = 0.9
+ rbpb = 50
+ rbpd = 50
+ pbsws = 0.9
+ rbps = 50
+ rbodymod = 0
+ rbsb = 50
+ pvag = 2.1
+ ckappad = 0.6
+ ckappas = 0.6
+ rdsw = 200
+ pdiblc1 = 0
+ pdiblc2 = 0.0014658889
+ pdiblcb = 0
+ tpbswg = 0.001
+ pdits = 0
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ bigbacc = 0.0054401
+ ptvoff = -2.2999757e-17
+ pk2we = 0.0
+ wpdiblc2 = 1.4741467e-10
+ rshg = 14.1
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ waigsd = 1.9716411e-12
+ kvth0we = -0.00022
+ diomod = 1
+ tnoia = 0
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ pditsd = 0
+ pditsl = 0
+ vtsswgd = 1.1
+ peta0 = 2.43224906e-17
+ vtsswgs = 1.1
+ cjswgd = 1.6832999999999998e-10
+ pku0we = 0.0
+ cjswgs = 1.6832999999999998e-10
+ petab = -2.558443e-17
+ wketa = 3.409679e-8
+ tpbsw = 0.0025
+ tnom = 25
+ cjswd = 4.743e-11
+ cjsws = 4.743e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ tvfbsdoff = 0.1
+ toxe = 2.6300000000000002e-9
+ toxm = 2.67e-9
+ wkvth0we = 0.0
+ mjswgd = 0.95
+ mjswgs = 0.95
+ wtvfbsdoff = 0
+ tcjswg = 0.00128
+ trnqsmod = 0
+ ltvfbsdoff = 0
+ wags = 2.5054667e-7
+ wcit = -1.09843482e-9
+ scref = 1e-6
+ voff = -0.1005239
+ pigcd = 2.572
+ acde = 0.5
+ aigsd = 0.0063632396
+ nfactor = 1
+ rgatemod = 0
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ tnjtsswg = 1
+ vsat = 107293.6
+ wint = 0
+ lvoff = -3.8177557e-9
+ vth0 = -0.17278243999999998
+ fprout = 200
+ wkt1 = 3.6711578e-8
+ wkt2 = 3.2153756e-9
+ wmax = 2.674e-7
+ xrcrg1 = 12
+ xrcrg2 = 1
+ aigc = 0.0068691843
+ wmin = 1.08e-7
+ lvsat = -0.00101193296
+ lvth0 = -8.0141177e-9
+ ptvfbsdoff = 0
+ delta = 0.018814
+ laigc = -1.683393e-11
+ wtvoff = 5.2119196e-10
+ wua1 = -3.864028e-16
+ wub1 = 3.2172349e-25
+ wuc1 = -2.0479093e-16
+ rnoia = 0
+ rnoib = 0
+ a0 = 3.0243356
+ a1 = 0
+ a2 = 1
+ nigbacc = 10
+ b0 = 0
+ b1 = 0
+ at = -187272.02
+ cf = 8.741900000000001e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.021495622
+ k3 = -2.5823
+ em = 20000000.0
+ bigc = 0.0012521
+ ll = 0
+ lw = 0
+ u0 = -0.0007545925899999995
+ w0 = 0
+ wwlc = 0
+ ua = -1.9655718e-9
+ ub = 1.2767046e-18
+ uc = -2.0243416e-10
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 2.33e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ pketa = -2.1465872e-15
+ ngate = 1.7e+20
+ ngcon = 1
+ capmod = 2
+ wpclm = -1.4226467e-7
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.2212350000000004e-11
+ cgdo = 2.8335740000000002e-11
+ wku0we = 1.5e-11
+ xtid = 3
+ xtis = 3
+ gbmin = 1e-12
+ nigbinv = 2.171
+ cgsl = 3.2212350000000004e-11
+ cgso = 2.8335740000000002e-11
+ cigc = 0.15259
+ jswgd = 3.69e-13
+ mobmod = 0
+ jswgs = 3.69e-13
+ )

.model pch_ff_40 pmos (
+ level = 54
+ fnoimod = 1
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ eigbinv = 1.1
+ laigsd = 6.1219753e-16
+ k2we = 5e-5
+ ijthsfwd = 0.01
+ tvoff = -0.00058332606
+ dsub = 0.5
+ dtox = 3.91e-10
+ xjbvd = 1
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ xjbvs = 1
+ lk2we = 0.0
+ eta0 = 0.11700471
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ etab = -0.15063456
+ ijthsrev = 0.01
+ cigbacc = 0.245
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = 2.3791388999999998e-9
+ letab = 4.3496496e-9
+ tnoimod = 0
+ ppclm = -3.5647768e-15
+ dlcig = 2.5e-9
+ cigbinv = 0.006
+ bgidl = 1834800000.0
+ ppdiblc2 = 0
+ toxref = 3e-9
+ version = 4.5
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ tempmod = 0
+ ags = 1.2522222
+ cjd = 0.0012517799999999999
+ cit = -0.0151232499
+ cjs = 0.0012517799999999999
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 4.0349e-9
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ aigbacc = 0.012071
+ bigsd = 0.0003327
+ pkvth0we = 0.0
+ la0 = -3.4726683e-8
+ ltvoff = 1.026653e-10
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0.0011579456999999999
+ kt1 = -0.60072817
+ kt2 = -0.12562663
+ lk2 = 5.8841473e-9
+ wvoff = 3.3909703e-9
+ llc = 0
+ lln = 1
+ lu0 = 5.1441728e-10
+ mjd = 0.335
+ mjs = 0.335
+ lua = 9.0470184e-17
+ lub = 2.1169426e-26
+ luc = 2.7216576e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 1.4761752e-15
+ nsd = 1e+20
+ pbd = 0.75
+ pat = -2.09104015e-10
+ wvsat = -0.009856557
+ pbs = 0.75
+ pk2 = -2.7720832e-16
+ aigbinv = 0.009974
+ wvth0 = 1.185091359e-8
+ pu0 = -6.1923224e-17
+ vfbsdoff = 0.01
+ prt = 0
+ pua = -4.2432063e-24
+ pub = -9.3890685e-33
+ puc = -1.7176927e-24
+ pud = 0
+ waigc = -4.0606639e-11
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 2.1566906e-9
+ ub1 = -1.4553545999999999e-18
+ pvfbsdoff = 0
+ uc1 = -1.7258848e-10
+ keta = 0.15497942
+ lku0we = 1.8e-11
+ tpb = 0.0016
+ wa0 = -1.421534e-7
+ epsrox = 3.9
+ ute = -1
+ wat = 0.0059122670000000006
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 1.0175701e-8
+ wlc = 0
+ wln = 1
+ wu0 = 1.2726735e-9
+ xgl = -8.2e-9
+ xgw = 0
+ wua = 4.3503521e-18
+ wub = 2.3289192e-25
+ wuc = 4.6446086e-17
+ wud = 0
+ lketa = -7.3399177e-9
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ paramchk = 1
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 7.725810299999999e-10
+ xpart = 1
+ rdsmod = 0
+ kt1l = 0
+ igbmod = 1
+ egidl = 0.001
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ lint = 0
+ poxedge = 1
+ pbswgd = 0.8
+ pbswgs = 0.8
+ lkt1 = 1.62709929e-8
+ lkt2 = 2.3369169e-9
+ lmax = 4.667e-8
+ lmin = 3.6e-8
+ ijthdfwd = 0.01
+ igcmod = 1
+ binunit = 2
+ lpe0 = 6.44e-8
+ lpeb = 0
+ minv = -0.33
+ lua1 = -7.3362164e-17
+ lub1 = 2.2595779999999982e-26
+ luc1 = 1.4382206e-17
+ ndep = 1e+18
+ lwlc = 0
+ ijthdrev = 0.01
+ moin = 5.5538
+ nigc = 2.291
+ paigsd = -6.9790518e-23
+ lpdiblc2 = 0
+ pvoff = -1.19138231e-16
+ cdscb = 0
+ cdscd = 0
+ pvsat = 4.6462985999999997e-10
+ noff = 2.2684
+ wk2we = 0.0
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ pvth0 = -4.0206497e-16
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ permod = 1
+ drout = 0.56
+ paigc = 8.520035e-19
+ voffl = 0
+ ntox = 2.958
+ pcit = -1.3690619999999969e-18
+ pclm = 0.41497396
+ weta0 = -9.956769999999999e-10
+ wetab = 1.1541057e-8
+ lpclm = 5.9549575e-9
+ lkvth0we = 3e-12
+ phin = 0.15
+ voffcv = -0.125
+ wpemod = 1
+ pkt1 = -3.3136614e-15
+ pkt2 = -7.0509572e-16
+ cgidl = 1
+ acnqsmod = 0
+ njtsswg = 6.489
+ rbdb = 50
+ pua1 = 3.2441676e-23
+ prwb = 0
+ pub1 = -4.1973804e-32
+ prwg = 0
+ puc1 = -1.3788915e-24
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ pbswd = 0.9
+ rbpb = 50
+ rbpd = 50
+ pbsws = 0.9
+ rbps = 50
+ rbodymod = 0
+ rbsb = 50
+ pvag = 2.1
+ ckappad = 0.6
+ ckappas = 0.6
+ rdsw = 200
+ pdiblc1 = 0
+ pdiblc2 = 0.0014658889
+ pdiblcb = 0
+ tpbswg = 0.001
+ pdits = 0
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ bigbacc = 0.0054401
+ ptvoff = -3.9364956e-17
+ pk2we = 0.0
+ wpdiblc2 = 1.4741467e-10
+ rshg = 14.1
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ waigsd = 1.9730654e-12
+ kvth0we = -0.00022
+ diomod = 1
+ tnoia = 0
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ pditsd = 0
+ pditsl = 0
+ vtsswgd = 1.1
+ peta0 = -1.4093622e-16
+ vtsswgs = 1.1
+ cjswgd = 1.6832999999999998e-10
+ pku0we = 0.0
+ cjswgs = 1.6832999999999998e-10
+ petab = -4.6421536e-16
+ wketa = -5.7187654e-8
+ tpbsw = 0.0025
+ tnom = 25
+ cjswd = 4.743e-11
+ cjsws = 4.743e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ tvfbsdoff = 0.1
+ toxe = 2.6300000000000002e-9
+ toxm = 2.67e-9
+ wkvth0we = 0.0
+ mjswgd = 0.95
+ mjswgs = 0.95
+ wtvfbsdoff = 0
+ tcjswg = 0.00128
+ trnqsmod = 0
+ ltvfbsdoff = 0
+ wags = 2.5054667e-7
+ wcit = -4.877341000000002e-11
+ scref = 1e-6
+ voff = -0.12231559
+ pigcd = 2.572
+ acde = 0.5
+ aigsd = 0.0063632271
+ nfactor = 1
+ rgatemod = 0
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ tnjtsswg = 1
+ vsat = 133672.58000000002
+ wint = 0
+ lvoff = -2.7499629e-9
+ vth0 = -0.42676907
+ fprout = 200
+ wkt1 = 7.0290182e-8
+ wkt2 = 1.5199615e-8
+ wmax = 2.674e-7
+ xrcrg1 = 12
+ xrcrg2 = 1
+ aigc = 0.0069354083
+ wmin = 1.08e-7
+ lvsat = -0.0023044963999999998
+ lvth0 = 4.431213099999999e-9
+ ptvfbsdoff = 0
+ delta = 0.018814
+ laigc = -2.0078906e-11
+ wtvoff = 8.5517561e-10
+ wua1 = -6.7415611e-16
+ wub1 = 9.128243e-25
+ wuc1 = 2.6781086e-17
+ rnoia = 0
+ rnoib = 0
+ a0 = 0.69140412
+ a1 = 0
+ a2 = 1
+ nigbacc = 10
+ b0 = 0
+ b1 = 0
+ at = -35954.44
+ cf = 8.741900000000001e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.06369048
+ k3 = -2.5823
+ em = 20000000.0
+ bigc = 0.0012521
+ ll = 0
+ lw = 0
+ u0 = -0.0029975803
+ w0 = 0
+ wwlc = 0
+ ua = -2.1984191e-9
+ ub = 5.914109e-19
+ uc = -1.4486626e-10
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 2.33e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ pketa = 2.3263506e-15
+ ngate = 1.7e+20
+ ngcon = 1
+ capmod = 2
+ wpclm = 8.9861524e-8
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.2212350000000004e-11
+ cgdo = 2.8335740000000002e-11
+ wku0we = 1.5e-11
+ xtid = 3
+ xtis = 3
+ gbmin = 1e-12
+ nigbinv = 2.171
+ cgsl = 3.2212350000000004e-11
+ cgso = 2.8335740000000002e-11
+ cigc = 0.15259
+ jswgd = 3.69e-13
+ mobmod = 0
+ jswgs = 3.69e-13
+ )

.model pch_fs_1 pmos (
+ level = 54
+ ppclm = 0
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ bigbacc = 0.0054401
+ wpdiblc2 = 0
+ tnom = 25
+ kvth0we = -0.00022
+ tvfbsdoff = 0.1
+ dmcgt = 0
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ tcjsw = 9.34e-5
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ toxref = 3e-9
+ bigsd = 0.0003327
+ wkvth0we = 0.0
+ wvoff = 0
+ trnqsmod = 0
+ voff = -0.11110337
+ acde = 0.5
+ wvsat = 0
+ wvfbsdoff = 0
+ wvth0 = -2.1600000000000004e-9
+ lvfbsdoff = 0
+ vsat = 120000
+ wint = 0
+ vth0 = -0.40913527
+ ltvoff = 0
+ wmax = 0.00090001
+ aigc = 0.0068307507
+ wmin = 9.0026e-6
+ a0 = 2.531
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 72000
+ cf = 8.17e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.00077592763
+ k3 = -2.5823
+ em = 20000000.0
+ lketa = 0
+ ll = 0
+ lw = 0
+ u0 = 0.009875
+ w0 = 0
+ rgatemod = 0
+ ua = 1.297e-10
+ ub = 1.182572e-18
+ uc = 2.014e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xpart = 1
+ xw = 3.4e-9
+ nfactor = 1
+ tnjtsswg = 1
+ lku0we = 1.8e-11
+ bigc = 0.0012521
+ egidl = 0.001
+ wwlc = 0
+ epsrox = 3.9
+ cdsc = 0
+ rdsmod = 0
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ igbmod = 1
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigc = 0.15259
+ nigbacc = 10
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ pbswgd = 0.8
+ pbswgs = 0.8
+ igcmod = 1
+ nigbinv = 2.171
+ pvoff = 2e-17
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ cdscb = 0
+ cdscd = 0
+ pvsat = 0
+ wk2we = 0.0
+ pvth0 = -1.2e-16
+ drout = 0.56
+ k2we = 5e-5
+ dsub = 0.5
+ dtox = 3.91e-10
+ voffl = 0
+ fnoimod = 1
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ eigbinv = 1.1
+ weta0 = -2.2400000000000003e-10
+ permod = 1
+ lpclm = 0
+ eta0 = 0.1672
+ etab = -0.23
+ ijthsfwd = 0.01
+ cgidl = 1
+ voffcv = -0.125
+ wpemod = 1
+ ijthsrev = 0.01
+ pbswd = 0.9
+ pbsws = 0.9
+ cigbacc = 0.245
+ tnoimod = 0
+ pdits = 0
+ cigsd = 0.013281
+ cigbinv = 0.006
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ ppdiblc2 = 0
+ tpbswg = 0.001
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ version = 4.5
+ tempmod = 0
+ tnoia = 0
+ peta0 = -1.6e-17
+ ptvoff = 0
+ aigbacc = 0.012071
+ tpbsw = 0.0025
+ pkvth0we = 0.0
+ pvfbsdoff = 0
+ keta = -0.042350111
+ cjswd = 5.3856e-11
+ cjsws = 5.3856e-11
+ diomod = 1
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ pditsd = 0
+ pditsl = 0
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ cjswgd = 1.9113600000000002e-10
+ pku0we = 0.0
+ cjswgs = 1.9113600000000002e-10
+ lcit = 1.6e-11
+ aigbinv = 0.009974
+ vfbsdoff = 0.01
+ wtvfbsdoff = 0
+ kt1l = 0
+ lint = 6.5375218e-9
+ ltvfbsdoff = 0
+ mjswgd = 0.95
+ mjswgs = 0.95
+ lkt1 = -4.8e-10
+ paramchk = 1
+ lmax = 2.001e-5
+ lmin = 8.9991e-6
+ tcjswg = 0.00128
+ scref = 1e-6
+ lpe0 = 6.44e-8
+ lpeb = 0
+ pigcd = 2.572
+ aigsd = 0.0063636
+ minv = -0.33
+ lvoff = 0
+ poxedge = 1
+ ndep = 1e+18
+ lwlc = 0
+ ijthdfwd = 0.01
+ lvsat = 8.000000000000001e-6
+ moin = 5.5538
+ lvth0 = -2.4e-10
+ binunit = 2
+ ptvfbsdoff = 0
+ nigc = 2.291
+ delta = 0.018814
+ rnoia = 0
+ rnoib = 0
+ fprout = 200
+ noff = 2.2684
+ ags = 0.8379228
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ ijthdrev = 0.01
+ ngate = 1.7e+20
+ cjd = 0.001421376
+ cit = 5e-6
+ cjs = 0.001421376
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 1.0572421799999999e-8
+ ngcon = 1
+ k3b = 2.1176
+ wpclm = 0
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ lpdiblc2 = 0
+ ntox = 1.0
+ wtvoff = 0
+ pcit = -8.000000000000001e-19
+ pclm = 1.484
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ la0 = 0
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0.00064
+ kt1 = -0.17107633
+ lk2 = 3.2000000000000003e-10
+ kt2 = -0.04747
+ jtsswgd = 1.75e-7
+ phin = 0.15
+ llc = 0
+ jtsswgs = 1.75e-7
+ lln = 1
+ lu0 = -8e-13
+ mjd = 0.335
+ mjs = 0.335
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 0
+ capmod = 2
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ pk2 = 0
+ pkt1 = -4e-17
+ pu0 = 0
+ prt = 0
+ wku0we = 1.5e-11
+ pud = 0
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 1.1969344e-9
+ ub1 = -1.3666143e-18
+ uc1 = 6.873e-11
+ mobmod = 0
+ tpb = 0.0016
+ wa0 = 0
+ lkvth0we = 3e-12
+ ute = -1
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 0
+ wlc = 0
+ wln = 1
+ rbdb = 50
+ prwb = 0
+ wu0 = 0
+ prwg = 0
+ xgl = -8.2e-9
+ xgw = 0
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ rdsw = 200
+ tvoff = 0.0026155642
+ acnqsmod = 0
+ njtsswg = 6.489
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ xtsswgd = 0.32
+ rbodymod = 0
+ xtsswgs = 0.32
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.0026729629
+ ku0we = -0.0007
+ pdiblcb = 0
+ beta0 = 13.32
+ rshg = 14.1
+ leta0 = -4.8e-10
+ )

.model pch_fs_2 pmos (
+ level = 54
+ aigbinv = 0.009974
+ eta0 = 0.1672
+ tnoia = 0
+ etab = -0.23
+ ijthdfwd = 0.01
+ peta0 = -1.6e-17
+ toxref = 3e-9
+ pvfbsdoff = 0
+ tpbsw = 0.0025
+ cjswd = 5.3856e-11
+ cjsws = 5.3856e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ ijthdrev = 0.01
+ lpdiblc2 = 7.1311563e-9
+ poxedge = 1
+ ltvoff = -4.7585658e-10
+ binunit = 2
+ scref = 1e-6
+ pigcd = 2.572
+ aigsd = 0.0063636
+ lku0we = 1.8e-11
+ epsrox = 3.9
+ lkvth0we = 3e-12
+ lvoff = -8.0044387e-9
+ lvsat = 8.000000000000001e-6
+ rdsmod = 0
+ lvth0 = -5.3667661e-9
+ ags = 0.80385259
+ igbmod = 1
+ delta = 0.018814
+ laigc = -4.8397409e-11
+ cjd = 0.001421376
+ cit = 5e-6
+ cjs = 0.001421376
+ clc = 1e-7
+ cle = 0.6
+ acnqsmod = 0
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 1.0572421799999999e-8
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ k3b = 2.1176
+ rnoia = 0
+ rnoib = 0
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ keta = -0.040853613
+ pbswgd = 0.8
+ pbswgs = 0.8
+ rbodymod = 0
+ a0 = 2.5747309
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 72000
+ lags = 3.062912e-7
+ ngate = 1.7e+20
+ cf = 8.17e-11
+ igcmod = 1
+ la0 = -3.9314047e-7
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.0012551498
+ k3 = -2.5823
+ em = 20000000.0
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0.00064
+ ll = 0
+ lw = 0
+ kt1 = -0.16652617
+ kt2 = -0.046491549
+ lk2 = 4.6282075e-9
+ u0 = 0.0098748901
+ ngcon = 1
+ w0 = 0
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ ua = 1.4083134e-10
+ ub = 1.1675774e-18
+ uc = 1.8373185e-11
+ ud = 0
+ llc = 0
+ wpclm = 0
+ lln = 1
+ lcit = 1.6e-11
+ wl = 0
+ wr = 1
+ lu0 = 1.8779011999999998e-13
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 3.4e-9
+ mjd = 0.335
+ mjs = 0.335
+ lua = -1.0007073e-16
+ lub = 1.3480174e-25
+ luc = 1.5883665e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ kt1l = 0
+ njs = 1.02
+ pa0 = 0
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ pk2 = 0
+ gbmin = 1e-12
+ pu0 = 0
+ jswgd = 3.69e-13
+ prt = 0
+ jswgs = 3.69e-13
+ pud = 0
+ lint = 6.5375218e-9
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 1.1817684e-9
+ ub1 = -1.3634053e-18
+ uc1 = 6.7786161e-11
+ tpb = 0.0016
+ lkt1 = -4.1386013000000005e-8
+ lkt2 = -8.7962711e-9
+ wa0 = 0
+ lmax = 8.9991e-6
+ ute = -1
+ lmin = 8.9908e-7
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 0
+ wlc = 0
+ wln = 1
+ wu0 = 0
+ xgl = -8.2e-9
+ xgw = 0
+ njtsswg = 6.489
+ lpe0 = 6.44e-8
+ wud = 0
+ wpdiblc2 = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ lpeb = 0
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ minv = -0.33
+ lua1 = 1.3634229e-16
+ lub1 = -2.8849398e-26
+ luc1 = 8.4851172e-18
+ permod = 1
+ ckappad = 0.6
+ ckappas = 0.6
+ ndep = 1e+18
+ pdiblc1 = 0
+ pdiblc2 = 0.0018797309
+ pdiblcb = 0
+ lwlc = 0
+ moin = 5.5538
+ nigc = 2.291
+ tvoff = 0.002668496
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ wkvth0we = 0.0
+ voffcv = -0.125
+ wpemod = 1
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ bigbacc = 0.0054401
+ trnqsmod = 0
+ ku0we = -0.0007
+ beta0 = 13.32
+ kvth0we = -0.00022
+ ntox = 1.0
+ pcit = -8.000000000000001e-19
+ pclm = 1.484
+ leta0 = -4.8e-10
+ lintnoi = -5e-9
+ ppclm = 0
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ phin = 0.15
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ pkt1 = -4e-17
+ rgatemod = 0
+ tpbswg = 0.001
+ tnjtsswg = 1
+ tvfbsdoff = 0.1
+ dmcgt = 0
+ rbdb = 50
+ tcjsw = 9.34e-5
+ prwb = 0
+ prwg = 0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ ptvoff = 0
+ wtvfbsdoff = 0
+ rdsw = 200
+ bigsd = 0.0003327
+ diomod = 1
+ ltvfbsdoff = 0
+ pditsd = 0
+ pditsl = 0
+ nfactor = 1
+ wvoff = 0
+ cjswgd = 1.9113600000000002e-10
+ pku0we = 0.0
+ cjswgs = 1.9113600000000002e-10
+ wvfbsdoff = 0
+ wvsat = 0
+ lvfbsdoff = 0
+ wvth0 = -2.1600000000000004e-9
+ rshg = 14.1
+ mjswgd = 0.95
+ mjswgs = 0.95
+ tcjswg = 0.00128
+ lketa = -1.3453518e-8
+ ptvfbsdoff = 0
+ nigbacc = 10
+ xpart = 1
+ tnom = 25
+ egidl = 0.001
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ ijthsfwd = 0.01
+ nigbinv = 2.171
+ fprout = 200
+ xrcrg1 = 12
+ xrcrg2 = 1
+ ijthsrev = 0.01
+ fnoimod = 1
+ voff = -0.110213
+ wtvoff = 0
+ acde = 0.5
+ eigbinv = 1.1
+ pvoff = 2e-17
+ vsat = 120000
+ wint = 0
+ vth0 = -0.408565
+ cdscb = 0
+ cdscd = 0
+ wmax = 0.00090001
+ pvsat = 0
+ aigc = 0.0068361342
+ wmin = 9.0026e-6
+ wk2we = 0.0
+ capmod = 2
+ pvth0 = -1.2e-16
+ drout = 0.56
+ wku0we = 1.5e-11
+ ppdiblc2 = 0
+ mobmod = 0
+ voffl = 0
+ bigc = 0.0012521
+ weta0 = -2.2400000000000003e-10
+ cigbacc = 0.245
+ wwlc = 0
+ lpclm = 0
+ cdsc = 0
+ tnoimod = 0
+ cgbo = 0
+ cgidl = 1
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigc = 0.15259
+ pkvth0we = 0.0
+ cigbinv = 0.006
+ pbswd = 0.9
+ pbsws = 0.9
+ vfbsdoff = 0.01
+ version = 4.5
+ tempmod = 0
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ pdits = 0
+ cigsd = 0.013281
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ dvt0w = 0
+ paramchk = 1
+ dvt1w = 0
+ dvt2w = 0
+ aigbacc = 0.012071
+ k2we = 5e-5
+ dsub = 0.5
+ dtox = 3.91e-10
+ pk2we = 0.0
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ )

.model pch_fs_3 pmos (
+ level = 54
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ nigbacc = 10
+ ijthsrev = 0.01
+ wvoff = 0
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ wvsat = 0
+ ntox = 1.0
+ wvth0 = -2.1600000000000004e-9
+ pcit = -8.000000000000001e-19
+ pclm = 1.484
+ ltvoff = -2.3123852e-10
+ nigbinv = 2.171
+ phin = 0.15
+ lketa = -1.5940244e-8
+ pkt1 = -4e-17
+ ppdiblc2 = 0
+ xpart = 1
+ lku0we = 1.8e-11
+ epsrox = 3.9
+ egidl = 0.001
+ rbdb = 50
+ fnoimod = 1
+ prwb = 0
+ prwg = 0
+ rdsmod = 0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ eigbinv = 1.1
+ igbmod = 1
+ rdsw = 200
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ pbswgd = 0.8
+ pbswgs = 0.8
+ pkvth0we = 0.0
+ igcmod = 1
+ vfbsdoff = 0.01
+ rshg = 14.1
+ cigbacc = 0.245
+ pvoff = 2e-17
+ cdscb = 0
+ cdscd = 0
+ pvsat = 0
+ tnoimod = 0
+ wk2we = 0.0
+ pvth0 = -1.2e-16
+ paramchk = 1
+ drout = 0.56
+ cigbinv = 0.006
+ voffl = 0
+ permod = 1
+ tnom = 25
+ weta0 = -2.2400000000000003e-10
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ a0 = 2.8917556
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ lpclm = 0
+ at = 72000
+ cf = 8.17e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = 0.0040664684
+ k3 = -2.5823
+ em = 20000000.0
+ ijthdfwd = 0.01
+ version = 4.5
+ ll = 0
+ lw = 0
+ u0 = 0.010106756
+ w0 = 0
+ ua = 1.1413788e-10
+ ub = 1.1978347e-18
+ uc = 4.3035111e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 3.4e-9
+ tempmod = 0
+ cgidl = 1
+ voffcv = -0.125
+ wpemod = 1
+ aigbacc = 0.012071
+ ijthdrev = 0.01
+ pbswd = 0.9
+ pbsws = 0.9
+ voff = -0.10886793
+ lpdiblc2 = 1.7469722e-9
+ acde = 0.5
+ vsat = 120000
+ aigbinv = 0.009974
+ wint = 0
+ vth0 = -0.41118963000000003
+ pdits = 0
+ cigsd = 0.013281
+ wmax = 0.00090001
+ aigc = 0.00683106
+ wmin = 9.0026e-6
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ wtvfbsdoff = 0
+ tpbswg = 0.001
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ ltvfbsdoff = 0
+ lkvth0we = 3e-12
+ bigc = 0.0012521
+ wwlc = 0
+ tnoia = 0
+ ptvoff = 0
+ poxedge = 1
+ cdsc = 0
+ peta0 = -1.6e-17
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ acnqsmod = 0
+ pvfbsdoff = 0
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigc = 0.15259
+ binunit = 2
+ diomod = 1
+ tpbsw = 0.0025
+ cjswd = 5.3856e-11
+ cjsws = 5.3856e-11
+ mjswd = 0.01
+ pditsd = 0
+ mjsws = 0.01
+ pditsl = 0
+ rbodymod = 0
+ agidl = 3.2166e-9
+ cjswgd = 1.9113600000000002e-10
+ pku0we = 0.0
+ cjswgs = 1.9113600000000002e-10
+ ptvfbsdoff = 0
+ dmcg = 3.1e-8
+ mjswgd = 0.95
+ dmci = 3.1e-8
+ dmdg = 0
+ mjswgs = 0.95
+ tcjswg = 0.00128
+ k2we = 5e-5
+ jtsswgd = 1.75e-7
+ scref = 1e-6
+ jtsswgs = 1.75e-7
+ wpdiblc2 = 0
+ dsub = 0.5
+ pigcd = 2.572
+ dtox = 3.91e-10
+ aigsd = 0.0063635603
+ ags = 0.82774541
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ lvoff = -9.201547e-9
+ cjd = 0.001421376
+ cit = -8.7888889e-5
+ cjs = 0.001421376
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 1.0572421799999999e-8
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ eta0 = 0.1672
+ etab = -0.23
+ lvsat = 8.000000000000001e-6
+ lvth0 = -3.0308401e-9
+ delta = 0.018814
+ laigc = -4.3881382e-11
+ la0 = -6.7529244e-7
+ fprout = 200
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0.00064
+ kt1 = -0.19559142
+ kt2 = -0.048919444
+ lk2 = -1.0803271999999996e-10
+ llc = 0
+ lln = 1
+ lu0 = -2.0617244e-10
+ rnoia = 0
+ rnoib = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ mjd = 0.335
+ mjs = 0.335
+ lua = -7.6313554e-17
+ lub = 1.0787275e-25
+ luc = -6.0654489e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ wkvth0we = 0.0
+ njs = 1.02
+ pa0 = 0
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ pk2 = 0
+ njtsswg = 6.489
+ pu0 = 0
+ prt = 0
+ pud = 0
+ ngate = 1.7e+20
+ trnqsmod = 0
+ wtvoff = 0
+ ngcon = 1
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 1.2804108e-9
+ ub1 = -1.1625424e-18
+ uc1 = 4.6637333e-11
+ wpclm = 0
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ tpb = 0.0016
+ wa0 = 0
+ ute = -1
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 0
+ ckappad = 0.6
+ ckappas = 0.6
+ gbmin = 1e-12
+ wlc = 0
+ wln = 1
+ wu0 = 0
+ xgl = -8.2e-9
+ xgw = 0
+ pdiblc1 = 0
+ pdiblc2 = 0.0079293759
+ wud = 0
+ jswgd = 3.69e-13
+ wwc = 0
+ jswgs = 3.69e-13
+ wwl = 0
+ wwn = 1
+ pdiblcb = 0
+ capmod = 2
+ wku0we = 1.5e-11
+ rgatemod = 0
+ mobmod = 0
+ tnjtsswg = 1
+ bigbacc = 0.0054401
+ kvth0we = -0.00022
+ lintnoi = -5e-9
+ tvoff = 0.0023936443
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ laigsd = 3.5374533e-14
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ keta = -0.03805954
+ lags = 2.8502658e-7
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 9.8671111e-11
+ ku0we = -0.0007
+ beta0 = 13.32
+ kt1l = 0
+ leta0 = -4.8e-10
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ ppclm = 0
+ lint = 6.5375218e-9
+ lkt1 = -1.5517938999999997e-8
+ lkt2 = -6.6354444e-9
+ dlcig = 2.5e-9
+ lmax = 8.9908e-7
+ bgidl = 1834800000.0
+ lmin = 4.4908e-7
+ lpe0 = 6.44e-8
+ lpeb = 0
+ tvfbsdoff = 0.1
+ minv = -0.33
+ lua1 = 4.8550568e-17
+ nfactor = 1
+ lub1 = -2.0761736e-25
+ luc1 = 2.7307573e-17
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ ndep = 1e+18
+ lwlc = 0
+ ijthsfwd = 0.01
+ moin = 5.5538
+ nigc = 2.291
+ toxref = 3e-9
+ bigsd = 0.0003327
+ )

.model pch_fs_4 pmos (
+ level = 54
+ aigc = 0.0067884199
+ wmin = 9.0026e-6
+ cjd = 0.001421376
+ cit = -0.00054497817
+ cjs = 0.001421376
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 1.38228675e-8
+ scref = 1e-6
+ k3b = 2.1176
+ rgatemod = 0
+ lku0we = 1.8e-11
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ pigcd = 2.572
+ tnjtsswg = 1
+ epsrox = 3.9
+ aigsd = 0.0063636407
+ njtsswg = 6.489
+ lvoff = -3.8830249e-9
+ bigc = 0.0012521
+ la0 = -4.3379389e-8
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0.00064
+ rdsmod = 0
+ kt1 = -0.2000222
+ kt2 = -0.054670852
+ lk2 = 1.6830221e-9
+ wwlc = 0
+ llc = -1.18e-13
+ xtsswgd = 0.32
+ lln = 0.7
+ xtsswgs = 0.32
+ lu0 = -4.840545000000001e-10
+ igbmod = 1
+ mjd = 0.335
+ mjs = 0.335
+ lua = -1.5477844e-16
+ lub = 5.0676856e-26
+ luc = -5.2541764e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ lvsat = 8.000000000000001e-6
+ njd = 1.02
+ njs = 1.02
+ pa0 = 0
+ lvth0 = 4.1004654e-9
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ ckappad = 0.6
+ pk2 = 0
+ ckappas = 0.6
+ cdsc = 0
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ pu0 = 0
+ pdiblc1 = 0
+ pdiblc2 = 0.013802718
+ delta = 0.018814
+ cgbo = 0
+ prt = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ pud = 0
+ pdiblcb = 0
+ xtid = 3
+ xtis = 3
+ laigc = -2.5119727e-11
+ pbswgd = 0.8
+ pbswgs = 0.8
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ rsh = 15.2
+ tcj = 0.000832
+ cigc = 0.15259
+ ua1 = 1.2553592e-9
+ ub1 = -1.2671808e-18
+ uc1 = 1.0455371e-10
+ rnoia = 0
+ rnoib = 0
+ tpb = 0.0016
+ wa0 = 0
+ igcmod = 1
+ ute = -1
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 0
+ wlc = 0
+ wln = 1
+ wu0 = 0
+ xgl = -8.2e-9
+ xgw = 0
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ ngate = 1.7e+20
+ ngcon = 1
+ wpclm = 0
+ bigbacc = 0.0054401
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ kvth0we = -0.00022
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ k2we = 5e-5
+ vtsswgs = 1.1
+ dsub = 0.5
+ dtox = 3.91e-10
+ permod = 1
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ eta0 = 0.1672
+ ijthsfwd = 0.01
+ etab = -0.23
+ tvoff = 0.002134918
+ voffcv = -0.125
+ wpemod = 1
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ ijthsrev = 0.01
+ wtvfbsdoff = 0
+ ku0we = -0.0007
+ beta0 = 13.32
+ nfactor = 1
+ leta0 = -4.8e-10
+ ltvfbsdoff = 0
+ ppclm = 0
+ a0 = 1.4555895
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 72000
+ cf = 8.17e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -4.1106394e-6
+ k3 = -2.5823
+ em = 20000000.0
+ ll = -1.18e-13
+ dlcig = 2.5e-9
+ lw = 0
+ u0 = 0.010738306
+ w0 = 0
+ tpbswg = 0.001
+ ua = 2.9246716e-10
+ ub = 1.3278253e-18
+ uc = 4.119131e-11
+ ud = 0
+ bgidl = 1834800000.0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 3.4e-9
+ ppdiblc2 = 0
+ tvfbsdoff = 0.1
+ nigbacc = 10
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ ptvoff = 0
+ ptvfbsdoff = 0
+ diomod = 1
+ nigbinv = 2.171
+ pkvth0we = 0.0
+ bigsd = 0.0003327
+ keta = -0.029364427
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.9113600000000002e-10
+ pku0we = 0.0
+ cjswgs = 1.9113600000000002e-10
+ wvoff = 0
+ lags = 5.4107004e-7
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 2.9979039e-10
+ vfbsdoff = 0.01
+ wvsat = 0
+ kt1l = 0
+ wvth0 = -2.1600000000000004e-9
+ mjswgd = 0.95
+ mjswgs = 0.95
+ fnoimod = 1
+ eigbinv = 1.1
+ tcjswg = 0.00128
+ lint = 9.7879675e-9
+ lkt1 = -1.3568393e-8
+ lkt2 = -4.1048253e-9
+ paramchk = 1
+ lmax = 4.4908e-7
+ lmin = 2.1577e-7
+ lketa = -1.9766093e-8
+ lpe0 = 6.44e-8
+ xpart = 1
+ lpeb = 0
+ minv = -0.33
+ lua1 = 5.9573279e-17
+ lub1 = -1.6157647e-25
+ egidl = 0.001
+ luc1 = 1.8243668e-18
+ ndep = 1e+18
+ lwlc = 0
+ ijthdfwd = 0.01
+ moin = 5.5538
+ cigbacc = 0.245
+ fprout = 200
+ nigc = 2.291
+ xrcrg1 = 12
+ xrcrg2 = 1
+ tnoimod = 0
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ ijthdrev = 0.01
+ cigbinv = 0.006
+ wtvoff = 0
+ lpdiblc2 = -8.3729822e-10
+ ntox = 1.0
+ pcit = -8.000000000000001e-19
+ pclm = 1.484
+ pvoff = 2e-17
+ capmod = 2
+ version = 4.5
+ cdscb = 0
+ cdscd = 0
+ pvsat = 0
+ phin = 0.15
+ wku0we = 1.5e-11
+ tempmod = 0
+ wk2we = 0.0
+ pvth0 = -1.2e-16
+ drout = 0.56
+ mobmod = 0
+ pkt1 = -4e-17
+ voffl = 0
+ aigbacc = 0.012071
+ lkvth0we = 3e-12
+ weta0 = -2.2400000000000003e-10
+ rbdb = 50
+ prwb = 0
+ prwg = 0
+ lpclm = 0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ rdsw = 200
+ aigbinv = 0.009974
+ cgidl = 1
+ acnqsmod = 0
+ rbodymod = 0
+ pbswd = 0.9
+ pbsws = 0.9
+ rshg = 14.1
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ pdits = 0
+ poxedge = 1
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ binunit = 2
+ wpdiblc2 = 0
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ tnom = 25
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ tnoia = 0
+ toxref = 3e-9
+ peta0 = -1.6e-17
+ pvfbsdoff = 0
+ tpbsw = 0.0025
+ wkvth0we = 0.0
+ cjswd = 5.3856e-11
+ cjsws = 5.3856e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ trnqsmod = 0
+ voff = -0.12095548
+ acde = 0.5
+ ltvoff = -1.1739897e-10
+ vsat = 120000
+ wint = 0
+ vth0 = -0.42739715
+ wmax = 0.00090001
+ ags = 0.24582847
+ )

.model pch_fs_5 pmos (
+ level = 54
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ pbswgd = 0.8
+ pbswgs = 0.8
+ acnqsmod = 0
+ version = 4.5
+ tempmod = 0
+ igcmod = 1
+ keta = -0.12863898
+ rbodymod = 0
+ lags = 3.2185083e-8
+ aigbacc = 0.012071
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 9.1945573e-11
+ kt1l = 0
+ pvoff = 2e-17
+ cdscb = 0
+ cdscd = 0
+ lint = 9.7879675e-9
+ pvsat = 0.0
+ wk2we = 0.0
+ pvth0 = -1.2e-16
+ aigbinv = 0.009974
+ lkt1 = -5.2209966e-9
+ lkt2 = -5.2805906e-10
+ drout = 0.56
+ lmax = 2.1577e-7
+ lmin = 9e-8
+ wpdiblc2 = 0
+ lpe0 = 6.44e-8
+ permod = 1
+ lpeb = 0
+ voffl = 0
+ minv = -0.33
+ lua1 = -1.5051887e-16
+ lub1 = 1.742578e-25
+ luc1 = 7.2216103e-18
+ weta0 = -2.2400000000000003e-10
+ ndep = 1e+18
+ lpclm = -1.4239795e-8
+ wtvfbsdoff = 0
+ lwlc = 0
+ moin = 5.5538
+ cgidl = 1
+ voffcv = -0.125
+ wpemod = 1
+ nigc = 2.291
+ ltvfbsdoff = 0
+ poxedge = 1
+ wkvth0we = 0.0
+ noff = 2.2684
+ binunit = 2
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ pbswd = 0.9
+ pbsws = 0.9
+ trnqsmod = 0
+ ntox = 1.0
+ pcit = -8.000000000000001e-19
+ pclm = 1.5514872
+ pdits = 0
+ cigsd = 0.013281
+ phin = 0.15
+ tpbswg = 0.001
+ ptvfbsdoff = 0
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ pkt1 = -4e-17
+ rgatemod = 0
+ tnjtsswg = 1
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ ptvoff = 0
+ rbdb = 50
+ prwb = 0
+ prwg = 0
+ tnoia = 0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ pvfbsdoff = 0
+ rdsw = 200
+ peta0 = -1.6e-17
+ diomod = 1
+ tpbsw = 0.0025
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.9113600000000002e-10
+ pku0we = 0.0
+ cjswgs = 1.9113600000000002e-10
+ cjswd = 5.3856e-11
+ a0 = 1.4508547
+ a1 = 0
+ a2 = 1
+ cjsws = 5.3856e-11
+ b0 = 0
+ b1 = 0
+ mjswd = 0.01
+ at = 72000
+ cf = 8.17e-11
+ mjsws = 0.01
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.013949949
+ k3 = -2.5823
+ agidl = 3.2166e-9
+ em = 20000000.0
+ ll = -1.18e-13
+ lw = 0
+ u0 = 0.009322119700000001
+ w0 = 0
+ ua = -3.1871506e-10
+ ub = 1.6925299e-18
+ uc = 2.1642376e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 3.4e-9
+ ags = 2.6576055
+ njtsswg = 6.489
+ mjswgd = 0.95
+ mjswgs = 0.95
+ cjd = 0.001421376
+ cit = 0.00044006838
+ cjs = 0.001421376
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ rshg = 14.1
+ bvs = 8.2
+ dlc = 1.38228675e-8
+ xtsswgd = 0.32
+ k3b = 2.1176
+ xtsswgs = 0.32
+ tcjswg = 0.00128
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.016932267
+ pdiblcb = 0
+ la0 = -4.2380342e-8
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0.00064
+ kt1 = -0.23958332
+ kt2 = -0.07162235
+ lk2 = 4.6255939e-9
+ scref = 1e-6
+ llc = -1.18e-13
+ lln = 0.7
+ lu0 = -1.8523925000000002e-10
+ mjd = 0.335
+ mjs = 0.335
+ lua = -2.581899e-17
+ lub = -2.6275812e-26
+ luc = -1.1293514e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ pigcd = 2.572
+ njd = 1.02
+ njs = 1.02
+ aigsd = 0.0063636407
+ pa0 = 0
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ pk2 = 0
+ pu0 = 0
+ prt = 0
+ pud = 0
+ tnom = 25
+ lvoff = -1.3382853e-9
+ rsh = 15.2
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ tcj = 0.000832
+ ua1 = 2.2510566e-9
+ ub1 = -2.8588123e-18
+ uc1 = 7.8974359e-11
+ bigbacc = 0.0054401
+ tpb = 0.0016
+ lvsat = 0.00085560684
+ ijthsfwd = 0.01
+ wa0 = 0
+ ute = -1
+ lvth0 = 4.9377832e-9
+ web = 6628.3
+ wec = -16935.0
+ fprout = 200
+ wk2 = 0
+ wlc = 0
+ wln = 1
+ wu0 = 0
+ xgl = -8.2e-9
+ xgw = 0
+ delta = 0.018814
+ wud = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ laigc = -2.0986759e-11
+ kvth0we = -0.00022
+ rnoia = 0
+ rnoib = 0
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ wtvoff = 0
+ vtsswgs = 1.1
+ ijthsrev = 0.01
+ ngate = 1.7e+20
+ wcit = 0.0
+ ngcon = 1
+ wpclm = 0
+ voff = -0.13301586
+ acde = 0.5
+ gbmin = 1e-12
+ capmod = 2
+ vsat = 115982.91
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ wint = 0
+ vth0 = -0.43136548
+ wku0we = 1.5e-11
+ wmax = 0.00090001
+ aigc = 0.0067688324
+ wmin = 9.0026e-6
+ mobmod = 0
+ ppdiblc2 = 0
+ bigc = 0.0012521
+ wwlc = 0
+ nfactor = 1
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ tvoff = 0.0018930751
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigc = 0.15259
+ xjbvd = 1
+ xjbvs = 1
+ pkvth0we = 0.0
+ lk2we = 0.0
+ vfbsdoff = 0.01
+ ku0we = -0.0007
+ nigbacc = 10
+ beta0 = 13.32
+ leta0 = -4.8e-10
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ ppclm = 0
+ paramchk = 1
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ nigbinv = 2.171
+ k2we = 5e-5
+ tvfbsdoff = 0.1
+ dsub = 0.5
+ dtox = 3.91e-10
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ eta0 = 0.1672
+ ijthdfwd = 0.01
+ etab = -0.23
+ toxref = 3e-9
+ fnoimod = 1
+ eigbinv = 1.1
+ bigsd = 0.0003327
+ ijthdrev = 0.01
+ wvfbsdoff = 0
+ wvoff = 0
+ lvfbsdoff = 0
+ ltvoff = -6.6370123e-11
+ lpdiblc2 = -1.4976331e-9
+ wvsat = 0.0
+ wvth0 = -2.1600000000000004e-9
+ cigbacc = 0.245
+ lku0we = 1.8e-11
+ lketa = 1.1808374e-9
+ tnoimod = 0
+ epsrox = 3.9
+ xpart = 1
+ rdsmod = 0
+ cigbinv = 0.006
+ egidl = 0.001
+ lkvth0we = 3e-12
+ igbmod = 1
+ )

.model pch_fs_6 pmos (
+ level = 54
+ wpclm = 0
+ vfbsdoff = 0.01
+ rshg = 14.1
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ nfactor = 1
+ wtvfbsdoff = 0
+ paramchk = 1
+ permod = 1
+ ltvfbsdoff = 0
+ tnom = 25
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ nigbacc = 10
+ ijthdfwd = 0.01
+ voffcv = -0.125
+ wpemod = 1
+ tvoff = 0.00091084129
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ nigbinv = 2.171
+ ptvfbsdoff = 0
+ ijthdrev = 0.01
+ wcit = 0.0
+ ku0we = -0.0007
+ lpdiblc2 = 0
+ voff = -0.11896044
+ beta0 = 13.32
+ acde = 0.5
+ leta0 = -1.5941465e-9
+ letab = 2.0255694e-8
+ vsat = 185878.73
+ wint = 0
+ vth0 = -0.36130292
+ ppclm = 0
+ tpbswg = 0.001
+ wmax = 0.00090001
+ fnoimod = 1
+ aigc = 0.0067067782
+ wmin = 9.0026e-6
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ eigbinv = 1.1
+ tvfbsdoff = 0.1
+ ptvoff = 0
+ lkvth0we = 3e-12
+ bigc = 0.0012521
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ wwlc = 0
+ diomod = 1
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ acnqsmod = 0
+ pditsd = 0
+ pditsl = 0
+ cgsl = 3.0105e-11
+ cjswgd = 1.9113600000000002e-10
+ pku0we = 0.0
+ cgso = 2.6482e-11
+ cigbacc = 0.245
+ cjswgs = 1.9113600000000002e-10
+ cigc = 0.15259
+ bigsd = 0.0003327
+ rbodymod = 0
+ wvfbsdoff = 0
+ tnoimod = 0
+ lvfbsdoff = 0
+ wvoff = 0
+ mjswgd = 0.95
+ mjswgs = 0.95
+ wvsat = 0.0
+ cigbinv = 0.006
+ wvth0 = -2.1600000000000004e-9
+ tcjswg = 0.00128
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ version = 4.5
+ lketa = 8.4925319e-9
+ k2we = 5e-5
+ tempmod = 0
+ wpdiblc2 = 0
+ xpart = 1
+ dsub = 0.5
+ dtox = 3.91e-10
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ egidl = 0.001
+ a0 = 3.4166667
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 140456.11
+ cf = 8.17e-11
+ aigbacc = 0.012071
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.010241786
+ k3 = -2.5823
+ em = 20000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.0053138889
+ w0 = 0
+ ua = -1.1682959e-9
+ ub = 1.3034444e-18
+ uc = -8.7638e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 3.4e-9
+ fprout = 200
+ eta0 = 0.17905262
+ etab = -0.44548611
+ xrcrg1 = 12
+ xrcrg2 = 1
+ aigbinv = 0.009974
+ wkvth0we = 0.0
+ wtvoff = 0
+ trnqsmod = 0
+ capmod = 2
+ pvoff = 2e-17
+ wku0we = 1.5e-11
+ cdscb = 0
+ cdscd = 0
+ mobmod = 0
+ pvsat = 0.0
+ wk2we = 0.0
+ pvth0 = -1.2e-16
+ drout = 0.56
+ poxedge = 1
+ rgatemod = 0
+ voffl = 0
+ tnjtsswg = 1
+ binunit = 2
+ weta0 = -2.2400000000000003e-10
+ lpclm = -9.8438889e-8
+ cgidl = 1
+ keta = -0.20642296
+ pbswd = 0.9
+ pbsws = 0.9
+ lags = -2.8753242e-8
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ lcit = 2.0151944e-10
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ kt1l = 0
+ pdits = 0
+ cigsd = 0.013281
+ lint = 0
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ lkt1 = -1.71119e-9
+ lkt2 = 1.5220167e-10
+ lmax = 9e-8
+ lmin = 5.4e-8
+ lpe0 = 6.44e-8
+ lpeb = 0
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ minv = -0.33
+ lua1 = -7.3062676e-18
+ lub1 = 1.0038041e-26
+ luc1 = 7.6176556e-18
+ ndep = 1e+18
+ toxref = 3e-9
+ njtsswg = 6.489
+ tnoia = 0
+ ijthsfwd = 0.01
+ lwlc = 0
+ pvfbsdoff = 0
+ moin = 5.5538
+ xtsswgd = 0.32
+ peta0 = -1.6e-17
+ xtsswgs = 0.32
+ nigc = 2.291
+ ckappad = 0.6
+ ckappas = 0.6
+ tpbsw = 0.0025
+ ags = 3.3058856
+ pdiblc1 = 0
+ pdiblc2 = 0.001
+ pdiblcb = 0
+ cjswd = 5.3856e-11
+ cjd = 0.001421376
+ cjsws = 5.3856e-11
+ cit = -0.00072561111
+ cjs = 0.001421376
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ dlc = 4.0349e-9
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ k3b = 2.1176
+ ijthsrev = 0.01
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ ltvoff = 2.5959859e-11
+ la0 = -2.2716667e-7
+ ntox = 1.0
+ pcit = -8.000000000000001e-19
+ jsd = 1.5e-7
+ pclm = 2.4472222
+ jss = 1.5e-7
+ lat = -0.0057948744
+ kt1 = -0.27692169
+ kt2 = -0.078859167
+ lk2 = 4.277026599999999e-9
+ llc = 0
+ lln = 1
+ lu0 = 1.9153444e-10
+ mjd = 0.335
+ bigbacc = 0.0054401
+ mjs = 0.335
+ lua = 5.4041604e-17
+ lub = 1.0298222e-26
+ luc = 9.143004e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 0
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ pk2 = 0
+ phin = 0.15
+ pu0 = 0
+ lku0we = 1.8e-11
+ prt = 0
+ pub = 0.0
+ pud = 0
+ kvth0we = -0.00022
+ epsrox = 3.9
+ ppdiblc2 = 0
+ rsh = 15.2
+ scref = 1e-6
+ pkt1 = -4e-17
+ tcj = 0.000832
+ ua1 = 7.2751825e-10
+ ub1 = -1.1117937e-18
+ uc1 = 7.4761111e-11
+ tpb = 0.0016
+ pigcd = 2.572
+ lintnoi = -5e-9
+ wa0 = 0
+ aigsd = 0.0063636407
+ ute = -1
+ web = 6628.3
+ wec = -16935.0
+ bigbinv = 0.00149
+ wk2 = 0
+ rdsmod = 0
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ wlc = 0
+ wln = 1
+ wu0 = 0
+ xgl = -8.2e-9
+ xgw = 0
+ wub = 0.0
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ igbmod = 1
+ lvoff = -2.6594942e-9
+ rbdb = 50
+ prwb = 0
+ prwg = 0
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ rbpb = 50
+ rbpd = 50
+ lvsat = -0.0057146009
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ lvth0 = -1.648097e-9
+ pbswgd = 0.8
+ pbswgs = 0.8
+ rdsw = 200
+ delta = 0.018814
+ laigc = -1.5153664e-11
+ igcmod = 1
+ rnoia = 0
+ rnoib = 0
+ pkvth0we = 0.0
+ ngate = 1.7e+20
+ ngcon = 1
+ )

.model pch_fs_7 pmos (
+ level = 54
+ voffl = 0
+ dsub = 0.5
+ dtox = 3.91e-10
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ weta0 = -2.2400000000000003e-10
+ ptvfbsdoff = 0
+ lpclm = -4.4240467e-8
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ eta0 = 0.18948293
+ ijthsfwd = 0.01
+ voffcv = -0.125
+ wpemod = 1
+ etab = -0.27185615
+ cgidl = 1
+ ijthsrev = 0.01
+ pbswd = 0.9
+ pbsws = 0.9
+ njtsswg = 6.489
+ tpbswg = 0.001
+ pdits = 0
+ cigsd = 0.013281
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ ppdiblc2 = 0
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.001
+ pdiblcb = 0
+ pk2we = 0.0
+ ptvoff = 0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ ags = 2.81014
+ pvfbsdoff = 0
+ tnoia = 0
+ diomod = 1
+ cjd = 0.001421376
+ cit = -0.0030912222
+ cjs = 0.001421376
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 4.0349e-9
+ peta0 = -1.6e-17
+ k3b = 2.1176
+ pditsd = 0
+ pditsl = 0
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ bigbacc = 0.0054401
+ dwj = 0
+ cjswgd = 1.9113600000000002e-10
+ pku0we = 0.0
+ cjswgs = 1.9113600000000002e-10
+ tpbsw = 0.0025
+ pkvth0we = 0.0
+ keta = 0.048888889
+ cjswd = 5.3856e-11
+ kvth0we = -0.00022
+ cjsws = 5.3856e-11
+ la0 = -1.5788889e-7
+ jsd = 1.5e-7
+ mjswd = 0.01
+ jss = 1.5e-7
+ lat = 0.0049061578
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ kt1 = -0.090229195
+ kt2 = -0.087042222
+ lk2 = 4.6553879e-9
+ llc = 0
+ lln = 1
+ lu0 = -7.3428889e-11
+ mjd = 0.335
+ mjs = 0.335
+ lua = -4.5270917e-17
+ lub = -1.9748742e-26
+ luc = -2.161341e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ lintnoi = -5e-9
+ njd = 1.02
+ mjswgd = 0.95
+ njs = 1.02
+ mjswgs = 0.95
+ pa0 = 0
+ bigbinv = 0.00149
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ jswd = 3.69e-13
+ vtsswgd = 1.1
+ pk2 = 0
+ jsws = 3.69e-13
+ vtsswgs = 1.1
+ vfbsdoff = 0.01
+ lcit = 3.3872489e-10
+ pu0 = 0
+ tcjswg = 0.00128
+ prt = 0
+ pub = 0.0
+ pud = 0
+ kt1l = 0
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 1.0031266e-9
+ ub1 = -2.5489021e-18
+ uc1 = 1.9738889e-10
+ tpb = 0.0016
+ wa0 = 0
+ ute = -1
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 0
+ lint = 0
+ wlc = 0
+ wln = 1
+ wu0 = 0
+ xgl = -8.2e-9
+ xgw = 0
+ paramchk = 1
+ wub = 0.0
+ wud = 0
+ wwc = 0
+ lkt1 = -1.2539355e-8
+ lkt2 = 6.2681889e-10
+ wwl = 0
+ wwn = 1
+ lmax = 5.4e-8
+ lmin = 4.5e-8
+ scref = 1e-6
+ lpe0 = 6.44e-8
+ lpeb = 0
+ pigcd = 2.572
+ aigsd = 0.0063636407
+ minv = -0.33
+ lvoff = -4.1866651e-9
+ lua1 = -2.3291554e-17
+ lub1 = 9.339033e-26
+ luc1 = 5.0524444e-19
+ fprout = 200
+ ndep = 1e+18
+ lvsat = -0.00013210428
+ ijthdfwd = 0.01
+ xrcrg1 = 12
+ xrcrg2 = 1
+ lwlc = 0
+ lvth0 = -2.5566339e-9
+ moin = 5.5538
+ delta = 0.018814
+ laigc = -9.9932362e-12
+ nigc = 2.291
+ nfactor = 1
+ rnoia = 0
+ rnoib = 0
+ wtvoff = 0
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ ijthdrev = 0.01
+ ngate = 1.7e+20
+ ngcon = 1
+ wpclm = 0
+ lpdiblc2 = 0
+ capmod = 2
+ ntox = 1.0
+ pcit = -8.000000000000001e-19
+ wku0we = 1.5e-11
+ pclm = 1.5127667
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ nigbacc = 10
+ a0 = 2.2222222
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = -44044.444
+ mobmod = 0
+ cf = 8.17e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.016765256
+ k3 = -2.5823
+ em = 20000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.0098822222
+ w0 = 0
+ ua = 5.4398899e-10
+ ub = 1.8214956e-18
+ uc = 4.42645e-10
+ ud = 0
+ phin = 0.15
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 3.4e-9
+ pkt1 = -4e-17
+ nigbinv = 2.171
+ lkvth0we = 3e-12
+ rbdb = 50
+ prwb = 0
+ prwg = 0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ rdsw = 200
+ tvoff = 0.0051729841
+ acnqsmod = 0
+ fnoimod = 1
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ eigbinv = 1.1
+ rbodymod = 0
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = -2.1991042999999997e-9
+ rshg = 14.1
+ letab = 1.0185157e-8
+ ppclm = 0
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ tvfbsdoff = 0.1
+ cigbacc = 0.245
+ wpdiblc2 = 0
+ tnoimod = 0
+ tnom = 25
+ dmcgt = 0
+ toxref = 3e-9
+ tcjsw = 9.34e-5
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ cigbinv = 0.006
+ bigsd = 0.0003327
+ wkvth0we = 0.0
+ version = 4.5
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ tempmod = 0
+ ltvoff = -2.2124443e-10
+ wvoff = 0
+ wcit = 0.0
+ trnqsmod = 0
+ voff = -0.092629909
+ wvsat = 0.0
+ acde = 0.5
+ wvth0 = -2.1600000000000004e-9
+ aigbacc = 0.012071
+ vsat = 89628.791
+ wint = 0
+ vth0 = -0.34563849
+ lku0we = 1.8e-11
+ wmax = 0.00090001
+ aigc = 0.0066178053
+ wmin = 9.0026e-6
+ epsrox = 3.9
+ lketa = -6.3155556e-9
+ rgatemod = 0
+ xpart = 1
+ aigbinv = 0.009974
+ tnjtsswg = 1
+ rdsmod = 0
+ igbmod = 1
+ egidl = 0.001
+ bigc = 0.0012521
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ wwlc = 0
+ pbswgd = 0.8
+ pbswgs = 0.8
+ cdsc = 0
+ cgbo = 0
+ igcmod = 1
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigc = 0.15259
+ wtvfbsdoff = 0
+ poxedge = 1
+ binunit = 2
+ ltvfbsdoff = 0
+ pvoff = 2e-17
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ cdscb = 0
+ cdscd = 0
+ pvsat = 0.0
+ wk2we = 0.0
+ pvth0 = -1.2e-16
+ drout = 0.56
+ permod = 1
+ k2we = 5e-5
+ )

.model pch_fs_8 pmos (
+ level = 54
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ wkvth0we = 0.0
+ cigbacc = 0.245
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ trnqsmod = 0
+ ku0we = -0.0007
+ tnoimod = 0
+ beta0 = 13.32
+ leta0 = 1.6523128000000001e-9
+ ntox = 1.0
+ letab = 3.9337702e-9
+ pcit = -8.000000000000001e-19
+ pclm = 1.0208333
+ tpbswg = 0.001
+ cigbinv = 0.006
+ ppclm = 0
+ phin = 0.15
+ dlcig = 2.5e-9
+ tvfbsdoff = 0.1
+ bgidl = 1834800000.0
+ pkt1 = -4e-17
+ rgatemod = 0
+ ptvoff = 0
+ tnjtsswg = 1
+ version = 4.5
+ tempmod = 0
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ diomod = 1
+ rbdb = 50
+ prwb = 0
+ prwg = 0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ aigbacc = 0.012071
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.9113600000000002e-10
+ pku0we = 0.0
+ cjswgs = 1.9113600000000002e-10
+ rdsw = 200
+ bigsd = 0.0003327
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ mjswgd = 0.95
+ mjswgs = 0.95
+ wvoff = 0
+ aigbinv = 0.009974
+ tcjswg = 0.00128
+ wvsat = 0.0
+ wvth0 = -2.1600000000000004e-9
+ rshg = 14.1
+ lketa = 8.0381778e-9
+ xpart = 1
+ poxedge = 1
+ egidl = 0.001
+ tnom = 25
+ fprout = 200
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ xrcrg1 = 12
+ xrcrg2 = 1
+ binunit = 2
+ ijthsfwd = 0.01
+ wtvoff = 0
+ ijthsrev = 0.01
+ wcit = 0.0
+ capmod = 2
+ voff = -0.10032114
+ wku0we = 1.5e-11
+ acde = 0.5
+ pvoff = 2e-17
+ mobmod = 0
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ vsat = 122520.32
+ wint = 0
+ vth0 = -0.39238557
+ cdscb = 0
+ cdscd = 0
+ wkt1 = 0.0
+ pvsat = 0.0
+ wmax = 0.00090001
+ wk2we = 0.0
+ pvth0 = -1.2e-16
+ aigc = 0.0065563017
+ wmin = 9.0026e-6
+ drout = 0.56
+ ppdiblc2 = 0
+ voffl = 0
+ weta0 = -2.2400000000000003e-10
+ wetab = 0
+ bigc = 0.0012521
+ wwlc = 0
+ lpclm = -2.0135733e-8
+ laigsd = -2.1777787e-18
+ cdsc = 0
+ cgidl = 1
+ njtsswg = 6.489
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigc = 0.15259
+ a0 = -0.19555556
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ xtsswgd = 0.32
+ pkvth0we = 0.0
+ xtsswgs = 0.32
+ at = 76220.0
+ cf = 8.17e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.012217534
+ k3 = -2.5823
+ em = 20000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.0053777778000000005
+ w0 = 0
+ ua = -1.1794951e-9
+ ub = 1.5005044e-18
+ uc = 5.0701667e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 3.4e-9
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.001
+ pbswd = 0.9
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ pbsws = 0.9
+ pdiblcb = 0
+ vfbsdoff = 0.01
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ pdits = 0
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ paramchk = 1
+ bigbacc = 0.0054401
+ k2we = 5e-5
+ ags = 1.0774289
+ dsub = 0.5
+ kvth0we = -0.00022
+ dtox = 3.91e-10
+ cjd = 0.001421376
+ cit = -0.00097166667
+ pk2we = 0.0
+ cjs = 0.001421376
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ dlc = 4.0349e-9
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ k3b = 2.1176
+ toxref = 3e-9
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ pvfbsdoff = 0
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ tnoia = 0
+ ijthdfwd = 0.01
+ eta0 = 0.11088258
+ etab = -0.14427684
+ la0 = -3.9417778e-8
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = -0.0009868
+ kt1 = -0.30391077
+ kt2 = -0.08425
+ lk2 = 4.432549499999999e-9
+ peta0 = -1.6e-17
+ llc = 0
+ lln = 1
+ lu0 = 1.4728888999999998e-10
+ petab = 0
+ mjd = 0.335
+ mjs = 0.335
+ lua = 3.9179804e-17
+ lub = -4.0201778e-27
+ luc = -2.4081867e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 0
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0.0
+ pbs = 0.75
+ tpbsw = 0.0025
+ pk2 = 0
+ pu0 = 0
+ prt = 0
+ pub = 0.0
+ pud = 0
+ cjswd = 5.3856e-11
+ cjsws = 5.3856e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ ltvoff = -2.4936809e-11
+ agidl = 3.2166e-9
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 1.4917512e-9
+ ub1 = -1.5908843e-18
+ uc1 = 1.6325556e-10
+ ijthdrev = 0.01
+ tpb = 0.0016
+ wa0 = 0
+ ute = -1
+ wat = 0.0
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 0
+ wlc = 0
+ wln = 1
+ lpdiblc2 = 0
+ wu0 = 0
+ xgl = -8.2e-9
+ xgw = 0
+ wub = 0.0
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ lku0we = 1.8e-11
+ epsrox = 3.9
+ nfactor = 1
+ scref = 1e-6
+ rdsmod = 0
+ pigcd = 2.572
+ aigsd = 0.0063636407
+ igbmod = 1
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ wtvfbsdoff = 0
+ lvoff = -3.8097951e-9
+ lkvth0we = 3e-12
+ pbswgd = 0.8
+ pbswgs = 0.8
+ lvsat = -0.0017437894
+ lvth0 = -2.66027058e-10
+ igcmod = 1
+ ltvfbsdoff = 0
+ delta = 0.018814
+ nigbacc = 10
+ laigc = -6.97956e-12
+ acnqsmod = 0
+ rnoia = 0
+ rnoib = 0
+ keta = -0.24404444
+ rbodymod = 0
+ ngate = 1.7e+20
+ lags = 8.4902844e-8
+ ngcon = 1
+ nigbinv = 2.171
+ wpclm = 0
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 2.3486667e-10
+ kt1l = 0
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ ptvfbsdoff = 0
+ lint = 0
+ permod = 1
+ lkt1 = -2.0689574e-9
+ lkt2 = 4.9e-10
+ lmax = 4.5e-8
+ lmin = 3.6e-8
+ fnoimod = 1
+ wpdiblc2 = 0
+ lpe0 = 6.44e-8
+ lpeb = 0
+ eigbinv = 1.1
+ minv = -0.33
+ lua1 = -4.7234158e-17
+ lub1 = 4.6447457e-26
+ luc1 = 2.1777778e-18
+ voffcv = -0.125
+ wpemod = 1
+ ndep = 1e+18
+ lwlc = 0
+ moin = 5.5538
+ tvoff = 0.0011667062
+ nigc = 2.291
+ )

.model pch_fs_9 pmos (
+ level = 54
+ vtsswgs = 1.1
+ ags = 0.82538676
+ vsat = 121084.96
+ wint = 0
+ vth0 = -0.40947733000000003
+ pdits = 0
+ cjd = 0.001421376
+ cit = 5e-6
+ cjs = 0.001421376
+ clc = 1e-7
+ cle = 0.6
+ cigsd = 0.013281
+ bvd = 8.2
+ bvs = 8.2
+ wkt1 = -1.0361455e-8
+ wkt2 = -3.8769913e-9
+ dlc = 1.0572421799999999e-8
+ wmax = 9.0026e-6
+ dvt0w = 0
+ k3b = 2.1176
+ dvt1w = 0
+ aigc = 0.0068303602
+ dvt2w = 0
+ wmin = 9.025999999999999e-7
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ ptvoff = 0
+ waigsd = 1.9139418e-12
+ la0 = 0
+ pk2we = 0.0
+ jsd = 1.5e-7
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ jss = 1.5e-7
+ lat = 0.00064
+ wua1 = -3.2799159e-16
+ kt1 = -0.16992583
+ lk2 = 3.2000000000000003e-10
+ kt2 = -0.04703951
+ wub1 = 5.9231251e-25
+ wuc1 = -8.7396626e-17
+ llc = 0
+ lln = 1
+ lu0 = -8e-13
+ mjd = 0.335
+ mjs = 0.335
+ lkvth0we = 3e-12
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ diomod = 1
+ pvfbsdoff = 0
+ njd = 1.02
+ bigc = 0.0012521
+ njs = 1.02
+ wute = -7.8572347e-8
+ pa0 = 0
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ wwlc = 0
+ pk2 = 0
+ tnoia = 0
+ pu0 = 0
+ pditsd = 0
+ pditsl = 0
+ prt = 0
+ pud = 0
+ cjswgd = 1.9113600000000002e-10
+ pku0we = 0.0
+ cjswgs = 1.9113600000000002e-10
+ rsh = 15.2
+ tcj = 0.000832
+ peta0 = -1.6e-17
+ cdsc = 0
+ ua1 = 1.2333536e-9
+ ub1 = -1.432383e-18
+ uc1 = 7.8434267e-11
+ cgbo = 0
+ tpb = 0.0016
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ acnqsmod = 0
+ xtid = 3
+ xtis = 3
+ wketa = 2.2362589e-8
+ wa0 = 3.3745816e-7
+ ute = -0.99127556
+ web = 6628.3
+ wec = -16935.0
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ wk2 = -2.287053e-9
+ tpbsw = 0.0025
+ cigc = 0.15259
+ wlc = 0
+ wln = 1
+ wu0 = -8.6631049e-11
+ xgl = -8.2e-9
+ xgw = 0
+ wua = -1.124189e-16
+ wub = -6.7100784e-26
+ wuc = -2.319496e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ cjswd = 5.3856e-11
+ nfactor = 1
+ cjsws = 5.3856e-11
+ mjswd = 0.01
+ mjswgd = 0.95
+ mjsws = 0.01
+ mjswgs = 0.95
+ agidl = 3.2166e-9
+ rbodymod = 0
+ tcjswg = 0.00128
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ nigbacc = 10
+ scref = 1e-6
+ k2we = 5e-5
+ wpdiblc2 = 3.6469361e-10
+ pigcd = 2.572
+ dsub = 0.5
+ aigsd = 0.0063633875
+ dtox = 3.91e-10
+ fprout = 200
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ lvoff = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ nigbinv = 2.171
+ lvsat = 8.000000000000001e-6
+ eta0 = 0.16744607
+ etab = -0.23671111
+ lvth0 = -2.4e-10
+ delta = 0.018814
+ wtvoff = -9.8925647e-11
+ rnoia = 0
+ rnoib = 0
+ wkvth0we = 0.0
+ fnoimod = 1
+ ngate = 1.7e+20
+ capmod = 2
+ trnqsmod = 0
+ eigbinv = 1.1
+ ngcon = 1
+ wpclm = -3.01194e-7
+ wku0we = 1.5e-11
+ mobmod = 0
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ rgatemod = 0
+ tnjtsswg = 1
+ cigbacc = 0.245
+ tnoimod = 0
+ tvoff = 0.0026265487
+ cigbinv = 0.006
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ keta = -0.044833188
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ version = 4.5
+ jswd = 3.69e-13
+ ku0we = -0.0007
+ jsws = 3.69e-13
+ lcit = 1.6e-11
+ tempmod = 0
+ beta0 = 13.32
+ leta0 = -4.8e-10
+ kt1l = 0
+ ppclm = 0
+ aigbacc = 0.012071
+ lint = 6.5375218e-9
+ tvfbsdoff = 0.1
+ dlcig = 2.5e-9
+ lkt1 = -4.8e-10
+ bgidl = 1834800000.0
+ lmax = 2.001e-5
+ lmin = 8.9991e-6
+ lpe0 = 6.44e-8
+ lpeb = 0
+ a0 = 2.4935296
+ a1 = 0
+ a2 = 1
+ toxref = 3e-9
+ b0 = 0
+ b1 = 0
+ at = 72000
+ cf = 8.17e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.00052197993
+ k3 = -2.5823
+ em = 20000000.0
+ aigbinv = 0.009974
+ minv = -0.33
+ ll = 0
+ lw = 0
+ u0 = 0.0098846193
+ w0 = 0
+ ua = 1.4218267e-10
+ ub = 1.1900227e-18
+ uc = 2.2715501e-11
+ ud = 0
+ dmcgt = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 3.4e-9
+ tcjsw = 9.34e-5
+ ndep = 1e+18
+ ijthsfwd = 0.01
+ lwlc = 0
+ moin = 5.5538
+ nigc = 2.291
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ bigsd = 0.0003327
+ ltvoff = 0
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ ijthsrev = 0.01
+ wvoff = 5.5905393e-9
+ poxedge = 1
+ wvsat = -0.0097711764
+ wvth0 = 9.205859999999996e-10
+ ntox = 1.0
+ pcit = -8.000000000000001e-19
+ pclm = 1.5174437
+ binunit = 2
+ lku0we = 1.8e-11
+ wtvfbsdoff = 0
+ waigc = 3.5172206e-12
+ epsrox = 3.9
+ phin = 0.15
+ lketa = 0
+ rdsmod = 0
+ ltvfbsdoff = 0
+ ppdiblc2 = 0
+ pkt1 = -4e-17
+ xpart = 1
+ igbmod = 1
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ egidl = 0.001
+ pbswgd = 0.8
+ pbswgs = 0.8
+ rbdb = 50
+ prwb = 0
+ prwg = 0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ igcmod = 1
+ rbsb = 50
+ pvag = 2.1
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ rdsw = 200
+ ptvfbsdoff = 0
+ pkvth0we = 0.0
+ vfbsdoff = 0.01
+ rshg = 14.1
+ pvoff = 2e-17
+ cdscb = 0
+ cdscd = 0
+ permod = 1
+ pvsat = 0
+ wk2we = 0.0
+ pvth0 = -1.2e-16
+ paramchk = 1
+ njtsswg = 6.489
+ drout = 0.56
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ voffl = 0
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.0026324684
+ weta0 = -2.4401431e-9
+ tnom = 25
+ pdiblcb = 0
+ wetab = 6.0440267e-8
+ voffcv = -0.125
+ wpemod = 1
+ lpclm = 0
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ ijthdfwd = 0.01
+ cgidl = 1
+ bigbacc = 0.0054401
+ wags = 1.128996e-7
+ ijthdrev = 0.01
+ pbswd = 0.9
+ pbsws = 0.9
+ kvth0we = -0.00022
+ lpdiblc2 = 0
+ voff = -0.11172412
+ tpbswg = 0.001
+ acde = 0.5
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ )

.model pch_fs_10 pmos (
+ level = 54
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ lags = 3.1017116e-7
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 1.6e-11
+ nfactor = 1
+ kt1l = 0
+ paramchk = 1
+ scref = 1e-6
+ pigcd = 2.572
+ aigsd = 0.0063633879
+ lint = 6.5375218e-9
+ lkt1 = -4.2387452e-8
+ lkt2 = -8.3161855e-9
+ lmax = 8.9991e-6
+ lvoff = -7.1040424e-9
+ lmin = 8.9908e-7
+ lpe0 = 6.44e-8
+ lpeb = 0
+ lvsat = 8.000000000000001e-6
+ lvth0 = -4.7217588e-9
+ ijthdfwd = 0.01
+ toxref = 3e-9
+ nigbacc = 10
+ minv = -0.33
+ delta = 0.018814
+ lua1 = 2.9697696e-17
+ lub1 = 1.2607181e-25
+ luc1 = -4.744495e-18
+ laigc = -4.752933e-11
+ wtvfbsdoff = 0
+ ndep = 1e+18
+ rnoia = 0
+ rnoib = 0
+ lute = -8.6179201e-9
+ lwlc = 0
+ tvfbsdoff = 0.1
+ moin = 5.5538
+ ltvfbsdoff = 0
+ pketa = -2.2807538e-14
+ nigc = 2.291
+ ngate = 1.7e+20
+ ijthdrev = 0.01
+ nigbinv = 2.171
+ ngcon = 1
+ wpclm = -3.01194e-7
+ lpdiblc2 = 7.3300428e-9
+ ltvoff = -4.2514859e-10
+ gbmin = 1e-12
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ pags = -3.4942959e-14
+ ntox = 1.0
+ pcit = -8.000000000000001e-19
+ pclm = 1.5174437
+ fnoimod = 1
+ wvfbsdoff = 0
+ lku0we = 1.8e-11
+ ptvfbsdoff = 0
+ eigbinv = 1.1
+ lvfbsdoff = 0
+ epsrox = 3.9
+ phin = 0.15
+ lkvth0we = 3e-12
+ pkt1 = 8.9789586e-15
+ pkt2 = -4.3236504e-15
+ rdsmod = 0
+ igbmod = 1
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ tvoff = 0.0026738399
+ pbswgd = 0.8
+ acnqsmod = 0
+ pbswgs = 0.8
+ rbdb = 50
+ pua1 = 9.6044121e-22
+ prwb = 0
+ pub1 = -1.3952204e-30
+ prwg = 0
+ puc1 = 1.1914589e-22
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ pute = 7.7612988e-14
+ igcmod = 1
+ cigbacc = 0.245
+ rdsw = 200
+ rbodymod = 0
+ tnoimod = 0
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = -4.8e-10
+ cigbinv = 0.006
+ ppclm = 0
+ paigsd = 3.3403436e-20
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ rshg = 14.1
+ version = 4.5
+ wpdiblc2 = 5.6393415e-10
+ permod = 1
+ tempmod = 0
+ ags = 0.79088496
+ dmcgt = 0
+ cjd = 0.001421376
+ cit = 5e-6
+ cjs = 0.001421376
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ tcjsw = 9.34e-5
+ dlc = 1.0572421799999999e-8
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ aigbacc = 0.012071
+ tnom = 25
+ la0 = -3.6651331e-7
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ jsd = 1.5e-7
+ voffcv = -0.125
+ wpemod = 1
+ jss = 1.5e-7
+ lat = 0.00064
+ kt1 = -0.16526426
+ kt2 = -0.046114462
+ lk2 = 4.8245047999999995e-9
+ llc = 0
+ lln = 1
+ bigsd = 0.0003327
+ lu0 = -1.2024212000000002e-10
+ mjd = 0.335
+ mjs = 0.335
+ lua = -1.1601528e-16
+ lub = 1.1870612e-25
+ luc = 1.7407612e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = -2.3980423e-13
+ wkvth0we = 0.0
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ pk2 = -1.7678537e-15
+ aigbinv = 0.009974
+ wvoff = 6.4925381e-9
+ pu0 = 1.0845918e-15
+ prt = 0
+ pua = 1.4359661e-22
+ pub = 1.4495718e-31
+ puc = -1.3724663e-23
+ pud = 0
+ trnqsmod = 0
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 1.2300502e-9
+ ub1 = -1.4464065e-18
+ uc1 = 7.8962019e-11
+ wvsat = -0.0097711764
+ tpb = 0.0016
+ wvth0 = 1.5667411999999999e-9
+ wa0 = 3.6413271e-7
+ ute = -0.99031694
+ wags = 1.1678647e-7
+ web = 6628.3
+ wec = -16935.0
+ wk2 = -2.0904063e-9
+ wlc = 0
+ wln = 1
+ wu0 = -2.0727529e-10
+ xgl = -8.2e-9
+ waigc = 4.3868453e-12
+ xgw = 0
+ wua = -1.2839182e-16
+ wub = -8.3225053e-26
+ wuc = -2.1668301e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ voff = -0.11093391
+ acde = 0.5
+ tpbswg = 0.001
+ lketa = -1.0921036e-8
+ vsat = 121084.96
+ wint = 0
+ xpart = 1
+ vth0 = -0.40897880000000003
+ rgatemod = 0
+ wkt1 = -1.1364676e-8
+ wkt2 = -3.3960513e-9
+ poxedge = 1
+ wmax = 9.0026e-6
+ tnjtsswg = 1
+ aigc = 0.0068356471
+ wmin = 9.025999999999999e-7
+ egidl = 0.001
+ binunit = 2
+ ptvoff = -4.5667618e-16
+ waigsd = 1.9102262e-12
+ wua1 = -4.3482598e-16
+ wub1 = 7.4750944e-25
+ wuc1 = -1.0064978e-16
+ bigc = 0.0012521
+ wute = -8.7205605e-8
+ diomod = 1
+ wwlc = 0
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.9113600000000002e-10
+ pku0we = 0.0
+ cjswgs = 1.9113600000000002e-10
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigc = 0.15259
+ pvoff = -8.088969200000001e-15
+ jtsswgd = 1.75e-7
+ pvfbsdoff = 0
+ mjswgd = 0.95
+ jtsswgs = 1.75e-7
+ mjswgs = 0.95
+ cdscb = 0
+ cdscd = 0
+ tcjswg = 0.00128
+ pvsat = 0
+ wk2we = 0.0
+ pvth0 = -5.9289351000000005e-15
+ drout = 0.56
+ paigc = -7.8179264e-18
+ a0 = 2.5342986
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 72000
+ cf = 8.17e-11
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.0010230372
+ k3 = -2.5823
+ em = 20000000.0
+ voffl = 0
+ ll = 0
+ lw = 0
+ u0 = 0.0098979054
+ w0 = 0
+ ua = 1.5508759e-10
+ ub = 1.1768184e-18
+ uc = 2.077917e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 3.4e-9
+ weta0 = -2.4401431e-9
+ wetab = 6.0440267e-8
+ k2we = 5e-5
+ lpclm = 0
+ dsub = 0.5
+ dtox = 3.91e-10
+ ijthsfwd = 0.01
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ njtsswg = 6.489
+ cgidl = 1
+ fprout = 200
+ xrcrg1 = 12
+ xrcrg2 = 1
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ eta0 = 0.16744607
+ etab = -0.23671111
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.0018171133
+ pdiblcb = 0
+ pbswd = 0.9
+ wtvoff = -4.8127407e-11
+ pbsws = 0.9
+ ijthsrev = 0.01
+ pdits = 0
+ capmod = 2
+ cigsd = 0.013281
+ wku0we = 1.5e-11
+ bigbacc = 0.0054401
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ mobmod = 0
+ ppdiblc2 = -1.7911725e-15
+ kvth0we = -0.00022
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ tnoia = 0
+ peta0 = -1.6e-17
+ wketa = 2.4899578e-8
+ laigsd = -3.7090202e-15
+ tpbsw = 0.0025
+ pkvth0we = 0.0
+ cjswd = 5.3856e-11
+ cjsws = 5.3856e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ keta = -0.04361839
+ vfbsdoff = 0.01
+ )

.model pch_fs_11 pmos (
+ level = 54
+ egidl = 0.001
+ ltvfbsdoff = 0
+ toxref = 3e-9
+ ijthsfwd = 0.01
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ tnom = 25
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ ijthsrev = 0.01
+ ptvfbsdoff = 0
+ ltvoff = -2.603747e-10
+ pvfbsdoff = 0
+ wags = -5.7105665e-9
+ pvoff = 6.0710934e-15
+ cdscb = 0
+ cdscd = 0
+ pvsat = 0
+ wk2we = 0.0
+ voff = -0.10782222
+ njtsswg = 6.489
+ pvth0 = 3.1263808e-15
+ drout = 0.56
+ acde = 0.5
+ paigc = 1.0166993e-17
+ lku0we = 1.8e-11
+ xtsswgd = 0.32
+ vsat = 121084.96
+ xtsswgs = 0.32
+ wint = 0
+ ppdiblc2 = 8.932051e-16
+ vth0 = -0.41047369
+ epsrox = 3.9
+ voffl = 0
+ wkt1 = 3.9882501e-9
+ wkt2 = -1.3862366e-8
+ ckappad = 0.6
+ wmax = 9.0026e-6
+ ckappas = 0.6
+ aigc = 0.0068328167
+ wmin = 9.025999999999999e-7
+ pdiblc1 = 0
+ pdiblc2 = 0.0082016634
+ pdiblcb = 0
+ weta0 = -2.4401431e-9
+ rdsmod = 0
+ wetab = 6.0440267e-8
+ igbmod = 1
+ lpclm = 0
+ wua1 = 1.0350058e-15
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ wub1 = -1.41997e-24
+ wuc1 = 5.1522417e-17
+ cgidl = 1
+ pbswgd = 0.8
+ bigc = 0.0012521
+ pbswgs = 0.8
+ wwlc = 0
+ bigbacc = 0.0054401
+ igcmod = 1
+ pkvth0we = 0.0
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ pbswd = 0.9
+ pbsws = 0.9
+ kvth0we = -0.00022
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigc = 0.15259
+ vfbsdoff = 0.01
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ pdits = 0
+ cigsd = 0.013281
+ paigsd = -3.7089273e-20
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ paramchk = 1
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ permod = 1
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ k2we = 5e-5
+ tnoia = 0
+ dsub = 0.5
+ dtox = 3.91e-10
+ ijthdfwd = 0.01
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ peta0 = -1.6e-17
+ voffcv = -0.125
+ wpemod = 1
+ wketa = -2.3248862e-8
+ tpbsw = 0.0025
+ eta0 = 0.16744607
+ nfactor = 1
+ etab = -0.23671111
+ cjswd = 5.3856e-11
+ cjsws = 5.3856e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ ijthdrev = 0.01
+ lpdiblc2 = 1.6477933e-9
+ nigbacc = 10
+ tpbswg = 0.001
+ scref = 1e-6
+ pigcd = 2.572
+ aigsd = 0.0063633394
+ lvoff = -9.8734428e-9
+ nigbinv = 2.171
+ ptvoff = 2.6240046e-16
+ lkvth0we = 3e-12
+ waigsd = 1.9894315e-12
+ lvsat = 8.000000000000001e-6
+ lvth0 = -3.3913088e-9
+ delta = 0.018814
+ diomod = 1
+ laigc = -4.5010295e-11
+ acnqsmod = 0
+ rnoia = 0
+ rnoib = 0
+ tvfbsdoff = 0.1
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.9113600000000002e-10
+ pku0we = 0.0
+ cjswgs = 1.9113600000000002e-10
+ fnoimod = 1
+ pketa = 2.0044574e-14
+ rbodymod = 0
+ ngate = 1.7e+20
+ eigbinv = 1.1
+ ngcon = 1
+ wpclm = -3.01194e-7
+ keta = -0.035478054
+ mjswgd = 0.95
+ mjswgs = 0.95
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ tcjswg = 0.00128
+ lags = 2.7680102e-7
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 9.8671111e-11
+ kt1l = 0
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ wpdiblc2 = -2.4522204e-9
+ lint = 6.5375218e-9
+ cigbacc = 0.245
+ lkt1 = -1.5002155e-8
+ lkt2 = -7.1896716e-9
+ lmax = 8.9908e-7
+ lmin = 4.4908e-7
+ tnoimod = 0
+ lpe0 = 6.44e-8
+ lpeb = 0
+ fprout = 200
+ minv = -0.33
+ cigbinv = 0.006
+ lua1 = 8.7159171e-17
+ lub1 = -2.6689299e-25
+ luc1 = 2.9116076e-17
+ tvoff = 0.0024887007
+ xrcrg1 = 12
+ xrcrg2 = 1
+ ndep = 1e+18
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ lwlc = 0
+ moin = 5.5538
+ wkvth0we = 0.0
+ wtvoff = -8.5607868e-10
+ nigc = 2.291
+ version = 4.5
+ a0 = 2.8862723
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ trnqsmod = 0
+ at = 72000
+ cf = 8.17e-11
+ tempmod = 0
+ ef = 1.15
+ ku0we = -0.0007
+ k1 = 0.30425
+ k2 = 0.0046668319
+ k3 = -2.5823
+ em = 20000000.0
+ ll = 0
+ lw = 0
+ beta0 = 13.32
+ u0 = 0.0098844338
+ w0 = 0
+ ua = 8.4190146e-11
+ ub = 1.1838278e-18
+ uc = 4.9200634e-11
+ ud = 0
+ leta0 = -4.8e-10
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 3.4e-9
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ capmod = 2
+ ppclm = 0
+ aigbacc = 0.012071
+ wku0we = 1.5e-11
+ pags = 7.4079401e-14
+ ags = 0.8283795
+ dlcig = 2.5e-9
+ mobmod = 0
+ bgidl = 1834800000.0
+ ntox = 1.0
+ pcit = -8.000000000000001e-19
+ pclm = 1.5174437
+ cjd = 0.001421376
+ cit = -8.7888889e-5
+ cjs = 0.001421376
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 1.0572421799999999e-8
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ rgatemod = 0
+ tnjtsswg = 1
+ phin = 0.15
+ aigbinv = 0.009974
+ dmcgt = 0
+ la0 = -6.797699e-7
+ pkt1 = -4.6851461e-15
+ jsd = 1.5e-7
+ pkt2 = 4.9913693e-15
+ tcjsw = 9.34e-5
+ jss = 1.5e-7
+ lat = 0.00064
+ kt1 = -0.19603426
+ kt2 = -0.047380208
+ lk2 = -2.394787e-10
+ llc = 0
+ lln = 1
+ lu0 = -1.0825246e-10
+ mjd = 0.335
+ mjs = 0.335
+ lua = -5.2916554e-17
+ lub = 1.1246778e-25
+ luc = -7.8874906e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 4.0323955e-14
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ pk2 = 1.1838025e-15
+ pu0 = -8.8186737e-16
+ laigsd = 3.9492818e-14
+ prt = 0
+ pua = -2.1071339e-22
+ pub = -4.1382897e-32
+ puc = 1.6409308e-23
+ pud = 0
+ rbdb = 50
+ pua1 = -3.4770908e-22
+ prwb = 0
+ pub1 = 5.3383631e-31
+ prwg = 0
+ rsh = 15.2
+ puc1 = -1.6287371e-23
+ tcj = 0.000832
+ ua1 = 1.1654868e-9
+ ub1 = -1.004873e-18
+ uc1 = 4.0916434e-11
+ bigsd = 0.0003327
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ tpb = 0.0016
+ wa0 = 4.9381936e-8
+ ute = -1
+ web = 6628.3
+ wec = -16935.0
+ wk2 = -5.406874e-9
+ rdsw = 200
+ wlc = 0
+ wln = 1
+ wu0 = 2.0022293e-9
+ xgl = -8.2e-9
+ wvoff = -9.4176445e-9
+ xgw = 0
+ wua = 2.6970929e-16
+ wub = 1.2614582e-25
+ wuc = -5.5526695e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ poxedge = 1
+ wvsat = -0.0097711764
+ wvth0 = -8.6077711e-9
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ binunit = 2
+ waigc = -1.5820929e-11
+ rshg = 14.1
+ lketa = -1.8165935e-8
+ xpart = 1
+ wtvfbsdoff = 0
+ )

.model pch_fs_12 pmos (
+ level = 54
+ wkvth0we = 0.0
+ pketa = 2.9922765e-15
+ ngate = 1.7e+20
+ ngcon = 1
+ cigbacc = 0.245
+ ltvoff = -1.0992228e-10
+ wpclm = -3.01194e-7
+ trnqsmod = 0
+ gbmin = 1e-12
+ tnoimod = 0
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ cigbinv = 0.006
+ lku0we = 1.8e-11
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ epsrox = 3.9
+ rgatemod = 0
+ tnjtsswg = 1
+ rdsmod = 0
+ version = 4.5
+ igbmod = 1
+ tempmod = 0
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ pbswgd = 0.8
+ pbswgs = 0.8
+ tvoff = 0.0021467634
+ aigbacc = 0.012071
+ igcmod = 1
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ ku0we = -0.0007
+ ags = 0.29253015
+ aigbinv = 0.009974
+ beta0 = 13.32
+ keta = -0.031086208
+ leta0 = -4.8e-10
+ cjd = 0.001421376
+ cit = -0.00056559017
+ cjs = 0.001421376
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 1.38228675e-8
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ lags = 5.1257474e-7
+ ppclm = 0
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 3.0885967e-10
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ kt1l = 0
+ la0 = -1.4357692e-8
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0.00064
+ kt1 = -0.19916819
+ kt2 = -0.054700402
+ lk2 = 1.7450990000000002e-9
+ permod = 1
+ llc = -1.18e-13
+ lln = 0.7
+ lu0 = -4.815604500000001e-10
+ mjd = 0.335
+ mjs = 0.335
+ lua = -1.6078561e-16
+ lub = 5.7693033e-26
+ luc = -4.8483261e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ lint = 9.7879675e-9
+ pa0 = -2.613694e-13
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ pk2 = -5.5906497e-16
+ lkt1 = -1.3623224e-8
+ lkt2 = -3.9687861e-9
+ pu0 = -2.2461433e-17
+ lmax = 4.4908e-7
+ prt = 0
+ pua = 5.4100623e-23
+ pub = -6.3187687e-32
+ puc = -3.6550877e-24
+ pud = 0
+ dmcgt = 0
+ lmin = 2.1577e-7
+ poxedge = 1
+ tcjsw = 9.34e-5
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 1.2176874e-9
+ ub1 = -1.2376668e-18
+ lpe0 = 6.44e-8
+ uc1 = 1.0272662e-10
+ lpeb = 0
+ tpb = 0.0016
+ wa0 = 7.3504866e-7
+ ijthsfwd = 0.01
+ ute = -1
+ web = 6628.3
+ wec = -16935.0
+ wk2 = -1.4458115e-9
+ binunit = 2
+ voffcv = -0.125
+ wpemod = 1
+ wlc = 0
+ wln = 1
+ minv = -0.33
+ wu0 = 4.9034036e-11
+ xgl = -8.2e-9
+ xgw = 0
+ lua1 = 6.4190903e-17
+ lub1 = -1.6446372e-25
+ wua = -3.3214073e-16
+ wub = 1.7570216e-25
+ wuc = -9.9257962e-18
+ wud = 0
+ luc1 = 1.9195943e-18
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ ndep = 1e+18
+ bigsd = 0.0003327
+ lwlc = 0
+ moin = 5.5538
+ wvoff = 6.3544834e-9
+ nigc = 2.291
+ ijthsrev = 0.01
+ wvsat = -0.0097711764
+ wvth0 = -1.7487296100000003e-9
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ waigc = 4.9938134e-12
+ tpbswg = 0.001
+ jtsswgd = 1.75e-7
+ pags = 2.5662868e-13
+ jtsswgs = 1.75e-7
+ ntox = 1.0
+ pcit = -8.2477938e-17
+ lketa = -2.0098347e-8
+ pclm = 1.5174437
+ xpart = 1
+ ppdiblc2 = -1.9289508e-16
+ phin = 0.15
+ ptvoff = -6.733506e-17
+ egidl = 0.001
+ waigsd = 1.9051377e-12
+ pkt1 = 4.5381461e-16
+ pkt2 = -1.2251691e-15
+ diomod = 1
+ pditsd = 0
+ pditsl = 0
+ rbdb = 50
+ cjswgd = 1.9113600000000002e-10
+ pku0we = 0.0
+ pua1 = -4.1586322e-23
+ prwb = 0
+ pub1 = 2.600258e-32
+ prwg = 0
+ cjswgs = 1.9113600000000002e-10
+ puc1 = -8.5761835e-25
+ njtsswg = 6.489
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ pkvth0we = 0.0
+ rdsw = 200
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ ckappad = 0.6
+ ckappas = 0.6
+ mjswgd = 0.95
+ mjswgs = 0.95
+ pdiblc1 = 0
+ pdiblc2 = 0.01380092
+ pvfbsdoff = 0
+ pdiblcb = 0
+ vfbsdoff = 0.01
+ pvoff = -8.686429e-16
+ tcjswg = 0.00128
+ cdscb = 0
+ cdscd = 0
+ pvsat = 0
+ wk2we = 0.0
+ pvth0 = 1.0840255e-16
+ drout = 0.56
+ paramchk = 1
+ rshg = 14.1
+ paigc = 1.0085061e-18
+ bigbacc = 0.0054401
+ voffl = 0
+ weta0 = -2.4401431e-9
+ kvth0we = -0.00022
+ wetab = 6.0440267e-8
+ lpclm = 0
+ lintnoi = -5e-9
+ fprout = 200
+ ijthdfwd = 0.01
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ xrcrg1 = 12
+ xrcrg2 = 1
+ cgidl = 1
+ tnom = 25
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ wtvoff = -1.0667978e-10
+ pbswd = 0.9
+ pbsws = 0.9
+ ijthdrev = 0.01
+ lpdiblc2 = -8.1587971e-10
+ capmod = 2
+ wags = -4.2059528e-7
+ wku0we = 1.5e-11
+ wcit = 1.8563168e-10
+ pdits = 0
+ cigsd = 0.013281
+ mobmod = 0
+ voff = -0.12166106
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ acde = 0.5
+ vsat = 121084.96
+ wint = 0
+ vth0 = -0.42744281
+ nfactor = 1
+ pk2we = 0.0
+ wkt1 = -7.6912059e-9
+ wkt2 = 2.6613072e-10
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ wmax = 9.0026e-6
+ aigc = 0.0067878654
+ wmin = 9.025999999999999e-7
+ lkvth0we = 3e-12
+ tnoia = 0
+ a0 = 1.3739719
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 72000
+ wua1 = 3.3927227e-16
+ cf = 8.17e-11
+ wub1 = -2.6580249e-25
+ wuc1 = 1.6454797e-17
+ ef = 1.15
+ k1 = 0.30425
+ k2 = 0.00015642806
+ k3 = -2.5823
+ em = 20000000.0
+ peta0 = -1.6e-17
+ ll = -1.18e-13
+ lw = 0
+ u0 = 0.010732861
+ w0 = 0
+ ua = 3.293471e-10
+ ub = 1.3083159e-18
+ uc = 4.2293442e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ bigc = 0.0012521
+ xw = 3.4e-9
+ wketa = 1.5506359e-8
+ wwlc = 0
+ acnqsmod = 0
+ tpbsw = 0.0025
+ nigbacc = 10
+ cjswd = 5.3856e-11
+ cjsws = 5.3856e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ cdsc = 0
+ cgbo = 0
+ rbodymod = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigc = 0.15259
+ wtvfbsdoff = 0
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ nigbinv = 2.171
+ ltvfbsdoff = 0
+ scref = 1e-6
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ pigcd = 2.572
+ wpdiblc2 = 1.6189099e-11
+ aigsd = 0.0063634291
+ fnoimod = 1
+ lvoff = -3.7843526e-9
+ eigbinv = 1.1
+ k2we = 5e-5
+ toxref = 3e-9
+ lvsat = 8.000000000000001e-6
+ dsub = 0.5
+ dtox = 3.91e-10
+ lvth0 = 4.0751043e-9
+ ptvfbsdoff = 0
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ delta = 0.018814
+ laigc = -2.5231709e-11
+ tvfbsdoff = 0.1
+ rnoia = 0
+ rnoib = 0
+ eta0 = 0.16744607
+ etab = -0.23671111
+ )

.model pch_fs_13 pmos (
+ level = 54
+ pags = 7.0037917e-14
+ lku0we = 1.8e-11
+ pvth0 = -8.4768891e-16
+ drout = 0.56
+ epsrox = 3.9
+ ntox = 1.0
+ pcit = 3.0450046e-17
+ pclm = 1.5924795
+ paigc = -7.3857349e-19
+ voffl = 0
+ rdsmod = 0
+ phin = 0.15
+ igbmod = 1
+ weta0 = -2.4401431e-9
+ wetab = 6.0440267e-8
+ lkvth0we = 3e-12
+ pkt1 = 2.4071967e-16
+ pkt2 = -8.6151083e-16
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ lpclm = -1.5832542e-8
+ pbswgd = 0.8
+ pbswgs = 0.8
+ cgidl = 1
+ igcmod = 1
+ acnqsmod = 0
+ rbdb = 50
+ pua1 = -5.7774504e-23
+ prwb = 0
+ pub1 = 1.0356474e-31
+ prwg = 0
+ puc1 = 6.0450908e-24
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ rdsw = 200
+ rbodymod = 0
+ pbswd = 0.9
+ pbsws = 0.9
+ nfactor = 1
+ pdits = 0
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ permod = 1
+ rshg = 14.1
+ nigbacc = 10
+ wpdiblc2 = -2.9527442e-9
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ tnoia = 0
+ voffcv = -0.125
+ wpemod = 1
+ nigbinv = 2.171
+ peta0 = -1.6e-17
+ tnom = 25
+ wketa = 2.8638443e-8
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ tpbsw = 0.0025
+ cjswd = 5.3856e-11
+ cjsws = 5.3856e-11
+ mjswd = 0.01
+ wkvth0we = 0.0
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ trnqsmod = 0
+ fnoimod = 1
+ eigbinv = 1.1
+ wags = 4.6372111e-7
+ tpbswg = 0.001
+ wcit = -3.4957204e-10
+ voff = -0.13366619
+ acde = 0.5
+ scref = 1e-6
+ vsat = 116618.55
+ wint = 0
+ vth0 = -0.43191428000000004
+ rgatemod = 0
+ pigcd = 2.572
+ aigsd = 0.0063634291
+ wkt1 = -6.6812774e-9
+ wkt2 = -1.4573681e-9
+ tnjtsswg = 1
+ ptvoff = -1.8786066e-17
+ wmax = 9.0026e-6
+ aigc = 0.0067673585
+ wmin = 9.025999999999999e-7
+ lvoff = -1.2512704e-9
+ waigsd = 1.9051377e-12
+ cigbacc = 0.245
+ lvsat = 0.0009504132299999999
+ diomod = 1
+ lvth0 = 5.0185836e-9
+ wua1 = 4.1599351e-16
+ wub1 = -6.3339564e-25
+ wuc1 = -1.6259465e-17
+ tnoimod = 0
+ delta = 0.018814
+ laigc = -2.090475e-11
+ pditsd = 0
+ pditsl = 0
+ tvfbsdoff = 0.1
+ bigc = 0.0012521
+ cjswgd = 1.9113600000000002e-10
+ pku0we = 0.0
+ cjswgs = 1.9113600000000002e-10
+ wwlc = 0
+ rnoia = 0
+ rnoib = 0
+ cigbinv = 0.006
+ cdsc = 0
+ pketa = 2.2140676e-16
+ ngate = 1.7e+20
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ ngcon = 1
+ mjswgd = 0.95
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ mjswgs = 0.95
+ wpclm = -3.6917638e-7
+ cigc = 0.15259
+ tcjswg = 0.00128
+ version = 4.5
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ tempmod = 0
+ jswgs = 3.69e-13
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ aigbacc = 0.012071
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ k2we = 5e-5
+ fprout = 200
+ aigbinv = 0.009974
+ dsub = 0.5
+ dtox = 3.91e-10
+ xrcrg1 = 12
+ xrcrg2 = 1
+ ijthsfwd = 0.01
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ tvoff = 0.0019304691
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ ags = 2.6061153
+ wtvoff = -3.3676979e-10
+ eta0 = 0.16744607
+ etab = -0.23671111
+ cjd = 0.001421376
+ cit = 0.00047888384
+ cjs = 0.001421376
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 1.38228675e-8
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ ijthsrev = 0.01
+ ku0we = -0.0007
+ beta0 = 13.32
+ capmod = 2
+ leta0 = -4.8e-10
+ la0 = -4.2186937e-8
+ poxedge = 1
+ wku0we = 1.5e-11
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0.00092821144
+ kt1 = -0.23884145
+ kt2 = -0.071460529
+ lk2 = 4.648829499999999e-9
+ llc = -1.18e-13
+ lln = 0.7
+ lu0 = -1.8531509e-10
+ mjd = 0.335
+ ppclm = 1.4344283e-14
+ mjs = 0.335
+ lua = -2.3141614e-17
+ lub = -3.0092793e-26
+ luc = -1.1168748e-18
+ lud = 0
+ lwc = 0
+ mobmod = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = -1.7418058e-15
+ nsd = 1e+20
+ binunit = 2
+ pbd = 0.75
+ pat = -2.5956322e-9
+ pbs = 0.75
+ pk2 = -2.0925962e-16
+ dlcig = 2.5e-9
+ pu0 = 6.8306111e-19
+ bgidl = 1834800000.0
+ prt = 0
+ pua = -2.4112447e-23
+ pub = 3.4375734e-32
+ puc = -1.1236355e-25
+ pud = 0
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 2.2048659e-9
+ ub1 = -2.7884819e-18
+ ppdiblc2 = 4.3354985e-16
+ uc1 = 8.0779763e-11
+ tpb = 0.0016
+ wa0 = -4.9541389e-7
+ ute = -1
+ wat = 0.012301575
+ web = 6628.3
+ wec = -16935.0
+ wk2 = -3.1036812e-9
+ wlc = 0
+ wln = 1
+ wu0 = -6.065551e-11
+ xgl = -8.2e-9
+ xgw = 0
+ wua = 3.8537331e-17
+ wub = -2.8668372e-25
+ wuc = -2.6715958e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ wtvfbsdoff = 0
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ bigsd = 0.0003327
+ ltvfbsdoff = 0
+ pkvth0we = 0.0
+ wvoff = 5.8569161e-9
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ wvsat = -0.0057246059
+ vfbsdoff = 0.01
+ keta = -0.13181891
+ wvth0 = 2.7825094999999996e-9
+ waigc = 1.3273811e-11
+ lags = 2.4408277e-8
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 8.8475659e-11
+ a0 = 1.505864
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ kt1l = 0
+ ptvfbsdoff = 0
+ at = 70634.069
+ paramchk = 1
+ cf = 8.17e-11
+ lketa = 1.156253e-9
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.013605325
+ k3 = -2.5823
+ em = 20000000.0
+ ll = -1.18e-13
+ lw = 0
+ u0 = 0.0093288547
+ w0 = 0
+ xpart = 1
+ ua = -3.2299413e-10
+ ub = 1.7243624e-18
+ uc = 2.4608838e-11
+ ud = 0
+ njtsswg = 6.489
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 3.4e-9
+ lint = 9.7879675e-9
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ lkt1 = -5.2521669e-9
+ lkt2 = -4.3239941e-10
+ egidl = 0.001
+ lmax = 2.1577e-7
+ lmin = 9e-8
+ toxref = 3e-9
+ ckappad = 0.6
+ ckappas = 0.6
+ lpe0 = 6.44e-8
+ pdiblc1 = 0
+ pdiblc2 = 0.017260131
+ lpeb = 0
+ pdiblcb = 0
+ ijthdfwd = 0.01
+ minv = -0.33
+ lua1 = -1.4410376e-16
+ lub1 = 1.6275827e-25
+ luc1 = 6.550381e-18
+ ndep = 1e+18
+ lwlc = 0
+ moin = 5.5538
+ bigbacc = 0.0054401
+ nigc = 2.291
+ ltvoff = -6.4284173e-11
+ ijthdrev = 0.01
+ pvfbsdoff = 0
+ lpdiblc2 = -1.5457732e-9
+ kvth0we = -0.00022
+ pvoff = -7.636562e-16
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ cdscb = 0
+ cdscd = 0
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ pvsat = -8.5382639e-10
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ wk2we = 0.0
+ )

.model pch_fs_14 pmos (
+ level = 54
+ cjd = 0.001421376
+ poxedge = 1
+ cit = -0.00080588346
+ wua1 = -1.4703955e-15
+ cjs = 0.001421376
+ clc = 1e-7
+ cle = 0.6
+ wub1 = 2.631826e-24
+ bvd = 8.2
+ wuc1 = 2.762344e-16
+ bvs = 8.2
+ igcmod = 1
+ dlc = 4.0349e-9
+ k3b = 2.1176
+ tvoff = 0.0011122833
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ bigc = 0.0012521
+ wwlc = 0
+ xjbvd = 1
+ binunit = 2
+ xjbvs = 1
+ lk2we = 0.0
+ pkvth0we = 0.0
+ la0 = -2.3326483e-7
+ jsd = 1.5e-7
+ cdsc = 0
+ jss = 1.5e-7
+ lat = -0.0059102639
+ kt1 = -0.2764195
+ kt2 = -0.075556865
+ lk2 = 4.2009156999999995e-9
+ llc = 0
+ cgbo = 0
+ lln = 1
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ lu0 = 2.0564492e-10
+ xtid = 3
+ xtis = 3
+ mjd = 0.335
+ mjs = 0.335
+ lua = 5.4621428e-17
+ lub = 1.4388057e-26
+ luc = 1.0238844e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ cgsl = 3.0105e-11
+ njs = 1.02
+ cgso = 2.6482e-11
+ pa0 = 5.4920056e-14
+ cigc = 0.15259
+ ku0we = -0.0007
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 1.0391973e-9
+ pbs = 0.75
+ pk2 = 6.854543e-16
+ beta0 = 13.32
+ vfbsdoff = 0.01
+ pu0 = -1.2707891e-16
+ leta0 = -1.1282603899999999e-9
+ prt = 0
+ pua = -5.2218942e-24
+ pub = -3.6833051e-32
+ puc = -9.869134e-24
+ pud = 0
+ letab = 2.0996791e-8
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 8.9078668e-10
+ ub1 = -1.404024e-18
+ uc1 = 4.4088848e-11
+ ppclm = 7.4853015e-14
+ tpb = 0.0016
+ wa0 = -1.0981997e-6
+ ute = -1
+ wat = -0.026366825
+ web = 6628.3
+ wec = -16935.0
+ wk2 = -1.2621914e-8
+ wlc = 0
+ dlcig = 2.5e-9
+ permod = 1
+ wln = 1
+ wu0 = 1.2985144e-9
+ xgl = -8.2e-9
+ xgw = 0
+ bgidl = 1834800000.0
+ wua = -1.62426e-16
+ wub = 4.7085654e-25
+ wuc = 7.7079472e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ paramchk = 1
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ k2we = 5e-5
+ voffcv = -0.125
+ wpemod = 1
+ dsub = 0.5
+ dtox = 3.91e-10
+ ijthdfwd = 0.01
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ bigsd = 0.0003327
+ eta0 = 0.17434246
+ etab = -0.46008122
+ njtsswg = 6.489
+ wvoff = -4.5993296e-9
+ ijthdrev = 0.01
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ wvsat = -0.039767366
+ wvth0 = -1.8578701e-8
+ lpdiblc2 = 0
+ ckappad = 0.6
+ tpbswg = 0.001
+ ckappas = 0.6
+ waigc = -2.1370578e-11
+ pdiblc1 = 0
+ pdiblc2 = 0.00081573526
+ pdiblcb = 0
+ lketa = 9.0137227e-9
+ xpart = 1
+ ptvoff = 1.200911e-16
+ waigsd = 1.9051377e-12
+ bigbacc = 0.0054401
+ egidl = 0.001
+ lkvth0we = 3e-12
+ diomod = 1
+ kvth0we = -0.00022
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.9113600000000002e-10
+ pku0we = 0.0
+ cjswgs = 1.9113600000000002e-10
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ acnqsmod = 0
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ rbodymod = 0
+ mjswgd = 0.95
+ mjswgs = 0.95
+ pvfbsdoff = 0
+ tcjswg = 0.00128
+ keta = -0.21540901
+ pvoff = 2.1923089e-16
+ cdscb = 0
+ cdscd = 0
+ lags = -3.1969346e-8
+ pvsat = 2.3461931e-9
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ wk2we = 0.0
+ pvth0 = 1.1602649e-15
+ lcit = 2.0924378e-10
+ drout = 0.56
+ kt1l = 0
+ paigc = 2.5179991e-18
+ voffl = 0
+ wpdiblc2 = 1.6594883e-9
+ lint = 0
+ lkt1 = -1.7198309e-9
+ lkt2 = -4.7343777e-11
+ weta0 = 4.2195709999999996e-8
+ nfactor = 1
+ lmax = 9e-8
+ wetab = 1.3144359e-7
+ fprout = 200
+ lmin = 5.4e-8
+ lpclm = -1.0675035e-7
+ xrcrg1 = 12
+ xrcrg2 = 1
+ lpe0 = 6.44e-8
+ lpeb = 0
+ cgidl = 1
+ minv = -0.33
+ lua1 = -2.0580314e-17
+ lub1 = 3.261922e-26
+ luc1 = 9.999327e-18
+ wtvoff = -1.8141864e-9
+ ndep = 1e+18
+ lwlc = 0
+ moin = 5.5538
+ wkvth0we = 0.0
+ nigbacc = 10
+ pbswd = 0.9
+ nigc = 2.291
+ pbsws = 0.9
+ capmod = 2
+ trnqsmod = 0
+ wku0we = 1.5e-11
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ mobmod = 0
+ pdits = 0
+ nigbinv = 2.171
+ cigsd = 0.013281
+ pags = 2.8964227e-14
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ wtvfbsdoff = 0
+ ntox = 1.0
+ pcit = -7.036540399999999e-17
+ pclm = 2.5596902
+ rgatemod = 0
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ tnjtsswg = 1
+ ltvfbsdoff = 0
+ phin = 0.15
+ pkt1 = 3.7820041e-17
+ pkt2 = 1.7971063e-15
+ fnoimod = 1
+ tnoia = 0
+ eigbinv = 1.1
+ peta0 = -4.2117702e-15
+ petab = -6.6743123e-15
+ wketa = 8.0928346e-8
+ tpbsw = 0.0025
+ rbdb = 50
+ pua1 = 1.1954606e-22
+ prwb = 0
+ pub1 = -2.033661e-31
+ prwg = 0
+ puc1 = -2.1449333e-23
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ cjswd = 5.3856e-11
+ pvag = 2.1
+ cjsws = 5.3856e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ rdsw = 200
+ ptvfbsdoff = 0
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ cigbacc = 0.245
+ tnoimod = 0
+ rshg = 14.1
+ scref = 1e-6
+ pigcd = 2.572
+ cigbinv = 0.006
+ aigsd = 0.0063634291
+ lvoff = -2.6816163e-9
+ toxref = 3e-9
+ lvsat = -0.0059751154
+ lvth0 = -1.7902539e-9
+ version = 4.5
+ ijthsfwd = 0.01
+ delta = 0.018814
+ tvfbsdoff = 0.1
+ tempmod = 0
+ laigc = -1.5433256e-11
+ tnom = 25
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ rnoia = 0
+ rnoib = 0
+ aigbacc = 0.012071
+ ltvoff = 1.2625293e-11
+ pketa = -4.6938441e-15
+ a0 = 3.5386076
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ ngate = 1.7e+20
+ at = 143383.81
+ cf = 8.17e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.0088402851
+ k3 = -2.5823
+ ijthsrev = 0.01
+ em = 20000000.0
+ ngcon = 1
+ ll = 0
+ lw = 0
+ u0 = 0.0051697056
+ wpclm = -1.0128863e-6
+ w0 = 0
+ ua = -1.1502605e-9
+ ub = 1.2511619e-18
+ uc = -9.619668e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 3.4e-9
+ gbmin = 1e-12
+ wags = 9.0067526e-7
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ aigbinv = 0.009974
+ wcit = 7.2293275e-10
+ lku0we = 1.8e-11
+ wvfbsdoff = 0
+ epsrox = 3.9
+ lvfbsdoff = 0
+ voff = -0.11844975
+ acde = 0.5
+ vsat = 190294.39
+ ppdiblc2 = 0
+ rdsmod = 0
+ wint = 0
+ vth0 = -0.35947984
+ igbmod = 1
+ wkt1 = -4.5227706e-9
+ wkt2 = -2.9740529e-8
+ wmax = 9.0026e-6
+ aigc = 0.0067091511
+ wmin = 9.025999999999999e-7
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ pbswgd = 0.8
+ ags = 3.2058772
+ pbswgs = 0.8
+ )

.model pch_fs_15 pmos (
+ level = 54
+ keta = 0.054978601
+ fnoimod = 1
+ pdits = 0
+ eigbinv = 1.1
+ cigsd = 0.013281
+ permod = 1
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 3.46566e-10
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ kt1l = 0
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ lint = 0
+ lkt1 = -1.4088112e-8
+ lkt2 = 1.0752811e-9
+ lmax = 5.4e-8
+ lmin = 4.5e-8
+ voffcv = -0.125
+ wpemod = 1
+ tnoia = 0
+ lpe0 = 6.44e-8
+ lpeb = 0
+ ijthsfwd = 0.01
+ cigbacc = 0.245
+ peta0 = 5.9336569e-15
+ petab = -1.9628815e-15
+ minv = -0.33
+ lua1 = -1.9488641e-18
+ lub1 = 6.8003561e-26
+ wketa = -5.4843946e-8
+ luc1 = -2.115524e-18
+ tpbsw = 0.0025
+ ndep = 1e+18
+ tnoimod = 0
+ cjswd = 5.3856e-11
+ lwlc = 0
+ cjsws = 5.3856e-11
+ moin = 5.5538
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ nigc = 2.291
+ cigbinv = 0.006
+ ijthsrev = 0.01
+ tpbswg = 0.001
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ version = 4.5
+ tempmod = 0
+ ntox = 1.0
+ pcit = -7.1417065e-17
+ pclm = 1.3082183
+ scref = 1e-6
+ ptvoff = 9.8606268e-17
+ ppdiblc2 = 0
+ pigcd = 2.572
+ aigsd = 0.0063634291
+ waigsd = 1.9051377e-12
+ aigbacc = 0.012071
+ phin = 0.15
+ lvoff = -4.1725981e-9
+ diomod = 1
+ pkt1 = 1.3908108999999999e-14
+ pkt2 = -4.0388508e-15
+ lvsat = -0.00018689407999999998
+ lvth0 = -2.2826855e-9
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.9113600000000002e-10
+ pku0we = 0.0
+ cjswgs = 1.9113600000000002e-10
+ tvfbsdoff = 0.1
+ delta = 0.018814
+ aigbinv = 0.009974
+ laigc = -9.3796225e-12
+ rnoia = 0
+ rnoib = 0
+ rbdb = 50
+ pua1 = -1.9221227e-22
+ prwb = 0
+ pub1 = 2.2863324e-31
+ prwg = 0
+ puc1 = 2.3602641e-23
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ pkvth0we = 0.0
+ rbsb = 50
+ pvag = 2.1
+ mjswgd = 0.95
+ mjswgs = 0.95
+ rdsw = 200
+ pketa = 3.1809489e-15
+ ngate = 1.7e+20
+ ngcon = 1
+ tcjswg = 0.00128
+ wpclm = 1.8421624e-6
+ vfbsdoff = 0.01
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ poxedge = 1
+ paramchk = 1
+ rshg = 14.1
+ binunit = 2
+ ags = 2.6546816
+ cjd = 0.001421376
+ cit = -0.0031735079
+ cjs = 0.001421376
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 4.0349e-9
+ fprout = 200
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ ijthdfwd = 0.01
+ la0 = -1.5436392e-7
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0.0049643403
+ kt1 = -0.063173267
+ kt2 = -0.094912467
+ lk2 = 4.598719299999999e-9
+ llc = 0
+ tvoff = 0.0053332949
+ lln = 1
+ lu0 = -6.2656189e-11
+ wtvoff = -1.4437583e-9
+ tnom = 25
+ mjd = 0.335
+ mjs = 0.335
+ lua = -3.3837758e-17
+ lub = -3.4072549e-26
+ luc = -2.4014309e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = -3.174587e-14
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ xjbvd = 1
+ xjbvs = 1
+ nsd = 1e+20
+ pbd = 0.75
+ pat = -5.2399134e-10
+ lk2we = 0.0
+ pbs = 0.75
+ pk2 = 5.1035691e-16
+ pu0 = -9.701894e-17
+ prt = 0
+ pua = -1.0296702e-22
+ pub = 1.290002e-31
+ puc = 2.16225e-23
+ pud = 0
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ rsh = 15.2
+ wtvfbsdoff = 0
+ tcj = 0.000832
+ ua1 = 5.6955479e-10
+ ub1 = -2.0140988e-18
+ uc1 = 2.5296559e-10
+ ijthdrev = 0.01
+ capmod = 2
+ tpb = 0.0016
+ wa0 = 3.9604044e-7
+ ute = -1
+ wat = 0.00058470362
+ ku0we = -0.0007
+ web = 6628.3
+ wec = -16935.0
+ wk2 = -9.6029938e-9
+ wku0we = 1.5e-11
+ wlc = 0
+ beta0 = 13.32
+ wln = 1
+ wu0 = 7.8023907e-10
+ xgl = -8.2e-9
+ xgw = 0
+ lpdiblc2 = 0
+ wua = 1.5228349e-15
+ wub = -2.3883374e-24
+ leta0 = -2.8597369e-9
+ wuc = -4.6587973e-16
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ letab = 1.0403109e-8
+ ltvfbsdoff = 0
+ mobmod = 0
+ wags = 1.4000585e-6
+ ppclm = -9.0739811e-14
+ wcit = 7.4106483e-10
+ voff = -0.092743162
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ acde = 0.5
+ vsat = 90497.467
+ wint = 0
+ vth0 = -0.35098964000000005
+ wkt1 = -2.4366569e-7
+ wkt2 = 7.087942e-8
+ wmax = 9.0026e-6
+ aigc = 0.0066047781
+ wmin = 9.025999999999999e-7
+ njtsswg = 6.489
+ dmcgt = 0
+ lkvth0we = 3e-12
+ tcjsw = 9.34e-5
+ ptvfbsdoff = 0
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ wua1 = 3.9047481e-15
+ wub1 = -4.8164385e-24
+ wuc1 = -5.0052376e-16
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.00081573526
+ pdiblcb = 0
+ bigc = 0.0012521
+ acnqsmod = 0
+ wwlc = 0
+ bigsd = 0.0003327
+ cdsc = 0
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ wvoff = 1.0199556e-9
+ rbodymod = 0
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigc = 0.15259
+ wvsat = -0.0078232946
+ bigbacc = 0.0054401
+ wvth0 = 4.6032398999999996e-8
+ waigc = 1.173226e-10
+ kvth0we = -0.00022
+ lintnoi = -5e-9
+ lketa = -6.6687589e-9
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ xpart = 1
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ wpdiblc2 = 1.6594883e-9
+ toxref = 3e-9
+ egidl = 0.001
+ k2we = 5e-5
+ dsub = 0.5
+ dtox = 3.91e-10
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ eta0 = 0.2041955
+ etab = -0.27743155
+ ltvoff = -2.3219338e-10
+ wkvth0we = 0.0
+ pvfbsdoff = 0
+ trnqsmod = 0
+ nfactor = 1
+ pvoff = -1.0668764999999999e-16
+ lku0we = 1.8e-11
+ cdscb = 0
+ cdscd = 0
+ epsrox = 3.9
+ pvsat = 4.9343693e-10
+ wk2we = 0.0
+ pvth0 = -2.5871789e-15
+ drout = 0.56
+ paigc = -5.5262052e-18
+ rdsmod = 0
+ igbmod = 1
+ rgatemod = 0
+ voffl = 0
+ tnjtsswg = 1
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ nigbacc = 10
+ weta0 = -1.3272544999999998e-7
+ wetab = 5.0212024e-8
+ pbswgd = 0.8
+ pbswgs = 0.8
+ lpclm = -3.4164983e-8
+ a0 = 2.1782471
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = -44109.368
+ cf = 8.17e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.015698968
+ k3 = -2.5823
+ em = 20000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.0097955868
+ w0 = 0
+ igcmod = 1
+ ua = 3.7489785e-10
+ ub = 2.0866896e-18
+ uc = 4.9437493e-10
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 3.4e-9
+ cgidl = 1
+ nigbinv = 2.171
+ pbswd = 0.9
+ pbsws = 0.9
+ )

.model pch_fs_16 pmos (
+ level = 54
+ wpdiblc2 = 1.6594883e-9
+ voffcv = -0.125
+ wpemod = 1
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ bigbacc = 0.0054401
+ tnom = 25
+ kvth0we = -0.00022
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ bigsd = 0.0003327
+ lintnoi = -5e-9
+ wkvth0we = 0.0
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ wvoff = -9.7608128e-9
+ trnqsmod = 0
+ wvsat = -0.0020201595
+ tpbswg = 0.001
+ wvth0 = 5.473123299999998e-9
+ wags = 3.1454838e-6
+ waigc = -1.1150212e-11
+ wcit = -4.2593599e-9
+ voff = -0.099237323
+ acde = 0.5
+ lketa = 8.2510741e-9
+ ptvoff = -1.3565734e-16
+ xpart = 1
+ waigsd = 2.0479558e-12
+ vsat = 122744.64
+ wint = 0
+ rgatemod = 0
+ vth0 = -0.39323313000000004
+ wkt1 = 3.1251908e-7
+ wkt2 = -1.0928272e-8
+ tnjtsswg = 1
+ wmax = 9.0026e-6
+ aigc = 0.0065575398
+ wmin = 9.025999999999999e-7
+ diomod = 1
+ egidl = 0.001
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.9113600000000002e-10
+ pku0we = 0.0
+ cjswgs = 1.9113600000000002e-10
+ nfactor = 1
+ wua1 = -3.8771176e-15
+ wub1 = 4.4904637e-24
+ wuc1 = 9.3089203e-17
+ bigc = 0.0012521
+ wwlc = 0
+ mjswgd = 0.95
+ mjswgs = 0.95
+ pvfbsdoff = 0
+ cdsc = 0
+ tcjswg = 0.00128
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigc = 0.15259
+ nigbacc = 10
+ pvoff = 4.2156999999999997e-16
+ cdscb = 0
+ cdscd = 0
+ pvsat = 2.0908331e-10
+ wk2we = 0.0
+ pvth0 = -5.997744e-16
+ drout = 0.56
+ paigc = 7.6896258e-19
+ nigbinv = 2.171
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ voffl = 0
+ dmdg = 0
+ fprout = 200
+ weta0 = 4.7064045e-9
+ xrcrg1 = 12
+ xrcrg2 = 1
+ wetab = 3.974597e-8
+ wtvfbsdoff = 0
+ lpclm = -2.1829165e-8
+ k2we = 5e-5
+ dsub = 0.5
+ dtox = 3.91e-10
+ ijthsfwd = 0.01
+ wtvoff = 3.3371317e-9
+ cgidl = 1
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ fnoimod = 1
+ ltvfbsdoff = 0
+ eigbinv = 1.1
+ eta0 = 0.11033512
+ etab = -0.14869011
+ capmod = 2
+ pbswd = 0.9
+ pbsws = 0.9
+ ijthsrev = 0.01
+ wku0we = 1.5e-11
+ mobmod = 0
+ pdits = 0
+ cigsd = 0.013281
+ ptvfbsdoff = 0
+ cigbacc = 0.245
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ ppdiblc2 = 0
+ tnoimod = 0
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ laigsd = 7.7486946e-16
+ cigbinv = 0.006
+ tnoia = 0
+ peta0 = -8.0050381e-16
+ petab = -1.4500449e-15
+ wketa = 4.9202854e-8
+ version = 4.5
+ tpbsw = 0.0025
+ tempmod = 0
+ cjswd = 5.3856e-11
+ pkvth0we = 0.0
+ cjsws = 5.3856e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ agidl = 3.2166e-9
+ aigbacc = 0.012071
+ vfbsdoff = 0.01
+ keta = -0.24950779
+ lags = 9.4399385e-8
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 2.1550138e-10
+ aigbinv = 0.009974
+ kt1l = 0
+ paramchk = 1
+ scref = 1e-6
+ pigcd = 2.572
+ aigsd = 0.0063634133
+ toxref = 3e-9
+ lint = 0
+ lvoff = -3.8543842e-9
+ lkt1 = -5.9161514e-10
+ lkt2 = 4.9336152e-10
+ lmax = 4.5e-8
+ lmin = 3.6e-8
+ lpe0 = 6.44e-8
+ lvsat = -0.0017670054
+ lpeb = 0
+ tvfbsdoff = 0.1
+ lvth0 = -2.12754306e-10
+ ijthdfwd = 0.01
+ delta = 0.018814
+ laigc = -7.0649434e-12
+ minv = -0.33
+ lua1 = -6.8231177e-17
+ lub1 = 7.1697841e-26
+ luc1 = 2.786749e-18
+ poxedge = 1
+ rnoia = 0
+ rnoib = 0
+ ndep = 1e+18
+ ltvoff = -9.8738127e-12
+ lwlc = 0
+ moin = 5.5538
+ binunit = 2
+ pketa = -1.9173443e-15
+ ngate = 1.7e+20
+ nigc = 2.291
+ ijthdrev = 0.01
+ ngcon = 1
+ wpclm = -3.2091624e-7
+ lpdiblc2 = 0
+ gbmin = 1e-12
+ lku0we = 1.8e-11
+ noff = 2.2684
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ epsrox = 3.9
+ ags = 0.72816353
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ cjd = 0.001421376
+ cit = -0.00049871975
+ cjs = 0.001421376
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ pags = -8.5525843e-14
+ dlc = 4.0349e-9
+ k3b = 2.1176
+ rdsmod = 0
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ ntox = 1.0
+ pcit = 1.7360375e-16
+ pclm = 1.0564669
+ igbmod = 1
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ la0 = -3.7737017e-8
+ jsd = 1.5e-7
+ phin = 0.15
+ jss = 1.5e-7
+ lat = -0.0012751021999999998
+ jtsswgd = 1.75e-7
+ kt1 = -0.33861198
+ kt2 = -0.083036557
+ lk2 = 4.3783258e-9
+ jtsswgs = 1.75e-7
+ llc = 0
+ lln = 1
+ pbswgd = 0.8
+ pbswgs = 0.8
+ lu0 = 1.5237989e-10
+ mjd = 0.335
+ mjs = 0.335
+ lua = 2.9640356e-17
+ lub = 1.5163389e-26
+ luc = -2.5002144e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ lkvth0we = 3e-12
+ njd = 1.02
+ njs = 1.02
+ pa0 = -1.5136929e-14
+ pkt1 = -1.3344944000000001e-14
+ pkt2 = -3.0273858e-17
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 2.5964497e-9
+ pbs = 0.75
+ pk2 = 4.883387e-16
+ igcmod = 1
+ pu0 = -4.5849539e-17
+ prt = 0
+ pua = 8.5912273e-23
+ pub = -1.727672e-31
+ puc = 8.2880171e-25
+ pud = 0
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 1.9222551e-9
+ ub1 = -2.0894923e-18
+ uc1 = 1.529192e-10
+ tvoff = 0.00079616085
+ tpb = 0.0016
+ wa0 = 5.7082474e-8
+ acnqsmod = 0
+ xjbvd = 1
+ ute = -1
+ wat = -0.063097766
+ xjbvs = 1
+ web = 6628.3
+ wec = -16935.0
+ rbdb = 50
+ wk2 = -9.1536426e-9
+ pua1 = 1.8909915e-22
+ prwb = 0
+ lk2we = 0.0
+ pub1 = -2.2740497e-31
+ prwg = 0
+ puc1 = -5.4843946e-24
+ wlc = 0
+ wln = 1
+ wu0 = -2.6403442e-10
+ xgl = -8.2e-9
+ rbpb = 50
+ rbpd = 50
+ xgw = 0
+ rbps = 50
+ rbsb = 50
+ wua = -2.3318447e-15
+ pvag = 2.1
+ wub = 3.770181e-24
+ wuc = -4.1518546e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ rdsw = 200
+ rbodymod = 0
+ paigsd = -6.9980875e-21
+ ku0we = -0.0007
+ beta0 = 13.32
+ njtsswg = 6.489
+ leta0 = 1.7394218e-9
+ letab = 4.094779e-9
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ ppclm = 1.5251044e-14
+ permod = 1
+ a0 = -0.20189383
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ ckappad = 0.6
+ at = 83226.192
+ cf = 8.17e-11
+ ckappas = 0.6
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.01120114
+ k3 = -2.5823
+ em = 20000000.0
+ dlcig = 2.5e-9
+ pdiblc1 = 0
+ pdiblc2 = 0.00081573526
+ ll = 0
+ lw = 0
+ bgidl = 1834800000.0
+ u0 = 0.0054070954
+ w0 = 0
+ pdiblcb = 0
+ ua = -9.2057386e-10
+ ub = 1.0818745e-18
+ uc = 5.5311765e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 3.4e-9
+ rshg = 14.1
+ )

.model pch_fs_17 pmos (
+ level = 54
+ tpbsw = 0.0025
+ aigbinv = 0.009974
+ eta0 = 0.191845
+ cjswd = 5.3856e-11
+ cjsws = 5.3856e-11
+ etab = -0.18516667
+ a0 = 2.6112
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ at = 72000
+ cf = 8.17e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.0045864754
+ k3 = -2.5823
+ em = 20000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.0097859667
+ w0 = 0
+ ua = 1.9119717e-10
+ ub = 1.0765761e-18
+ uc = -8.28048e-12
+ ud = 0
+ ijthdrev = 0.01
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 3.4e-9
+ tpbswg = 0.001
+ lpdiblc2 = 0
+ ptvoff = 0
+ waigsd = 1.9350626e-12
+ scref = 1e-6
+ poxedge = 1
+ pigcd = 2.572
+ aigsd = 0.0063633642
+ diomod = 1
+ binunit = 2
+ lvoff = 0
+ pditsd = 0
+ lkvth0we = 3e-12
+ pditsl = 0
+ cjswgd = 1.9113600000000002e-10
+ pku0we = 0.0
+ cjswgs = 1.9113600000000002e-10
+ tvfbsdoff = 0.1
+ lvsat = 8.000000000000001e-6
+ lvth0 = -2.4e-10
+ delta = 0.018814
+ acnqsmod = 0
+ rnoia = 0
+ rnoib = 0
+ mjswgd = 0.95
+ mjswgs = 0.95
+ tcjswg = 0.00128
+ ngate = 1.7e+20
+ rbodymod = 0
+ ags = 0.98525249
+ ngcon = 1
+ wpclm = -5.08417e-8
+ cjd = 0.001421376
+ cit = 5e-6
+ cjs = 0.001421376
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ dlc = 1.0572421799999999e-8
+ k3b = 2.1176
+ dwb = 0
+ keta = -0.016063969
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ gbmin = 1e-12
+ wvfbsdoff = 0
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ lvfbsdoff = 0
+ wtvfbsdoff = 0
+ la0 = 0
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0.00064
+ lcit = 1.6e-11
+ kt1 = -0.18299632
+ lk2 = 3.2000000000000003e-10
+ kt2 = -0.042133438
+ llc = 0
+ lln = 1
+ lu0 = -8e-13
+ mjd = 0.335
+ kt1l = 0
+ mjs = 0.335
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 0
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ ltvfbsdoff = 0
+ pk2 = 0
+ wpdiblc2 = -1.7580235e-10
+ fprout = 200
+ pu0 = 0
+ prt = 0
+ pud = 0
+ lint = 6.5375218e-9
+ xrcrg1 = 12
+ xrcrg2 = 1
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 1.45515e-9
+ ub1 = -1.5029257e-18
+ uc1 = -4.3667733e-11
+ lkt1 = -4.8e-10
+ lmax = 2.001e-5
+ tpb = 0.0016
+ wa0 = 2.308488e-7
+ lmin = 8.9991e-6
+ ute = -0.96728333
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 1.3953799e-9
+ njtsswg = 6.489
+ lpe0 = 6.44e-8
+ wlc = 0
+ wln = 1
+ wu0 = 2.7482e-12
+ xgl = -8.2e-9
+ lpeb = 0
+ xgw = 0
+ wua = -1.5682603e-16
+ wub = 3.5681818e-26
+ wuc = 4.8873989e-18
+ wud = 0
+ wtvoff = -7.2458121e-11
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ tvoff = 0.0025973351
+ minv = -0.33
+ xjbvd = 1
+ xjbvs = 1
+ ckappad = 0.6
+ ckappas = 0.6
+ lk2we = 0.0
+ ndep = 1e+18
+ pdiblc1 = 0
+ pdiblc2 = 0.0032290423
+ pdiblcb = 0
+ lwlc = 0
+ ptvfbsdoff = 0
+ capmod = 2
+ wkvth0we = 0.0
+ moin = 5.5538
+ wku0we = 1.5e-11
+ nigc = 2.291
+ trnqsmod = 0
+ mobmod = 0
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = -4.8e-10
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ bigbacc = 0.0054401
+ ppclm = 0
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ kvth0we = -0.00022
+ ntox = 1.0
+ pcit = -8.000000000000001e-19
+ pclm = 1.2411167
+ rgatemod = 0
+ lintnoi = -5e-9
+ tnjtsswg = 1
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ phin = 0.15
+ vtsswgs = 1.1
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ pkt1 = -4e-17
+ bigsd = 0.0003327
+ rbdb = 50
+ prwb = 0
+ prwg = 0
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ rdsw = 200
+ wvoff = 3.276885e-9
+ wvsat = -0.017628054
+ wvth0 = -1.1005744000000004e-9
+ waigc = -7.2361068e-12
+ nfactor = 1
+ lketa = 0
+ rshg = 14.1
+ xpart = 1
+ toxref = 3e-9
+ egidl = 0.001
+ nigbacc = 10
+ ijthsfwd = 0.01
+ tnom = 25
+ ltvoff = 0
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ pvfbsdoff = 0
+ nigbinv = 2.171
+ ijthsrev = 0.01
+ lku0we = 1.8e-11
+ pvoff = 2e-17
+ epsrox = 3.9
+ wags = -3.1938756e-8
+ cdscb = 0
+ cdscd = 0
+ pvsat = 0
+ wk2we = 0.0
+ rdsmod = 0
+ pvth0 = -1.2e-16
+ fnoimod = 1
+ drout = 0.56
+ voff = -0.10917042
+ igbmod = 1
+ acde = 0.5
+ eigbinv = 1.1
+ ppdiblc2 = 0
+ vsat = 129757.01
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ wint = 0
+ voffl = 0
+ vth0 = -0.40724647
+ wkt1 = 1.4804073e-9
+ wkt2 = -8.3218931e-9
+ pbswgd = 0.8
+ pbswgs = 0.8
+ wmax = 9.025999999999999e-7
+ aigc = 0.0068422292
+ wmin = 5.426e-7
+ weta0 = -2.454557e-8
+ wetab = 1.3741e-8
+ igcmod = 1
+ lpclm = 0
+ wua1 = -5.289391e-16
+ wub1 = 6.5622425e-25
+ wuc1 = 2.3227786e-17
+ cgidl = 1
+ bigc = 0.0012521
+ wute = -1.003093e-7
+ cigbacc = 0.245
+ wwlc = 0
+ pkvth0we = 0.0
+ cdsc = 0
+ tnoimod = 0
+ pbswd = 0.9
+ pbsws = 0.9
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigc = 0.15259
+ vfbsdoff = 0.01
+ cigbinv = 0.006
+ permod = 1
+ pdits = 0
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ paramchk = 1
+ version = 4.5
+ tempmod = 0
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ voffcv = -0.125
+ wpemod = 1
+ aigbacc = 0.012071
+ k2we = 5e-5
+ tnoia = 0
+ dsub = 0.5
+ dtox = 3.91e-10
+ ijthdfwd = 0.01
+ peta0 = -1.6e-17
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ wketa = -3.7023239e-9
+ )

.model pch_fs_18 pmos (
+ level = 54
+ waigc = -9.2878513e-12
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ nigbacc = 10
+ ptvoff = 6.0745993e-16
+ pags = -1.6587566e-14
+ waigsd = 1.93751e-12
+ lketa = -8.0782883e-8
+ ntox = 1.0
+ pcit = -8.000000000000001e-19
+ pclm = 1.2411167
+ xpart = 1
+ ppdiblc2 = 2.0750737e-15
+ diomod = 1
+ nigbinv = 2.171
+ phin = 0.15
+ egidl = 0.001
+ pditsd = 0
+ pditsl = 0
+ a0 = 2.6572474
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ cjswgd = 1.9113600000000002e-10
+ pku0we = 0.0
+ cjswgs = 1.9113600000000002e-10
+ at = 72000
+ cf = 8.17e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.0050849127
+ k3 = -2.5823
+ em = 20000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.0096657581
+ pkt1 = 7.4478862e-15
+ pkt2 = 7.624365e-15
+ w0 = 0
+ ua = 1.8022848e-10
+ ub = 1.0497212e-18
+ uc = -5.9216956e-12
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 3.4e-9
+ mjswgd = 0.95
+ mjswgs = 0.95
+ rbdb = 50
+ pua1 = 3.0135942e-22
+ prwb = 0
+ pub1 = -6.7644414e-31
+ prwg = 0
+ fnoimod = 1
+ puc1 = -4.7294542e-23
+ pvfbsdoff = 0
+ wtvfbsdoff = 0
+ tcjswg = 0.00128
+ pkvth0we = 0.0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ eigbinv = 1.1
+ pute = 3.5290383e-14
+ rdsw = 200
+ ltvfbsdoff = 0
+ vfbsdoff = 0.01
+ pvoff = 8.1887382e-16
+ cdscb = 0
+ cdscd = 0
+ pvsat = 0
+ wk2we = 0.0
+ pvth0 = -1.2864923999999999e-15
+ drout = 0.56
+ paramchk = 1
+ paigc = 1.8445184e-17
+ rshg = 14.1
+ cigbacc = 0.245
+ fprout = 200
+ voffl = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ tnoimod = 0
+ ptvfbsdoff = 0
+ weta0 = -2.454557e-8
+ wetab = 1.3741e-8
+ lpclm = 0
+ wtvoff = -1.4002875e-10
+ cigbinv = 0.006
+ ijthdfwd = 0.01
+ cgidl = 1
+ tnom = 25
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ capmod = 2
+ version = 4.5
+ wku0we = 1.5e-11
+ tempmod = 0
+ pbswd = 0.9
+ pbsws = 0.9
+ ijthdrev = 0.01
+ mobmod = 0
+ lpdiblc2 = 3.0626629e-9
+ aigbacc = 0.012071
+ wags = -3.0093643e-8
+ pdits = 0
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ voff = -0.10728654
+ acde = 0.5
+ vsat = 129757.01
+ aigbinv = 0.009974
+ wint = 0
+ vth0 = -0.40617796
+ laigsd = 5.7445099e-14
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ wkt1 = 6.4749443e-10
+ wkt2 = -9.1699871e-9
+ wmax = 9.025999999999999e-7
+ aigc = 0.0068507406
+ wmin = 5.426e-7
+ lkvth0we = 3e-12
+ tnoia = 0
+ peta0 = -1.6e-17
+ wua1 = -5.6246072e-16
+ wub1 = 7.3146831e-25
+ wuc1 = 2.8488581e-17
+ wketa = -8.2059163e-9
+ bigc = 0.0012521
+ wute = -1.0423482e-7
+ acnqsmod = 0
+ tpbsw = 0.0025
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ wwlc = 0
+ cjswd = 5.3856e-11
+ cjsws = 5.3856e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ poxedge = 1
+ cdsc = 0
+ rbodymod = 0
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigc = 0.15259
+ binunit = 2
+ toxref = 3e-9
+ scref = 1e-6
+ pigcd = 2.572
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ wpdiblc2 = -4.0662257e-10
+ aigsd = 0.0063633578
+ dmdg = 0
+ lvoff = -1.6936099e-8
+ tvfbsdoff = 0.1
+ k2we = 5e-5
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ lvsat = 8.000000000000001e-6
+ lvth0 = -9.845867799999999e-9
+ dsub = 0.5
+ dtox = 3.91e-10
+ delta = 0.018814
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ laigc = -7.651731e-11
+ ltvoff = -1.5996918e-9
+ ags = 0.95300429
+ rnoia = 0
+ rnoib = 0
+ cjd = 0.001421376
+ cit = 5e-6
+ cjs = 0.001421376
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 1.0572421799999999e-8
+ k3b = 2.1176
+ eta0 = 0.191845
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ etab = -0.18516667
+ dwj = 0
+ wkvth0we = 0.0
+ pketa = 4.0487295e-14
+ ngate = 1.7e+20
+ ngcon = 1
+ wpclm = -5.08417e-8
+ trnqsmod = 0
+ la0 = -4.1396638e-7
+ lku0we = 1.8e-11
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0.00064
+ kt1 = -0.17852273
+ kt2 = -0.039741464
+ lk2 = 4.8009517e-9
+ llc = 0
+ lln = 1
+ epsrox = 3.9
+ lu0 = 1.0798753e-9
+ mjd = 0.335
+ wvfbsdoff = 0
+ mjs = 0.335
+ lua = 9.8608496e-17
+ lub = 2.4142536e-25
+ luc = -2.1205472e-17
+ lud = 0
+ gbmin = 1e-12
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ lvfbsdoff = 0
+ njd = 1.02
+ njs = 1.02
+ pa0 = -1.9681175e-13
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ pk2 = -1.7465146e-15
+ njtsswg = 6.489
+ pu0 = -2.7146448e-18
+ rdsmod = 0
+ prt = 0
+ pua = -5.0852536e-23
+ pub = 3.3773548e-32
+ puc = 2.1258791e-23
+ pud = 0
+ igbmod = 1
+ xtsswgd = 0.32
+ rsh = 15.2
+ xtsswgs = 0.32
+ tcj = 0.000832
+ ua1 = 1.3709274e-9
+ ub1 = -1.4287011e-18
+ uc1 = -6.3574807e-11
+ tpb = 0.0016
+ wa0 = 2.527411e-7
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ ute = -0.97152091
+ ckappad = 0.6
+ ckappas = 0.6
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 1.5896529e-9
+ wlc = 0
+ rgatemod = 0
+ wln = 1
+ pdiblc1 = 0
+ pdiblc2 = 0.0028883679
+ wu0 = 3.0501627e-12
+ xgl = -8.2e-9
+ xgw = 0
+ pbswgd = 0.8
+ pdiblcb = 0
+ wua = -1.5116947e-16
+ pbswgs = 0.8
+ wub = 3.1925028e-26
+ wuc = 2.5226836e-18
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ tnjtsswg = 1
+ igcmod = 1
+ tvoff = 0.0027752763
+ bigbacc = 0.0054401
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ kvth0we = -0.00022
+ paigsd = -2.2002196e-20
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ ku0we = -0.0007
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ beta0 = 13.32
+ leta0 = -4.8e-10
+ keta = -0.0070781088
+ permod = 1
+ ppclm = 0
+ lags = 2.8991134e-7
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ dlcig = 2.5e-9
+ lcit = 1.6e-11
+ bgidl = 1834800000.0
+ kt1l = 0
+ voffcv = -0.125
+ wpemod = 1
+ lint = 6.5375218e-9
+ lkt1 = -4.0697527e-8
+ lkt2 = -2.1503841e-8
+ dmcgt = 0
+ lmax = 8.9991e-6
+ tcjsw = 9.34e-5
+ lmin = 8.9908e-7
+ lpe0 = 6.44e-8
+ lpeb = 0
+ ijthsfwd = 0.01
+ minv = -0.33
+ lua1 = 7.5716104e-16
+ lub1 = -6.6727951e-25
+ luc1 = 1.7896459e-16
+ nfactor = 1
+ bigsd = 0.0003327
+ ndep = 1e+18
+ lute = 3.8095772e-8
+ lwlc = 0
+ moin = 5.5538
+ wvoff = 3.1880225e-9
+ tpbswg = 0.001
+ ijthsrev = 0.01
+ nigc = 2.291
+ wvsat = -0.017628054
+ wvth0 = -9.708200000000004e-10
+ noff = 2.2684
+ )

.model pch_fs_19 pmos (
+ level = 54
+ cjd = 0.001421376
+ cit = -8.7888889e-5
+ cjs = 0.001421376
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ lvsat = 8.000000000000001e-6
+ dlc = 1.0572421799999999e-8
+ k3b = 2.1176
+ lvth0 = -4.0657388e-10
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ ltvfbsdoff = 0
+ wua1 = -6.1430214e-16
+ wub1 = 1.1920544e-25
+ delta = 0.018814
+ wuc1 = -4.9561039e-17
+ laigc = -1.8208261e-11
+ mjswgd = 0.95
+ mjswgs = 0.95
+ njtsswg = 6.489
+ bigc = 0.0012521
+ wute = -1.2773023e-7
+ rnoia = 0
+ rnoib = 0
+ la0 = -9.6086602e-7
+ wwlc = 0
+ tcjswg = 0.00128
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0.00064
+ kt1 = -0.20738899
+ kt2 = -0.065812764
+ lk2 = 8.919589000000003e-11
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ llc = 0
+ lln = 1
+ lu0 = -1.5290408e-9
+ mjd = 0.335
+ mjs = 0.335
+ lua = -3.205013e-16
+ lub = -3.7552526e-26
+ luc = 5.1848161e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 2.9499704e-13
+ pketa = -2.8529622e-14
+ ckappad = 0.6
+ cdsc = 0
+ ckappas = 0.6
+ ngate = 1.7e+20
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ pk2 = 8.8602334e-16
+ pdiblc1 = 0
+ pdiblc2 = -8.9657994e-6
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ ngcon = 1
+ xtis = 3
+ pdiblcb = 0
+ pu0 = 4.0536683e-16
+ wpclm = -5.08417e-8
+ prt = 0
+ pua = 3.1718399e-23
+ pub = 9.4535502e-32
+ puc = -3.7711192e-23
+ pud = 0
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigc = 0.15259
+ rsh = 15.2
+ wvfbsdoff = 0
+ tcj = 0.000832
+ ua1 = 2.985915e-9
+ ub1 = -2.7037422e-18
+ uc1 = 1.5248758e-10
+ lvfbsdoff = 0
+ gbmin = 1e-12
+ tpb = 0.0016
+ wa0 = -2.9985305e-7
+ jswgd = 3.69e-13
+ ptvfbsdoff = 0
+ jswgs = 3.69e-13
+ ute = -0.85901741
+ web = 6628.3
+ wec = -16935.0
+ wk2 = -1.3682549e-9
+ a0 = 3.2717414
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ wlc = 0
+ wln = 1
+ wu0 = -4.5546835e-10
+ at = 72000
+ cf = 8.17e-11
+ xgl = -8.2e-9
+ ef = 1.15
+ k1 = 0.30425
+ k2 = 0.00020919492
+ xgw = 0
+ k3 = -2.5823
+ em = 20000000.0
+ wua = -2.439458e-16
+ wub = -3.6346832e-26
+ wuc = 6.8781092e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ ll = 0
+ lw = 0
+ u0 = 0.012597124
+ w0 = 0
+ ua = 6.5113837e-10
+ ub = 1.3631795e-18
+ uc = -8.8004429e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 3.4e-9
+ bigbacc = 0.0054401
+ fprout = 200
+ xrcrg1 = 12
+ xrcrg2 = 1
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ kvth0we = -0.00022
+ lintnoi = -5e-9
+ wtvoff = 9.9743807e-10
+ bigbinv = 0.00149
+ k2we = 5e-5
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ dsub = 0.5
+ dtox = 3.91e-10
+ ijthsfwd = 0.01
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ tvoff = 0.00044287651
+ capmod = 2
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ wku0we = 1.5e-11
+ eta0 = 0.191845
+ etab = -0.18516667
+ mobmod = 0
+ ijthsrev = 0.01
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = -4.8e-10
+ ppclm = 0
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ nfactor = 1
+ laigsd = -3.6354984e-15
+ ppdiblc2 = -2.7249029e-15
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ nigbacc = 10
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ bigsd = 0.0003327
+ pkvth0we = 0.0
+ wvoff = 1.2743983e-8
+ nigbinv = 2.171
+ wvsat = -0.017628054
+ vfbsdoff = 0.01
+ wvth0 = -2.8907114200000004e-9
+ keta = -0.13767457
+ waigc = 2.7297355e-11
+ lags = 8.1183869e-8
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 9.8671111e-11
+ toxref = 3e-9
+ paramchk = 1
+ lketa = 3.5447968e-8
+ kt1l = 0
+ xpart = 1
+ fnoimod = 1
+ eigbinv = 1.1
+ lint = 6.5375218e-9
+ egidl = 0.001
+ lkt1 = -1.5006561e-8
+ lkt2 = 1.6996159e-9
+ lmax = 8.9908e-7
+ lmin = 4.4908e-7
+ lpe0 = 6.44e-8
+ lpeb = 0
+ ijthdfwd = 0.01
+ ltvoff = 4.7614406e-10
+ minv = -0.33
+ lua1 = -6.8017788e-16
+ lub1 = 4.6750711e-25
+ luc1 = -1.3330934e-17
+ pvfbsdoff = 0
+ ndep = 1e+18
+ lute = -6.2032341e-8
+ lwlc = 0
+ moin = 5.5538
+ cigbacc = 0.245
+ ijthdrev = 0.01
+ nigc = 2.291
+ lku0we = 1.8e-11
+ epsrox = 3.9
+ tnoimod = 0
+ lpdiblc2 = 5.64129e-9
+ pvoff = -7.6859313e-15
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ rdsmod = 0
+ cdscb = 0
+ cdscd = 0
+ cigbinv = 0.006
+ igbmod = 1
+ pvsat = 0
+ wk2we = 0.0
+ pvth0 = 4.2221102000000002e-16
+ drout = 0.56
+ pags = 2.5130854e-13
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ paigc = -1.411565e-17
+ ntox = 1.0
+ pcit = -8.000000000000001e-19
+ pclm = 1.2411167
+ pbswgd = 0.8
+ pbswgs = 0.8
+ voffl = 0
+ version = 4.5
+ igcmod = 1
+ phin = 0.15
+ tempmod = 0
+ weta0 = -2.454557e-8
+ wetab = 1.3741e-8
+ lkvth0we = 3e-12
+ lpclm = 0
+ pkt1 = -4.6811548e-15
+ pkt2 = -3.0623252e-15
+ aigbacc = 0.012071
+ cgidl = 1
+ acnqsmod = 0
+ rbdb = 50
+ pua1 = 3.4749829e-22
+ prwb = 0
+ pub1 = -1.3153018e-31
+ prwg = 0
+ puc1 = 2.216962e-23
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ paigsd = 1.9849821e-21
+ rbsb = 50
+ pvag = 2.1
+ pute = 5.6201301e-14
+ rdsw = 200
+ rbodymod = 0
+ pbswd = 0.9
+ pbsws = 0.9
+ aigbinv = 0.009974
+ permod = 1
+ pdits = 0
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ rshg = 14.1
+ voffcv = -0.125
+ wpemod = 1
+ wpdiblc2 = 4.9866096e-9
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ poxedge = 1
+ tnoia = 0
+ binunit = 2
+ peta0 = -1.6e-17
+ wketa = 6.9341182e-8
+ tnom = 25
+ tpbsw = 0.0025
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ cjswd = 5.3856e-11
+ cjsws = 5.3856e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ wkvth0we = 0.0
+ agidl = 3.2166e-9
+ tpbswg = 0.001
+ trnqsmod = 0
+ wags = -3.311005e-7
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ ptvoff = -4.0488554e-16
+ waigsd = 1.9105581e-12
+ voff = -0.13228318
+ acde = 0.5
+ scref = 1e-6
+ diomod = 1
+ vsat = 129757.01
+ pigcd = 2.572
+ rgatemod = 0
+ wint = 0
+ aigsd = 0.0063634264
+ vth0 = -0.41678391000000004
+ tnjtsswg = 1
+ wkt1 = 1.4275631e-8
+ wkt2 = 2.8375299e-9
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.9113600000000002e-10
+ pku0we = 0.0
+ wmax = 9.025999999999999e-7
+ wtvfbsdoff = 0
+ cjswgs = 1.9113600000000002e-10
+ aigc = 0.0067852248
+ lvoff = 5.3109112e-9
+ wmin = 5.426e-7
+ ags = 1.1875295
+ tvfbsdoff = 0.1
+ )

.model pch_fs_20 pmos (
+ level = 54
+ cjd = 0.001421376
+ cit = -0.00041212495
+ cjs = 0.001421376
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ lvsat = 8.000000000000001e-6
+ dlc = 1.38228675e-8
+ k3b = 2.1176
+ lvth0 = 6.2654743e-9
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ ltvfbsdoff = 0
+ wua1 = 2.4012676e-16
+ wub1 = -6.2487918e-26
+ delta = 0.018814
+ wuc1 = -3.9943707e-17
+ laigc = -2.2400472e-11
+ mjswgd = 0.95
+ mjswgs = 0.95
+ njtsswg = 6.489
+ bigc = 0.0012521
+ rnoia = 0
+ rnoib = 0
+ la0 = -7.2511148e-8
+ wwlc = 0
+ tcjswg = 0.00128
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0.00064
+ kt1 = -0.20886849
+ kt2 = -0.049681978
+ lk2 = 1.5317426e-9
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ llc = -1.18e-13
+ lln = 0.7
+ lu0 = -4.8175715e-10
+ mjd = 0.335
+ mjs = 0.335
+ lua = -5.9775833e-17
+ lub = -8.2990392e-26
+ luc = -8.4878869e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = -2.0868237e-13
+ pketa = -1.8963071e-15
+ ckappad = 0.6
+ cdsc = 0
+ ckappas = 0.6
+ ngate = 1.7e+20
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ pk2 = -3.6576402e-16
+ pdiblc1 = 0
+ pdiblc2 = 0.01788848
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ ngcon = 1
+ xtis = 3
+ pdiblcb = 0
+ pu0 = -2.2283222e-17
+ wpclm = -5.08417e-8
+ prt = 0
+ pua = -3.7414239e-23
+ pub = 6.4271496e-32
+ puc = -3.5764571e-25
+ pud = 0
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigc = 0.15259
+ rsh = 15.2
+ wvfbsdoff = 0
+ tcj = 0.000832
+ ua1 = 1.3271195e-9
+ ub1 = -1.4620758e-18
+ uc1 = 1.6497662e-10
+ lvfbsdoff = 0
+ gbmin = 1e-12
+ tpb = 0.0016
+ wa0 = 8.4487289e-7
+ jswgd = 3.69e-13
+ ptvfbsdoff = 0
+ jswgs = 3.69e-13
+ ute = -1
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 1.4767164e-9
+ a0 = 1.2527531
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ wlc = 0
+ wln = 1
+ wu0 = 5.1646359e-10
+ at = 72000
+ cf = 8.17e-11
+ xgl = -8.2e-9
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.0030693202
+ xgw = 0
+ k3 = -2.5823
+ em = 20000000.0
+ wua = -8.6826164e-17
+ wub = 3.2435001e-26
+ wuc = -1.6113333e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ ll = -1.18e-13
+ lw = 0
+ u0 = 0.010216934
+ w0 = 0
+ ua = 5.8580479e-11
+ ub = 1.4664474e-18
+ uc = 4.9122952e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 3.4e-9
+ bigbacc = 0.0054401
+ fprout = 200
+ xrcrg1 = 12
+ xrcrg2 = 1
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ kvth0we = -0.00022
+ lintnoi = -5e-9
+ wtvoff = -3.604609e-11
+ bigbinv = 0.00149
+ k2we = 5e-5
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ dsub = 0.5
+ dtox = 3.91e-10
+ ijthsfwd = 0.01
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ tvoff = 0.0020688013
+ capmod = 2
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ wku0we = 1.5e-11
+ eta0 = 0.191845
+ etab = -0.18516667
+ mobmod = 0
+ ijthsrev = 0.01
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = -4.8e-10
+ ppclm = 0
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ nfactor = 1
+ ppdiblc2 = 1.0915468e-15
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ nigbacc = 10
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ bigsd = 0.0003327
+ pkvth0we = 0.0
+ wvoff = -5.0330429e-9
+ nigbinv = 2.171
+ wvsat = -0.017628054
+ vfbsdoff = 0.01
+ wvth0 = 2.3326608e-9
+ keta = -0.023696099
+ waigc = -1.2459534e-12
+ lags = 6.5053339e-7
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 2.4133498e-10
+ toxref = 3e-9
+ paramchk = 1
+ lketa = -1.4702559e-8
+ kt1l = 0
+ xpart = 1
+ fnoimod = 1
+ eigbinv = 1.1
+ lint = 9.7879675e-9
+ egidl = 0.001
+ lkt1 = -1.4355579e-8
+ lkt2 = -5.3979298e-9
+ lmax = 4.4908e-7
+ lmin = 2.1577e-7
+ lpe0 = 6.44e-8
+ lpeb = 0
+ ijthdfwd = 0.01
+ ltvoff = -2.3926284e-10
+ minv = -0.33
+ lua1 = 4.9692128e-17
+ lub1 = -7.8826099e-26
+ luc1 = -1.8826114e-17
+ pvfbsdoff = 0
+ ndep = 1e+18
+ lwlc = 0
+ moin = 5.5538
+ cigbacc = 0.245
+ ijthdrev = 0.01
+ nigc = 2.291
+ lku0we = 1.8e-11
+ epsrox = 3.9
+ tnoimod = 0
+ lpdiblc2 = -2.233586e-9
+ pvoff = 1.3596021e-16
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ rdsmod = 0
+ cdscb = 0
+ cdscd = 0
+ cigbinv = 0.006
+ igbmod = 1
+ pvsat = 0
+ wk2we = 0.0
+ pvth0 = -1.8760727e-15
+ drout = 0.56
+ pags = 1.3163813e-13
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ paigc = -1.5565945e-18
+ ntox = 1.0
+ pcit = -2.1300563999999998e-17
+ pclm = 1.2411167
+ pbswgd = 0.8
+ pbswgs = 0.8
+ voffl = 0
+ version = 4.5
+ igcmod = 1
+ phin = 0.15
+ tempmod = 0
+ weta0 = -2.454557e-8
+ wetab = 1.3741e-8
+ lkvth0we = 3e-12
+ lpclm = 0
+ pkt1 = 1.1173276e-15
+ pkt2 = 6.9635068e-17
+ aigbacc = 0.012071
+ cgidl = 1
+ acnqsmod = 0
+ rbdb = 50
+ pua1 = -2.8450432e-23
+ prwb = 0
+ pub1 = -5.1585101e-32
+ prwg = 0
+ puc1 = 1.7937993e-23
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ rdsw = 200
+ rbodymod = 0
+ pbswd = 0.9
+ pbsws = 0.9
+ aigbinv = 0.009974
+ permod = 1
+ pdits = 0
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ rshg = 14.1
+ voffcv = -0.125
+ wpemod = 1
+ wpdiblc2 = -3.6871397e-9
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ poxedge = 1
+ tnoia = 0
+ binunit = 2
+ peta0 = -1.6e-17
+ wketa = 8.8109206e-9
+ tnom = 25
+ tpbsw = 0.0025
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ cjswd = 5.3856e-11
+ cjsws = 5.3856e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ wkvth0we = 0.0
+ agidl = 3.2166e-9
+ tpbswg = 0.001
+ trnqsmod = 0
+ wags = -5.9122303e-8
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ ptvoff = 4.9847489e-17
+ wcit = 4.6592191e-11
+ waigsd = 1.9150694e-12
+ voff = -0.10909205
+ acde = 0.5
+ scref = 1e-6
+ diomod = 1
+ vsat = 129757.01
+ pigcd = 2.572
+ rgatemod = 0
+ wint = 0
+ aigsd = 0.0063634182
+ vth0 = -0.43194766
+ tnjtsswg = 1
+ wkt1 = 1.0972613e-9
+ wkt2 = -4.2805615e-9
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.9113600000000002e-10
+ pku0we = 0.0
+ wmax = 9.025999999999999e-7
+ wtvfbsdoff = 0
+ cjswgs = 1.9113600000000002e-10
+ aigc = 0.0067947526
+ lvoff = -4.893186e-9
+ wmin = 5.426e-7
+ ags = -0.10644665
+ tvfbsdoff = 0.1
+ )

.model pch_fs_21 pmos (
+ level = 54
+ rbodymod = 0
+ version = 4.5
+ tempmod = 0
+ keta = -0.074839654
+ pvoff = 2.997289e-16
+ cdscb = 0
+ cdscd = 0
+ lags = 2.5597727e-7
+ pvsat = 0
+ aigbacc = 0.012071
+ wk2we = 0.0
+ pvth0 = 3.0710494e-16
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ drout = 0.56
+ fprout = 200
+ lcit = 1.6312816e-10
+ kt1l = 0
+ paigc = 3.3660127e-18
+ xrcrg1 = 12
+ xrcrg2 = 1
+ voffl = 0
+ wpdiblc2 = 2.1803424e-9
+ lint = 9.7879675e-9
+ weta0 = -2.454557e-8
+ wtvoff = -4.3702924e-10
+ aigbinv = 0.009974
+ wetab = 1.3741e-8
+ lkt1 = -6.6443471e-9
+ lkt2 = -3.8990903e-9
+ lmax = 2.1577e-7
+ lpclm = 5.4900145e-8
+ lmin = 9e-8
+ lpe0 = 6.44e-8
+ lpeb = 0
+ cgidl = 1
+ minv = -0.33
+ capmod = 2
+ lua1 = -2.9544713e-16
+ lub1 = 3.7855773e-25
+ luc1 = 4.6029572e-17
+ wku0we = 1.5e-11
+ a0 = 0.98313605
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ ndep = 1e+18
+ at = 41320.114
+ cf = 8.17e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.016096302
+ k3 = -2.5823
+ em = 20000000.0
+ ll = -1.18e-13
+ lwlc = 0
+ lw = 0
+ u0 = 0.008766993
+ mobmod = 0
+ w0 = 0
+ wkvth0we = 0.0
+ ua = 2.7312462e-10
+ ub = 6.1180894e-19
+ uc = 6.0007215e-11
+ ud = 0
+ moin = 5.5538
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 3.4e-9
+ pbswd = 0.9
+ pbsws = 0.9
+ nigc = 2.291
+ trnqsmod = 0
+ poxedge = 1
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ binunit = 2
+ pdits = 0
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ pags = -1.3976359e-13
+ ntox = 1.0
+ pcit = -3.7185120000000004e-17
+ pclm = 0.98092641
+ rgatemod = 0
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ tnjtsswg = 1
+ phin = 0.15
+ pkt1 = 1.502035e-15
+ pkt2 = 2.2793112e-15
+ tnoia = 0
+ peta0 = -1.6e-17
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ wketa = -2.2984762e-8
+ tpbsw = 0.0025
+ rbdb = 50
+ pua1 = 7.9342593e-23
+ prwb = 0
+ pub1 = -9.194958e-32
+ prwg = 0
+ puc1 = -2.9723056e-23
+ cjswd = 5.3856e-11
+ cjsws = 5.3856e-11
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ mjswd = 0.01
+ rbsb = 50
+ pvag = 2.1
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ rdsw = 200
+ toxref = 3e-9
+ njtsswg = 6.489
+ ags = 1.7634876
+ scref = 1e-6
+ rshg = 14.1
+ cjd = 0.001421376
+ cit = -4.1476524e-5
+ cjs = 0.001421376
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ xtsswgd = 0.32
+ pigcd = 2.572
+ xtsswgs = 0.32
+ dlc = 1.38228675e-8
+ aigsd = 0.0063634182
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ tvfbsdoff = 0.1
+ ckappad = 0.6
+ ckappas = 0.6
+ lvoff = -2.4249846e-9
+ pdiblc1 = 0
+ pdiblc2 = 0.011594472
+ pdiblcb = 0
+ la0 = -1.5621959e-8
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0.007113456
+ lvsat = 8.000000000000001e-6
+ kt1 = -0.24541461
+ kt2 = -0.056785482
+ lk2 = 4.2804228e-9
+ llc = -1.18e-13
+ lvth0 = 3.7439767e-9
+ lln = 0.7
+ ltvoff = -2.3342435e-10
+ lu0 = -1.7581951e-10
+ mjd = 0.335
+ mjs = 0.335
+ lua = -1.0504465e-16
+ ijthsfwd = 0.01
+ lub = 9.7338322e-26
+ luc = -1.0784466e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ delta = 0.018814
+ pa0 = -2.5809676e-14
+ nsd = 1e+20
+ laigc = -2.5435198e-11
+ pbd = 0.75
+ pat = -8.1994638e-9
+ pbs = 0.75
+ pk2 = 1.2451684e-16
+ tnom = 25
+ pu0 = -7.9199366e-18
+ prt = 0
+ pua = 5.00917e-23
+ pub = -8.1076857e-32
+ puc = 8.6464743e-24
+ pud = 0
+ rnoia = 0
+ rnoib = 0
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 2.9628506e-9
+ ub1 = -3.6297717e-18
+ uc1 = -1.423963e-10
+ bigbacc = 0.0054401
+ tpb = 0.0016
+ wa0 = -2.1822352e-8
+ pketa = 4.8125819e-15
+ ute = -1
+ wat = 0.038860018
+ ngate = 1.7e+20
+ web = 6628.3
+ wec = -16935.0
+ lku0we = 1.8e-11
+ wk2 = -8.468563e-10
+ wlc = 0
+ wln = 1
+ ijthsrev = 0.01
+ wu0 = 4.4839114e-10
+ xgl = -8.2e-9
+ ngcon = 1
+ xgw = 0
+ epsrox = 3.9
+ wua = -5.0154626e-16
+ wub = 7.2128975e-25
+ wuc = -5.8786887e-17
+ wud = 0
+ wpclm = 1.8489068e-7
+ wwc = 0
+ kvth0we = -0.00022
+ wwl = 0
+ wwn = 1
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ gbmin = 1e-12
+ lintnoi = -5e-9
+ rdsmod = 0
+ jswgd = 3.69e-13
+ bigbinv = 0.00149
+ jswgs = 3.69e-13
+ wags = 1.2271418e-6
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ igbmod = 1
+ wcit = 1.2187445e-10
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ voff = -0.12078969
+ acde = 0.5
+ pbswgd = 0.8
+ pbswgs = 0.8
+ ppdiblc2 = -1.4649193e-16
+ vsat = 129757.01
+ wint = 0
+ vth0 = -0.41999743
+ igcmod = 1
+ wkt1 = -7.259963e-10
+ wkt2 = -1.475296e-8
+ wmax = 9.025999999999999e-7
+ aigc = 0.0068091352
+ wmin = 5.426e-7
+ wua1 = -2.7074066e-16
+ wub1 = 1.2881293e-25
+ wuc1 = 1.8593804e-16
+ tvoff = 0.0020411307
+ bigc = 0.0012521
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ wwlc = 0
+ pkvth0we = 0.0
+ nfactor = 1
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ permod = 1
+ ku0we = -0.0007
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigc = 0.15259
+ beta0 = 13.32
+ vfbsdoff = 0.01
+ leta0 = -4.8e-10
+ ppclm = -4.9739531e-14
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ nigbacc = 10
+ paramchk = 1
+ voffcv = -0.125
+ wpemod = 1
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ nigbinv = 2.171
+ k2we = 5e-5
+ dsub = 0.5
+ ijthdfwd = 0.01
+ dtox = 3.91e-10
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ bigsd = 0.0003327
+ eta0 = 0.191845
+ tpbswg = 0.001
+ etab = -0.18516667
+ wvoff = -5.8091978e-9
+ fnoimod = 1
+ ijthdrev = 0.01
+ eigbinv = 1.1
+ wvsat = -0.017628054
+ wvth0 = -8.0141529e-9
+ lpdiblc2 = -9.0555048e-10
+ wtvfbsdoff = 0
+ ptvoff = 1.3445493e-16
+ waigc = -2.4575845e-11
+ waigsd = 1.9150694e-12
+ ltvfbsdoff = 0
+ lketa = -3.9112692e-9
+ diomod = 1
+ xpart = 1
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.9113600000000002e-10
+ pku0we = 0.0
+ cjswgs = 1.9113600000000002e-10
+ cigbacc = 0.245
+ egidl = 0.001
+ lkvth0we = 3e-12
+ tnoimod = 0
+ mjswgd = 0.95
+ mjswgs = 0.95
+ cigbinv = 0.006
+ tcjswg = 0.00128
+ pvfbsdoff = 0
+ ptvfbsdoff = 0
+ acnqsmod = 0
+ )

.model pch_fs_22 pmos (
+ level = 54
+ xrcrg1 = 12
+ xrcrg2 = 1
+ paramchk = 1
+ rshg = 14.1
+ nfactor = 1
+ wtvoff = 2.0697628e-9
+ ijthdfwd = 0.01
+ capmod = 2
+ tvoff = -0.0031746364
+ tnom = 25
+ wku0we = 1.5e-11
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ mobmod = 0
+ nigbacc = 10
+ ijthdrev = 0.01
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = -1.0531895e-8
+ lpdiblc2 = 0
+ letab = 1.4778454e-8
+ nigbinv = 2.171
+ wags = -2.597049e-7
+ ppclm = 2.5985382e-14
+ wcit = -2.4970451e-10
+ dlcig = 2.5e-9
+ laigsd = 2.2969081e-18
+ bgidl = 1834800000.0
+ voff = -0.11952627
+ acde = 0.5
+ vsat = 226790.48
+ wint = 0
+ vth0 = -0.38544588
+ a0 = 2.9368155
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ wkt1 = -1.289882e-8
+ wkt2 = 2.7006409e-8
+ at = 192293.99
+ cf = 8.17e-11
+ wmax = 9.025999999999999e-7
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.02088367
+ k3 = -2.5823
+ em = 20000000.0
+ fnoimod = 1
+ aigc = 0.0066428307
+ wmin = 5.426e-7
+ ll = 0
+ lw = 0
+ u0 = 0.008363541700000001
+ dmcgt = 0
+ w0 = 0
+ ua = -1.5734149e-9
+ ub = 3.4167628e-18
+ uc = -1.3540772e-10
+ ud = 0
+ tcjsw = 9.34e-5
+ wl = 0
+ lkvth0we = 3e-12
+ wr = 1
+ xj = 1.1e-7
+ eigbinv = 1.1
+ xl = 4e-9
+ ww = 0
+ xw = 3.4e-9
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ wua1 = 6.2697239e-16
+ wub1 = -9.8389336e-25
+ wuc1 = -5.3295995e-16
+ bigc = 0.0012521
+ acnqsmod = 0
+ bigsd = 0.0003327
+ wwlc = 0
+ wvoff = -3.6240027e-9
+ cdsc = 0
+ rbodymod = 0
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigbacc = 0.245
+ wvsat = -0.072832829
+ cigc = 0.15259
+ wvth0 = 4.946536399999999e-9
+ waigc = 3.8715701e-11
+ tnoimod = 0
+ toxref = 3e-9
+ lketa = 1.7736502e-8
+ cigbinv = 0.006
+ xpart = 1
+ wpdiblc2 = 6.2191766e-10
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ egidl = 0.001
+ version = 4.5
+ ltvoff = 2.5685776e-10
+ k2we = 5e-5
+ tempmod = 0
+ dsub = 0.5
+ dtox = 3.91e-10
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ pvfbsdoff = 0
+ aigbacc = 0.012071
+ eta0 = 0.29878005
+ etab = -0.34238426
+ wkvth0we = 0.0
+ lku0we = 1.8e-11
+ epsrox = 3.9
+ trnqsmod = 0
+ rdsmod = 0
+ aigbinv = 0.009974
+ pvoff = 9.4320558e-17
+ igbmod = 1
+ cdscb = 0
+ cdscd = 0
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ pvsat = 5.1892488e-9
+ wk2we = 0.0
+ pvth0 = -9.111998500000001e-16
+ drout = 0.56
+ pbswgd = 0.8
+ pbswgs = 0.8
+ paigc = -2.5833927e-18
+ igcmod = 1
+ voffl = 0
+ rgatemod = 0
+ tnjtsswg = 1
+ weta0 = -7.0544749e-8
+ wetab = 2.4810139e-8
+ lpclm = -5.2812564e-8
+ poxedge = 1
+ cgidl = 1
+ binunit = 2
+ paigsd = -2.080997e-24
+ pbswd = 0.9
+ pbsws = 0.9
+ permod = 1
+ keta = -0.30513509
+ pdits = 0
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ jtsswgd = 1.75e-7
+ lcit = 1.3406861e-10
+ jtsswgs = 1.75e-7
+ voffcv = -0.125
+ wpemod = 1
+ kt1l = 0
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ lint = 0
+ lkt1 = -4.5989262e-9
+ lkt2 = 3.753071e-9
+ lmax = 9e-8
+ lmin = 5.4e-8
+ tnoia = 0
+ lpe0 = 6.44e-8
+ lpeb = 0
+ ijthsfwd = 0.01
+ peta0 = 4.3079228999999995e-15
+ petab = -1.0404991e-15
+ wketa = 1.6222018e-7
+ minv = -0.33
+ wtvfbsdoff = 0
+ lua1 = 1.1693458e-16
+ lub1 = -2.0580342e-25
+ luc1 = -5.5456179e-17
+ tpbsw = 0.0025
+ tpbswg = 0.001
+ ndep = 1e+18
+ cjswd = 5.3856e-11
+ njtsswg = 6.489
+ cjsws = 5.3856e-11
+ mjswd = 0.01
+ lwlc = 0
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ moin = 5.5538
+ ltvfbsdoff = 0
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ ijthsrev = 0.01
+ nigc = 2.291
+ ckappad = 0.6
+ ckappas = 0.6
+ ags = 4.48665
+ pdiblc1 = 0
+ pdiblc2 = 0.0019609567
+ ptvoff = -1.0118352e-16
+ pdiblcb = 0
+ cjd = 0.001421376
+ cit = 0.00026766759
+ waigsd = 1.9150916e-12
+ cjs = 0.001421376
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ noff = 2.2684
+ bvs = 8.2
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ dlc = 4.0349e-9
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ diomod = 1
+ scref = 1e-6
+ ntox = 1.0
+ pcit = -2.2566987e-18
+ pclm = 2.1268063
+ la0 = -1.9926782e-7
+ pditsd = 0
+ pditsl = 0
+ ppdiblc2 = 0
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = -0.0070780887
+ cjswgd = 1.9113600000000002e-10
+ pku0we = 0.0
+ pigcd = 2.572
+ kt1 = -0.26717441
+ cjswgs = 1.9113600000000002e-10
+ kt2 = -0.13819145
+ lk2 = 4.7304354e-9
+ aigsd = 0.0063634181
+ bigbacc = 0.0054401
+ llc = 0
+ ptvfbsdoff = 0
+ lln = 1
+ lu0 = -1.3789508000000001e-10
+ mjd = 0.335
+ mjs = 0.335
+ lua = 6.8530064e-17
+ lub = -1.6632734e-25
+ luc = 7.5845372e-18
+ lud = 0
+ tvfbsdoff = 0.1
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 2.4118768e-14
+ phin = 0.15
+ lvoff = -2.5437461e-9
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 2.0972465e-9
+ pbs = 0.75
+ pk2 = 2.0570947e-16
+ pu0 = 1.8416833e-16
+ kvth0we = -0.00022
+ prt = 0
+ pua = -1.7823119e-23
+ pub = 1.268951e-31
+ puc = -7.4643321e-24
+ pud = 0
+ pkt1 = 2.6462803e-15
+ pkt2 = -1.6460695e-15
+ lvsat = -0.009113146
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = -1.4241889e-9
+ ub1 = 2.5868363e-18
+ mjswgd = 0.95
+ lvth0 = 4.9613109e-10
+ uc1 = 9.3723935e-10
+ mjswgs = 0.95
+ lintnoi = -5e-9
+ tpb = 0.0016
+ wa0 = -5.5297601e-7
+ delta = 0.018814
+ bigbinv = 0.00149
+ ute = -1
+ vtsswgd = 1.1
+ wat = -0.070679454
+ laigc = -9.8025804e-12
+ vtsswgs = 1.1
+ tcjswg = 0.00128
+ web = 6628.3
+ wec = -16935.0
+ wk2 = -1.7106076e-9
+ wlc = 0
+ wln = 1
+ wu0 = -1.5951011e-9
+ xgl = -8.2e-9
+ xgw = 0
+ wua = 2.2095182e-16
+ wub = -1.4911779e-24
+ wuc = 1.1260467e-16
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ rnoia = 0
+ rnoib = 0
+ rbdb = 50
+ pua1 = -5.0424332e-24
+ prwb = 0
+ pub1 = 1.2644812e-32
+ prwg = 0
+ puc1 = 3.7853356e-23
+ pkvth0we = 0.0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ pketa = -1.2596682e-14
+ ngate = 1.7e+20
+ rdsw = 200
+ ngcon = 1
+ wvfbsdoff = 0
+ wpclm = -6.2069351e-7
+ lvfbsdoff = 0
+ vfbsdoff = 0.01
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ fprout = 200
+ )

.model pch_fs_23 pmos (
+ level = 54
+ ijthsfwd = 0.01
+ dtox = 3.91e-10
+ cgidl = 1
+ wku0we = 1.5e-11
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ mobmod = 0
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ eta0 = 7.956713e-6
+ etab = -0.26192508
+ pbswd = 0.9
+ pbsws = 0.9
+ ijthsrev = 0.01
+ pdits = 0
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ ppdiblc2 = 0
+ njtsswg = 6.489
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ tnoia = 0
+ ckappad = 0.6
+ ckappas = 0.6
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ pdiblc1 = 0
+ pdiblc2 = 0.0019609567
+ pdiblcb = 0
+ peta0 = -2.8152439e-15
+ petab = -1.6989745e-15
+ wketa = -4.2902456e-7
+ tpbsw = 0.0025
+ cjswd = 5.3856e-11
+ cjsws = 5.3856e-11
+ pkvth0we = 0.0
+ ags = 4.48665
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ cjd = 0.001421376
+ cit = -0.002877963
+ cjs = 0.001421376
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 4.0349e-9
+ bigbacc = 0.0054401
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ vfbsdoff = 0.01
+ a0 = 5.6551822
+ a1 = 0
+ a2 = 1
+ keta = 0.46798148
+ b0 = 0
+ b1 = 0
+ kvth0we = -0.00022
+ at = -40561.437
+ cf = 8.17e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.018874979
+ k3 = -2.5823
+ em = 20000000.0
+ la0 = -3.569331e-7
+ toxref = 3e-9
+ ll = 0
+ jsd = 1.5e-7
+ lw = 0
+ jss = 1.5e-7
+ lat = 0.0064275263
+ u0 = 0.0073684759
+ w0 = 0
+ kt1 = -0.46532049
+ kt2 = 0.0072316444
+ lk2 = 4.6139313e-9
+ ua = 5.3944309e-9
+ ub = -7.8004593e-18
+ uc = 1.0922891e-10
+ ud = 0
+ llc = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ lln = 1
+ xw = 3.4e-9
+ lu0 = -8.018127e-11
+ mjd = 0.335
+ lintnoi = -5e-9
+ mjs = 0.335
+ lua = -3.3560499e-16
+ lub = 4.8427154e-25
+ luc = -6.604387e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ bigbinv = 0.00149
+ njs = 1.02
+ pa0 = 1.517818e-13
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ nsd = 1e+20
+ lcit = 3.1651519e-10
+ pbd = 0.75
+ pat = -1.8496379e-9
+ pbs = 0.75
+ pk2 = 4.9657487e-16
+ paramchk = 1
+ pu0 = -8.1141216e-17
+ scref = 1e-6
+ kt1l = 0
+ prt = 0
+ pua = 1.7043409e-22
+ pub = -3.4061954e-31
+ puc = 5.8491101e-24
+ pud = 0
+ pigcd = 2.572
+ rsh = 15.2
+ aigsd = 0.0063634182
+ tcj = 0.000832
+ ua1 = 9.464156e-9
+ tvfbsdoff = 0.1
+ ub1 = -1.352433e-17
+ uc1 = -1.5339544e-9
+ tpb = 0.0016
+ wa0 = -2.7540628e-6
+ lint = 0
+ ute = -1
+ wat = -0.002629722
+ lvoff = -5.520199e-9
+ web = 6628.3
+ wec = -16935.0
+ wk2 = -6.7255282e-9
+ wlc = 0
+ wln = 1
+ lkt1 = 6.8935466e-9
+ lkt2 = -4.6814687e-9
+ wu0 = 2.9792015e-9
+ xgl = -8.2e-9
+ xgw = 0
+ ltvoff = -2.6406105e-10
+ wua = -3.0248621e-15
+ wub = 6.5694194e-24
+ wuc = -1.1693744e-16
+ wud = 0
+ lmax = 5.4e-8
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ lmin = 4.5e-8
+ lvsat = 0.0051221042
+ lpe0 = 6.44e-8
+ lvth0 = -6.9814368e-9
+ lpeb = 0
+ ijthdfwd = 0.01
+ delta = 0.018814
+ laigc = -1.6050622e-11
+ minv = -0.33
+ lua1 = -5.1458943e-16
+ lub1 = 7.2864421e-25
+ luc1 = 8.7873061e-17
+ rnoia = 0
+ rnoib = 0
+ ndep = 1e+18
+ lku0we = 1.8e-11
+ lwlc = 0
+ epsrox = 3.9
+ moin = 5.5538
+ pketa = 2.1695512e-14
+ ngate = 1.7e+20
+ wvfbsdoff = 0
+ ijthdrev = 0.01
+ lvfbsdoff = 0
+ ngcon = 1
+ nigc = 2.291
+ wpclm = -1.0386396e-6
+ nfactor = 1
+ rdsmod = 0
+ igbmod = 1
+ lpdiblc2 = 0
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ noff = 2.2684
+ pscbe1 = 926400000.0
+ noia = 2.86e+42
+ pscbe2 = 1e-20
+ noib = 2.5e+24
+ noic = 31000000000.0
+ pbswgd = 0.8
+ pbswgs = 0.8
+ igcmod = 1
+ ntox = 1.0
+ pcit = -4.4191024e-17
+ pclm = 4.4879115
+ nigbacc = 10
+ phin = 0.15
+ lkvth0we = 3e-12
+ pkt1 = -5.1012735999999995e-15
+ pkt2 = 1.1767646e-15
+ nigbinv = 2.171
+ tvoff = 0.0058067224
+ acnqsmod = 0
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ rbdb = 50
+ pua1 = 2.7224008e-22
+ prwb = 0
+ pub1 = -3.6990718e-31
+ prwg = 0
+ puc1 = -5.7927018e-23
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ permod = 1
+ rbodymod = 0
+ rdsw = 200
+ ku0we = -0.0007
+ beta0 = 13.32
+ fnoimod = 1
+ leta0 = 6.7968866e-9
+ letab = 1.0111821e-8
+ eigbinv = 1.1
+ ppclm = 5.0226256e-14
+ voffcv = -0.125
+ wpemod = 1
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ rshg = 14.1
+ wtvfbsdoff = 0
+ wpdiblc2 = 6.2191766e-10
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ ltvfbsdoff = 0
+ cigbacc = 0.245
+ tnoimod = 0
+ tnom = 25
+ tpbswg = 0.001
+ bigsd = 0.0003327
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ cigbinv = 0.006
+ wkvth0we = 0.0
+ wvoff = -2.1208799e-8
+ trnqsmod = 0
+ wvsat = 0.09105966
+ ptvoff = 1.2747838e-16
+ ptvfbsdoff = 0
+ wvth0 = -3.9555008e-8
+ waigsd = 1.9150557e-12
+ version = 4.5
+ waigc = -1.4751759e-11
+ wags = -2.597049e-7
+ tempmod = 0
+ wcit = 4.7330111e-10
+ diomod = 1
+ voff = -0.068208113
+ lketa = -2.7104259e-8
+ acde = 0.5
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.9113600000000002e-10
+ pku0we = 0.0
+ cjswgs = 1.9113600000000002e-10
+ aigbacc = 0.012071
+ xpart = 1
+ rgatemod = 0
+ vsat = -18644.867
+ wint = 0
+ vth0 = -0.2565223
+ tnjtsswg = 1
+ wkt1 = 1.206797e-7
+ wkt2 = -2.1663145e-8
+ egidl = 0.001
+ wmax = 9.025999999999999e-7
+ aigc = 0.0067505556
+ wmin = 5.426e-7
+ mjswgd = 0.95
+ mjswgs = 0.95
+ aigbinv = 0.009974
+ tcjswg = 0.00128
+ pvfbsdoff = 0
+ wua1 = -4.1537606e-15
+ wub1 = 5.6118307e-24
+ wuc1 = 1.1184258e-15
+ bigc = 0.0012521
+ wwlc = 0
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigc = 0.15259
+ pvoff = 1.1142388e-15
+ poxedge = 1
+ cdscb = 0
+ cdscd = 0
+ fprout = 200
+ pvsat = -4.3165155e-9
+ wk2we = 0.0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ pvth0 = 1.6698897e-15
+ drout = 0.56
+ binunit = 2
+ paigc = 5.1772001e-19
+ voffl = 0
+ dmcg = 3.1e-8
+ wtvoff = -1.8726837e-9
+ dmci = 3.1e-8
+ dmdg = 0
+ weta0 = 5.2268470999999997e-8
+ wetab = 3.6163164e-8
+ lpclm = -1.8975667e-7
+ k2we = 5e-5
+ capmod = 2
+ dsub = 0.5
+ )

.model pch_fs_24 pmos (
+ level = 54
+ beta0 = 13.32
+ leta0 = -2.4191759999999978e-11
+ letab = 2.8639817e-9
+ cigbacc = 0.245
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ ppclm = -6.983762e-15
+ laigsd = -1.7489044e-14
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ tnoimod = 0
+ ntox = 1.0
+ pcit = -2.4019874999999997e-16
+ pclm = 0.55996802
+ rgatemod = 0
+ cigbinv = 0.006
+ tnjtsswg = 1
+ phin = 0.15
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ pkt1 = 8.0039909e-15
+ pkt2 = -6.3201272e-16
+ version = 4.5
+ tempmod = 0
+ bigsd = 0.0003327
+ rbdb = 50
+ pua1 = -2.7866327e-22
+ prwb = 0
+ pub1 = 3.2786288e-31
+ prwg = 0
+ puc1 = 2.5974765e-23
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ aigbacc = 0.012071
+ wvoff = -2.6959456e-8
+ rdsw = 200
+ wvsat = 0.037826603
+ wvth0 = -7.2775681e-9
+ toxref = 3e-9
+ waigc = -9.7737582e-11
+ aigbinv = 0.009974
+ lketa = 1.4220453e-8
+ rshg = 14.1
+ xpart = 1
+ egidl = 0.001
+ ltvoff = -2.5344658e-10
+ pvfbsdoff = 0
+ ijthsfwd = 0.01
+ poxedge = 1
+ a0 = -2.5402778
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ tnom = 25
+ at = 213109.93
+ cf = 8.17e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.022656115
+ k3 = -2.5823
+ em = 20000000.0
+ lku0we = 1.8e-11
+ ll = 0
+ lw = 0
+ u0 = 0.0014778574
+ w0 = 0
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ ua = -6.0379704e-9
+ ub = 8.1069989e-18
+ uc = -2.2784413e-10
+ ud = 0
+ binunit = 2
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ epsrox = 3.9
+ xw = 3.4e-9
+ ijthsrev = 0.01
+ rdsmod = 0
+ igbmod = 1
+ pvoff = 1.396021e-15
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ wags = -2.597049e-7
+ cdscb = 0
+ cdscd = 0
+ pbswgd = 0.8
+ pbswgs = 0.8
+ pvsat = -1.7080957e-9
+ wcit = 4.4734589e-9
+ wk2we = 0.0
+ pvth0 = 8.829517000000001e-17
+ drout = 0.56
+ igcmod = 1
+ voff = -0.080254273
+ paigc = 4.5840253e-18
+ acde = 0.5
+ ppdiblc2 = 0
+ voffl = 0
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ vsat = 78763.66
+ wint = 0
+ vth0 = -0.37915952
+ wkt1 = -1.4677468e-7
+ wkt2 = 1.5250678e-8
+ wmax = 9.025999999999999e-7
+ weta0 = -2.1457527999999998e-8
+ aigc = 0.0066531108
+ wetab = 8.325777e-9
+ wmin = 5.426e-7
+ lpclm = 2.7125638e-9
+ cgidl = 1
+ paigsd = 9.5490179e-21
+ wua1 = 7.089165e-15
+ wub1 = -8.6283747e-24
+ wuc1 = -5.9385548e-16
+ bigc = 0.0012521
+ wwlc = 0
+ pkvth0we = 0.0
+ permod = 1
+ cdsc = 0
+ pbswd = 0.9
+ pbsws = 0.9
+ njtsswg = 6.489
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ wtvfbsdoff = 0
+ cigc = 0.15259
+ vfbsdoff = 0.01
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ ckappad = 0.6
+ ckappas = 0.6
+ pdits = 0
+ voffcv = -0.125
+ wpemod = 1
+ pdiblc1 = 0
+ pdiblc2 = 0.0019609567
+ cigsd = 0.013281
+ ltvfbsdoff = 0
+ pdiblcb = 0
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ paramchk = 1
+ pk2we = 0.0
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ bigbacc = 0.0054401
+ tnoia = 0
+ k2we = 5e-5
+ ags = 4.48665
+ ijthdfwd = 0.01
+ dsub = 0.5
+ dtox = 3.91e-10
+ kvth0we = -0.00022
+ peta0 = 7.973300400000001e-16
+ ptvfbsdoff = 0
+ petab = -3.349425e-16
+ cjd = 0.001421376
+ cit = -0.010137593
+ cjs = 0.001421376
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dvt0 = 3.48
+ tpbswg = 0.001
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ wketa = 1.6324308e-7
+ dlc = 4.0349e-9
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ tpbsw = 0.0025
+ dwg = 0
+ lintnoi = -5e-9
+ dwj = 0
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ cjswd = 5.3856e-11
+ cjsws = 5.3856e-11
+ mjswd = 0.01
+ eta0 = 0.13921364
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ etab = -0.11400999
+ la0 = 4.4644444e-8
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = -0.0060023707
+ kt1 = 0.16833478
+ kt2 = -0.11193164
+ lk2 = 4.7992069999999995e-9
+ ijthdrev = 0.01
+ llc = 0
+ lln = 1
+ lu0 = 2.0845903999999999e-10
+ mjd = 0.335
+ ptvoff = 8.5019581e-17
+ mjs = 0.335
+ lua = 2.2458267e-16
+ lub = -2.9519392e-25
+ luc = 9.9121919e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = -8.9774533e-14
+ waigsd = 1.7201778e-12
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 6.8793549e-9
+ pbs = 0.75
+ lpdiblc2 = 0
+ pk2 = 1.0702031e-16
+ pu0 = -9.6657248e-17
+ prt = 0
+ pua = -9.0705467e-23
+ pub = 1.0841652e-31
+ puc = -1.0416838e-23
+ pud = 0
+ diomod = 1
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = -1.018181e-8
+ ub1 = 1.2390462e-17
+ uc1 = 9.111363e-10
+ tpb = 0.0016
+ wa0 = 2.1756583e-6
+ ute = -1
+ wat = -0.18077244
+ pditsd = 0
+ web = 6628.3
+ wec = -16935.0
+ pditsl = 0
+ wk2 = 1.2245648e-9
+ cjswgd = 1.9113600000000002e-10
+ pku0we = 0.0
+ cjswgs = 1.9113600000000002e-10
+ wlc = 0
+ wln = 1
+ wu0 = 3.2958552e-9
+ xgl = -8.2e-9
+ xgw = 0
+ scref = 1e-6
+ wua = 2.3045166e-15
+ wub = -2.5945817e-24
+ wuc = 2.150207e-16
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ tvfbsdoff = 0.1
+ pigcd = 2.572
+ aigsd = 0.0063637751
+ lvoff = -4.9299372e-9
+ mjswgd = 0.95
+ mjswgs = 0.95
+ lkvth0we = 3e-12
+ nfactor = 1
+ lvsat = 0.00034908628
+ tcjswg = 0.00128
+ lvth0 = -9.7221299e-10
+ delta = 0.018814
+ laigc = -1.1275829e-11
+ acnqsmod = 0
+ rnoia = 0
+ rnoib = 0
+ wvfbsdoff = 0
+ pketa = -7.3256019e-15
+ ngate = 1.7e+20
+ lvfbsdoff = 0
+ rbodymod = 0
+ nigbacc = 10
+ ngcon = 1
+ wpclm = 1.2891178e-7
+ gbmin = 1e-12
+ keta = -0.37538
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ fprout = 200
+ xrcrg1 = 12
+ xrcrg2 = 1
+ nigbinv = 2.171
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 6.722370400000001e-10
+ kt1l = 0
+ wtvoff = -1.0061777e-9
+ wpdiblc2 = 6.2191766e-10
+ lint = 0
+ lkt1 = -2.4155560999999997e-8
+ lkt2 = 1.1575324e-9
+ lmax = 4.5e-8
+ lmin = 3.6e-8
+ capmod = 2
+ fnoimod = 1
+ lpe0 = 6.44e-8
+ lpeb = 0
+ wku0we = 1.5e-11
+ eigbinv = 1.1
+ tvoff = 0.0055901005
+ mobmod = 0
+ minv = -0.33
+ lua1 = 4.4806289e-16
+ lub1 = -5.4118058e-25
+ luc1 = -3.1936385e-17
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ ndep = 1e+18
+ wkvth0we = 0.0
+ lwlc = 0
+ moin = 5.5538
+ nigc = 2.291
+ trnqsmod = 0
+ ku0we = -0.0007
+ )

.model pch_fs_25 pmos (
+ level = 54
+ wint = 0
+ ags = 0.93810347
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ vth0 = -0.40198248000000003
+ wkt1 = -1.5318394e-9
+ wkt2 = 2.21858e-9
+ cjd = 0.001421376
+ cit = 5e-6
+ cjs = 0.001421376
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ wmax = 5.426e-7
+ bvs = 8.2
+ aigc = 0.0068215676
+ wmin = 2.726e-7
+ dlc = 1.0572421799999999e-8
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ k3b = 2.1176
+ lkvth0we = 3e-12
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ tnoia = 0
+ peta0 = -1.6e-17
+ la0 = 0
+ wua1 = 1.6452204e-16
+ wub1 = -6.9710259e-26
+ wuc1 = 2.1709154e-17
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0.00064
+ wketa = 2.2687563e-8
+ kt1 = -0.17747938
+ lk2 = 3.2000000000000003e-10
+ kt2 = -0.061438333
+ llc = 0
+ lln = 1
+ lu0 = -8e-13
+ tpbsw = 0.0025
+ acnqsmod = 0
+ mjd = 0.335
+ bigc = 0.0012521
+ mjs = 0.335
+ wute = 3.2371733e-8
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ wwlc = 0
+ pa0 = 0
+ cjswd = 5.3856e-11
+ nsd = 1e+20
+ cjsws = 5.3856e-11
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ pk2 = 0
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ pu0 = 0
+ prt = 0
+ pud = 0
+ rbodymod = 0
+ cdsc = 0
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 1.8507467e-10
+ ub1 = -1.7337534e-19
+ uc1 = -4.0886356e-11
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ tpb = 0.0016
+ wa0 = -1.5013787e-7
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigc = 0.15259
+ ute = -1.2102889
+ toxref = 3e-9
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 4.440518e-10
+ wlc = 0
+ wln = 1
+ wu0 = 3.7953067e-11
+ xgl = -8.2e-9
+ xgw = 0
+ nfactor = 1
+ wua = -1.5196107e-16
+ wub = 9.0507286e-26
+ wuc = 5.3799588e-18
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ scref = 1e-6
+ tvfbsdoff = 0.1
+ pigcd = 2.572
+ aigsd = 0.0063632886
+ wpdiblc2 = -7.7579138e-11
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ ltvoff = 0
+ lvoff = 0
+ nigbacc = 10
+ lvsat = 8.000000000000001e-6
+ k2we = 5e-5
+ lvth0 = -2.4e-10
+ dsub = 0.5
+ dtox = 3.91e-10
+ delta = 0.018814
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ lku0we = 1.8e-11
+ rnoia = 0
+ rnoib = 0
+ epsrox = 3.9
+ nigbinv = 2.171
+ eta0 = 0.17962267
+ wvfbsdoff = 0
+ wkvth0we = 0.0
+ etab = -0.19577778
+ lvfbsdoff = 0
+ ngate = 1.7e+20
+ rdsmod = 0
+ ngcon = 1
+ igbmod = 1
+ wpclm = -1.1447315e-8
+ trnqsmod = 0
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ pbswgd = 0.8
+ pbswgs = 0.8
+ fnoimod = 1
+ eigbinv = 1.1
+ igcmod = 1
+ a0 = 3.3089778
+ a1 = 0
+ a2 = 1
+ rgatemod = 0
+ b0 = 0
+ b1 = 0
+ at = 72000
+ cf = 8.17e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.0028441163
+ k3 = -2.5823
+ em = 20000000.0
+ tnjtsswg = 1
+ ll = 0
+ lw = 0
+ u0 = 0.0097214889
+ w0 = 0
+ ua = 1.8228697e-10
+ ub = 9.7616315e-19
+ uc = -9.1826044e-12
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 3.4e-9
+ wtvfbsdoff = 0
+ cigbacc = 0.245
+ tvoff = 0.0026578776
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ permod = 1
+ ltvfbsdoff = 0
+ tnoimod = 0
+ cigbinv = 0.006
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = -4.8e-10
+ keta = -0.064397096
+ voffcv = -0.125
+ wpemod = 1
+ ppclm = 0
+ version = 4.5
+ dlcig = 2.5e-9
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ bgidl = 1834800000.0
+ lcit = 1.6e-11
+ tempmod = 0
+ ptvfbsdoff = 0
+ kt1l = 0
+ aigbacc = 0.012071
+ lint = 6.5375218e-9
+ dmcgt = 0
+ lkt1 = -4.8e-10
+ tcjsw = 9.34e-5
+ lmax = 2.001e-5
+ lmin = 8.9991e-6
+ lpe0 = 6.44e-8
+ lpeb = 0
+ ijthsfwd = 0.01
+ tpbswg = 0.001
+ minv = -0.33
+ aigbinv = 0.009974
+ bigsd = 0.0003327
+ ndep = 1e+18
+ lwlc = 0
+ moin = 5.5538
+ wvoff = 2.5521431e-9
+ ptvoff = 0
+ ijthsrev = 0.01
+ nigc = 2.291
+ waigsd = 1.9763167e-12
+ wvsat = 0.0034765009
+ wvth0 = -3.974714700000001e-9
+ diomod = 1
+ waigc = 4.045116e-12
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.9113600000000002e-10
+ pku0we = 0.0
+ cjswgs = 1.9113600000000002e-10
+ poxedge = 1
+ lketa = 0
+ ntox = 1.0
+ xpart = 1
+ pcit = -8.000000000000001e-19
+ pclm = 1.1689658
+ ppdiblc2 = 0
+ binunit = 2
+ egidl = 0.001
+ mjswgd = 0.95
+ mjswgs = 0.95
+ phin = 0.15
+ tcjswg = 0.00128
+ pkt1 = -4e-17
+ pvfbsdoff = 0
+ rbdb = 50
+ prwb = 0
+ prwg = 0
+ pkvth0we = 0.0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ jtsswgd = 1.75e-7
+ rdsw = 200
+ jtsswgs = 1.75e-7
+ vfbsdoff = 0.01
+ fprout = 200
+ pvoff = 2e-17
+ xrcrg1 = 12
+ xrcrg2 = 1
+ cdscb = 0
+ cdscd = 0
+ pvsat = 0
+ wk2we = 0.0
+ pvth0 = -1.2e-16
+ drout = 0.56
+ paramchk = 1
+ wtvoff = -1.0551434e-10
+ rshg = 14.1
+ voffl = 0
+ weta0 = -1.7872176e-8
+ wetab = 1.9534667e-8
+ njtsswg = 6.489
+ capmod = 2
+ lpclm = 0
+ wku0we = 1.5e-11
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ ijthdfwd = 0.01
+ cgidl = 1
+ mobmod = 0
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.0030491463
+ tnom = 25
+ pdiblcb = 0
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ pbswd = 0.9
+ pbsws = 0.9
+ ijthdrev = 0.01
+ lpdiblc2 = 0
+ bigbacc = 0.0054401
+ wags = -6.1953916e-9
+ pdits = 0
+ cigsd = 0.013281
+ kvth0we = -0.00022
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ voff = -0.10784306
+ acde = 0.5
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ vsat = 91103.982
+ pk2we = 0.0
+ )

.model pch_fs_26 pmos (
+ level = 54
+ bigsd = 0.0003327
+ poxedge = 1
+ pkvth0we = 0.0
+ wvoff = 2.9007224e-9
+ binunit = 2
+ toxref = 3e-9
+ wvsat = 0.0034765009
+ wvth0 = -4.0362892e-9
+ vfbsdoff = 0.01
+ keta = -0.06875265
+ waigc = 4.3476029e-12
+ lags = 1.0877241e-7
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 1.6e-11
+ lketa = 3.9156432e-8
+ paramchk = 1
+ kt1l = 0
+ xpart = 1
+ ltvoff = -4.4286369e-10
+ egidl = 0.001
+ lint = 6.5375218e-9
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ lkt1 = -3.5333729e-8
+ lkt2 = -1.4641311e-8
+ lmax = 8.9991e-6
+ pvfbsdoff = 0
+ lmin = 8.9908e-7
+ lpe0 = 6.44e-8
+ ijthdfwd = 0.01
+ lpeb = 0
+ lku0we = 1.8e-11
+ minv = -0.33
+ epsrox = 3.9
+ lua1 = 1.4818924e-15
+ lub1 = -2.0711788e-24
+ luc1 = 2.2491171e-16
+ ndep = 1e+18
+ lute = 1.330224e-7
+ rdsmod = 0
+ lwlc = 0
+ moin = 5.5538
+ igbmod = 1
+ ijthdrev = 0.01
+ nigc = 2.291
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ lpdiblc2 = 8.2033961e-9
+ njtsswg = 6.489
+ pbswgd = 0.8
+ pvoff = -3.1137282e-15
+ pbswgs = 0.8
+ noff = 2.2684
+ cdscb = 0
+ cdscd = 0
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ igcmod = 1
+ pvsat = 0
+ wk2we = 0.0
+ pvth0 = 4.3355474000000005e-16
+ drout = 0.56
+ ckappad = 0.6
+ ckappas = 0.6
+ pags = 8.2314292e-14
+ wtvfbsdoff = 0
+ pdiblc1 = 0
+ pdiblc2 = 0.002136644
+ paigc = -2.7193569e-18
+ pdiblcb = 0
+ ntox = 1.0
+ pcit = -8.000000000000001e-19
+ pclm = 1.1689658
+ voffl = 0
+ ltvfbsdoff = 0
+ weta0 = -1.7872176e-8
+ phin = 0.15
+ wetab = 1.9534667e-8
+ lkvth0we = 3e-12
+ lpclm = 0
+ paigsd = -4.5957918e-20
+ pkt1 = 4.5192526e-15
+ pkt2 = 3.8774237e-15
+ bigbacc = 0.0054401
+ cgidl = 1
+ permod = 1
+ acnqsmod = 0
+ kvth0we = -0.00022
+ rbdb = 50
+ pua1 = -9.4343892e-23
+ prwb = 0
+ pub1 = 9.0084871e-32
+ prwg = 0
+ puc1 = -7.238167e-23
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ lintnoi = -5e-9
+ pute = -1.6539558e-14
+ bigbinv = 0.00149
+ rbodymod = 0
+ pbswd = 0.9
+ pbsws = 0.9
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ rdsw = 200
+ ptvfbsdoff = 0
+ a0 = 3.4253346
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 72000
+ cf = 8.17e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.0024652651
+ k3 = -2.5823
+ em = 20000000.0
+ ll = 0
+ voffcv = -0.125
+ lw = 0
+ wpemod = 1
+ u0 = 0.0096054275
+ w0 = 0
+ ua = 1.8429003e-10
+ ub = 9.3982253e-19
+ uc = -1.1498405e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 3.4e-9
+ pdits = 0
+ cigsd = 0.013281
+ ags = 0.9260042
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ cjd = 0.001421376
+ cit = 5e-6
+ cjs = 0.001421376
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 1.0572421799999999e-8
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ rshg = 14.1
+ wpdiblc2 = 3.818702e-12
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ la0 = -1.0460478e-6
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0.00064
+ kt1 = -0.17360244
+ kt2 = -0.059809712
+ lk2 = -3.0858721e-9
+ llc = 0
+ lln = 1
+ lu0 = 1.0425917e-9
+ mjd = 0.335
+ mjs = 0.335
+ lua = -1.8007487e-17
+ lub = 3.2670219e-25
+ luc = 2.0819042e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ tnoia = 0
+ njd = 1.02
+ njs = 1.02
+ pa0 = 1.483047e-13
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ tpbswg = 0.001
+ pk2 = 2.5596912e-15
+ pu0 = 1.7642195e-17
+ nfactor = 1
+ peta0 = -1.6e-17
+ prt = 0
+ pua = 1.2819791e-23
+ pub = -1.2787603e-32
+ puc = -1.6865938e-24
+ pud = 0
+ wketa = 2.5468383e-8
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 2.0236805e-11
+ ub1 = 5.7011626e-20
+ uc1 = -6.5904343e-11
+ tnom = 25
+ tpbsw = 0.0025
+ tpb = 0.0016
+ wa0 = -1.666345e-7
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ ute = -1.2250856
+ cjswd = 5.3856e-11
+ cjsws = 5.3856e-11
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 1.5932531e-10
+ mjswd = 0.01
+ wlc = 0
+ mjsws = 0.01
+ wln = 1
+ agidl = 3.2166e-9
+ wu0 = 3.5990642e-11
+ wkvth0we = 0.0
+ xgl = -8.2e-9
+ xgw = 0
+ wua = -1.5338707e-16
+ wub = 9.1929712e-26
+ wuc = 5.5675666e-18
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ ptvoff = -2.4168192e-17
+ waigsd = 1.9814288e-12
+ trnqsmod = 0
+ nigbacc = 10
+ diomod = 1
+ wags = -1.5351598e-8
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.9113600000000002e-10
+ pku0we = 0.0
+ cjswgs = 1.9113600000000002e-10
+ tvfbsdoff = 0.1
+ voff = -0.10676035
+ scref = 1e-6
+ acde = 0.5
+ nigbinv = 2.171
+ pigcd = 2.572
+ rgatemod = 0
+ aigsd = 0.0063632773
+ vsat = 91103.982
+ wint = 0
+ vth0 = -0.40056355000000005
+ tnjtsswg = 1
+ mjswgd = 0.95
+ mjswgs = 0.95
+ wkt1 = -2.0389865e-9
+ wkt2 = 1.7872759e-9
+ lvoff = -9.7335308e-9
+ wmax = 5.426e-7
+ aigc = 0.0068257672
+ wmin = 2.726e-7
+ tcjswg = 0.00128
+ lvsat = 8.000000000000001e-6
+ lvth0 = -1.2996137e-8
+ delta = 0.018814
+ laigc = -3.7754415e-11
+ wua1 = 1.7501635e-16
+ wub1 = -7.9730823e-26
+ wuc1 = 2.9760508e-17
+ fnoimod = 1
+ rnoia = 0
+ rnoib = 0
+ bigc = 0.0012521
+ eigbinv = 1.1
+ wute = 3.4211506e-8
+ wwlc = 0
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ pketa = -2.4999571e-14
+ ngate = 1.7e+20
+ cdsc = 0
+ ngcon = 1
+ cgbo = 0
+ wpclm = -1.1447315e-8
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ fprout = 200
+ cigc = 0.15259
+ gbmin = 1e-12
+ xrcrg1 = 12
+ xrcrg2 = 1
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ cigbacc = 0.245
+ wtvoff = -1.02826e-10
+ tnoimod = 0
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ capmod = 2
+ cigbinv = 0.006
+ wku0we = 1.5e-11
+ k2we = 5e-5
+ mobmod = 0
+ ijthsfwd = 0.01
+ dsub = 0.5
+ dtox = 3.91e-10
+ tvoff = 0.0027071394
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ xjbvd = 1
+ xjbvs = 1
+ version = 4.5
+ lk2we = 0.0
+ tempmod = 0
+ eta0 = 0.17962267
+ etab = -0.19577778
+ ijthsrev = 0.01
+ ku0we = -0.0007
+ aigbacc = 0.012071
+ beta0 = 13.32
+ leta0 = -4.8e-10
+ laigsd = 1.0132005e-13
+ ppclm = 0
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ aigbinv = 0.009974
+ ppdiblc2 = -7.3176658e-16
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ )

.model pch_fs_27 pmos (
+ level = 54
+ tvfbsdoff = 0.1
+ fnoimod = 1
+ scref = 1e-6
+ eigbinv = 1.1
+ rshg = 14.1
+ ltvoff = -3.7535707e-10
+ pigcd = 2.572
+ aigsd = 0.0063633912
+ lvoff = -1.1639377e-8
+ lvsat = 8.000000000000001e-6
+ lvth0 = 8.106701000000001e-10
+ ijthsfwd = 0.01
+ lku0we = 1.8e-11
+ delta = 0.018814
+ laigc = -5.5983746e-11
+ epsrox = 3.9
+ tnom = 25
+ rnoia = 0
+ rnoib = 0
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ cigbacc = 0.245
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ rdsmod = 0
+ igbmod = 1
+ pketa = 5.6398736e-15
+ ngate = 1.7e+20
+ wtvfbsdoff = 0
+ ijthsrev = 0.01
+ ngcon = 1
+ tnoimod = 0
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ wpclm = -1.1447315e-8
+ pbswgd = 0.8
+ pbswgs = 0.8
+ gbmin = 1e-12
+ cigbinv = 0.006
+ jswgd = 3.69e-13
+ ltvfbsdoff = 0
+ jswgs = 3.69e-13
+ igcmod = 1
+ wags = 3.4820603e-7
+ voff = -0.10461895
+ acde = 0.5
+ version = 4.5
+ ppdiblc2 = 9.4893758e-16
+ vsat = 91103.982
+ tempmod = 0
+ wint = 0
+ vth0 = -0.41607682
+ wkt1 = 1.4552168e-8
+ wkt2 = 6.9668931e-9
+ wmax = 5.426e-7
+ aigc = 0.0068462496
+ wmin = 2.726e-7
+ aigbacc = 0.012071
+ ptvfbsdoff = 0
+ tvoff = 0.0026312893
+ wua1 = 1.777316e-16
+ wub1 = 1.5048515e-26
+ wuc1 = -3.1929257e-17
+ permod = 1
+ xjbvd = 1
+ xjbvs = 1
+ bigc = 0.0012521
+ wute = 6.965504e-8
+ lk2we = 0.0
+ wwlc = 0
+ pkvth0we = 0.0
+ aigbinv = 0.009974
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ ku0we = -0.0007
+ beta0 = 13.32
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ voffcv = -0.125
+ wpemod = 1
+ cigc = 0.15259
+ vfbsdoff = 0.01
+ leta0 = -4.8e-10
+ ppclm = 0
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ paramchk = 1
+ poxedge = 1
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ binunit = 2
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ tpbswg = 0.001
+ k2we = 5e-5
+ ijthdfwd = 0.01
+ dsub = 0.5
+ dtox = 3.91e-10
+ a0 = 2.4559917
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 72000
+ cf = 8.17e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.0065510297
+ k3 = -2.5823
+ em = 20000000.0
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ ll = 0
+ lw = 0
+ u0 = 0.011139968
+ w0 = 0
+ ua = 2.2475737e-10
+ ub = 1.3971204e-18
+ uc = 8.9671176e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 3.4e-9
+ bigsd = 0.0003327
+ ptvoff = 6.0034078e-17
+ eta0 = 0.17962267
+ etab = -0.19577778
+ waigsd = 1.9297907e-12
+ wvoff = -2.3606869e-9
+ ijthdrev = 0.01
+ wvsat = 0.0034765009
+ diomod = 1
+ wvth0 = -3.2767848000000002e-9
+ lpdiblc2 = -1.0873556e-9
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ waigc = -6.0221967e-12
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.9113600000000002e-10
+ pku0we = 0.0
+ cjswgs = 1.9113600000000002e-10
+ lketa = -2.7133526e-8
+ xpart = 1
+ mjswgd = 0.95
+ mjswgs = 0.95
+ egidl = 0.001
+ tcjswg = 0.00128
+ pvfbsdoff = 0
+ lkvth0we = 3e-12
+ njtsswg = 6.489
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ acnqsmod = 0
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.012575691
+ pdiblcb = 0
+ rbodymod = 0
+ fprout = 200
+ xrcrg1 = 12
+ xrcrg2 = 1
+ pvoff = 1.5689261e-15
+ keta = 0.0057304489
+ cdscb = 0
+ cdscd = 0
+ pvsat = 0
+ bigbacc = 0.0054401
+ lags = 9.833094e-7
+ wk2we = 0.0
+ pvth0 = -2.4240418e-16
+ wtvoff = -1.9743529e-10
+ drout = 0.56
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 9.8671111e-11
+ paigc = 6.5097646e-18
+ kt1l = 0
+ kvth0we = -0.00022
+ voffl = 0
+ wpdiblc2 = -1.8846129e-9
+ lintnoi = -5e-9
+ capmod = 2
+ lint = 6.5375218e-9
+ bigbinv = 0.00149
+ weta0 = -1.7872176e-8
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ wetab = 1.9534667e-8
+ wku0we = 1.5e-11
+ lkt1 = -4.8129349e-9
+ lkt2 = -2.567581e-9
+ lpclm = 0
+ lmax = 8.9908e-7
+ lmin = 4.4908e-7
+ mobmod = 0
+ lpe0 = 6.44e-8
+ lpeb = 0
+ cgidl = 1
+ minv = -0.33
+ lua1 = 1.3348283e-16
+ lub1 = 2.1611253e-25
+ luc1 = 5.928335e-17
+ ndep = 1e+18
+ lute = 1.2896693e-7
+ wkvth0we = 0.0
+ lwlc = 0
+ moin = 5.5538
+ pbswd = 0.9
+ pbsws = 0.9
+ ags = -0.056621626
+ nigc = 2.291
+ trnqsmod = 0
+ cjd = 0.001421376
+ cit = -8.7888889e-5
+ cjs = 0.001421376
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 1.0572421799999999e-8
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ pdits = 0
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ cigsd = 0.013281
+ nfactor = 1
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ la0 = -1.8333262e-7
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0.00064
+ pags = -2.41252e-13
+ kt1 = -0.20789546
+ kt2 = -0.0733757
+ lk2 = 5.5045842e-10
+ llc = 0
+ lln = 1
+ lu0 = -3.2314965e-10
+ mjd = 0.335
+ mjs = 0.335
+ lua = -5.402342e-17
+ lub = -8.029291e-26
+ luc = -6.9221885e-17
+ lud = 0
+ ntox = 1.0
+ lwc = 0
+ lwl = 0
+ pcit = -8.000000000000001e-19
+ lwn = 1
+ pclm = 1.1689658
+ njd = 1.02
+ njs = 1.02
+ pa0 = -1.295362e-13
+ rgatemod = 0
+ nsd = 1e+20
+ pbd = 0.75
+ pk2we = 0.0
+ pat = 0
+ pbs = 0.75
+ pk2 = 6.34174e-16
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ tnjtsswg = 1
+ pu0 = -2.5304972e-16
+ prt = 0
+ pua = -1.1377853e-22
+ pub = 1.1787175e-31
+ puc = 2.8393052e-23
+ pud = 0
+ phin = 0.15
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 1.5353037e-9
+ ub1 = -2.5129786e-18
+ uc1 = 1.2019494e-10
+ tpb = 0.0016
+ tnoia = 0
+ wa0 = 1.4554629e-7
+ pkt1 = -1.0246874e-14
+ pkt2 = -7.3243565e-16
+ ute = -1.2205289
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 2.3228278e-9
+ nigbacc = 10
+ wlc = 0
+ wln = 1
+ wu0 = 3.4013886e-10
+ xgl = -8.2e-9
+ xgw = 0
+ peta0 = -1.6e-17
+ wua = -1.1141771e-17
+ wub = -5.4878553e-26
+ wuc = -2.8229789e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ wketa = -8.9579586e-9
+ tpbsw = 0.0025
+ cjswd = 5.3856e-11
+ cjsws = 5.3856e-11
+ rbdb = 50
+ pua1 = -9.6760461e-23
+ prwb = 0
+ pub1 = 5.7312604e-33
+ prwg = 0
+ puc1 = -1.747778e-23
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ nigbinv = 2.171
+ pute = -4.8084303e-14
+ rdsw = 200
+ toxref = 3e-9
+ )

.model pch_fs_28 pmos (
+ level = 54
+ wtvfbsdoff = 0
+ lku0we = 1.8e-11
+ k2we = 5e-5
+ epsrox = 3.9
+ dsub = 0.5
+ dtox = 3.91e-10
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ ltvfbsdoff = 0
+ bigbacc = 0.0054401
+ rdsmod = 0
+ igbmod = 1
+ wkvth0we = 0.0
+ eta0 = 0.17962267
+ etab = -0.19577778
+ kvth0we = -0.00022
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ trnqsmod = 0
+ pbswgd = 0.8
+ lintnoi = -5e-9
+ pbswgs = 0.8
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ pvoff = -2.0654209e-16
+ igcmod = 1
+ cdscb = 0
+ cdscd = 0
+ pvsat = 0
+ wk2we = 0.0
+ pvth0 = -8.1676914e-16
+ ptvfbsdoff = 0
+ drout = 0.56
+ paigc = -3.9499473e-18
+ voffl = 0
+ rgatemod = 0
+ tnjtsswg = 1
+ weta0 = -1.7872176e-8
+ wetab = 1.9534667e-8
+ lpclm = 0
+ cgidl = 1
+ permod = 1
+ ags = -1.2539967
+ nfactor = 1
+ cjd = 0.001421376
+ cit = -0.00036538451
+ cjs = 0.001421376
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 1.38228675e-8
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ pbswd = 0.9
+ pbsws = 0.9
+ voffcv = -0.125
+ wpemod = 1
+ la0 = -4.7253353e-7
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0.00064
+ kt1 = -0.16257215
+ kt2 = -0.066291072
+ lk2 = 1.24447077e-9
+ llc = -1.18e-13
+ lln = 0.7
+ lu0 = -5.437045400000001e-10
+ keta = -0.0061234738
+ mjd = 0.335
+ mjs = 0.335
+ lua = -1.0290148e-16
+ lub = -5.3060964e-27
+ luc = -4.0794824e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pdits = 0
+ pa0 = 9.7298482e-15
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ cigsd = 0.013281
+ pk2 = -2.0891363e-16
+ nigbacc = 10
+ lags = 1.5101544e-6
+ pu0 = 1.1540053e-17
+ dvt0w = 0
+ dvt1w = 0
+ prt = 0
+ dvt2w = 0
+ pua = -1.3867635e-23
+ pub = 2.1855871e-32
+ puc = -2.7646346e-24
+ pud = 0
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 2.2076918e-10
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 1.7313241e-9
+ ub1 = -1.3316629e-18
+ uc1 = 2.2670111e-10
+ kt1l = 0
+ tpb = 0.0016
+ wa0 = -1.7096745e-7
+ ute = -0.86054925
+ web = 6628.3
+ wec = -16935.0
+ pk2we = 0.0
+ wk2 = 4.238936e-9
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ wlc = 0
+ wln = 1
+ wu0 = -2.6120153e-10
+ xgl = -8.2e-9
+ xgw = 0
+ wua = -2.3821198e-16
+ wub = 1.6333936e-25
+ wuc = 4.2583136e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ nigbinv = 2.171
+ lint = 9.7879675e-9
+ tpbswg = 0.001
+ lkt1 = -2.4755192e-8
+ lkt2 = -5.6848171e-9
+ lmax = 4.4908e-7
+ tnoia = 0
+ lmin = 2.1577e-7
+ lpe0 = 6.44e-8
+ ijthsfwd = 0.01
+ lpeb = 0
+ peta0 = -1.6e-17
+ wketa = -7.8373297e-10
+ minv = -0.33
+ tpbsw = 0.0025
+ lua1 = 4.723388e-17
+ lub1 = -3.0366637e-25
+ luc1 = 1.2420632e-17
+ ptvoff = 5.0195791e-17
+ cjswd = 5.3856e-11
+ cjsws = 5.3856e-11
+ ndep = 1e+18
+ fnoimod = 1
+ mjswd = 0.01
+ lute = -2.9424109e-8
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ waigsd = 1.9297907e-12
+ lwlc = 0
+ eigbinv = 1.1
+ moin = 5.5538
+ ijthsrev = 0.01
+ nigc = 2.291
+ diomod = 1
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.9113600000000002e-10
+ pku0we = 0.0
+ cjswgs = 1.9113600000000002e-10
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ tvfbsdoff = 0.1
+ pags = -3.3771496e-13
+ scref = 1e-6
+ a0 = 3.1132665
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 72000
+ cf = 8.17e-11
+ ntox = 1.0
+ mjswgd = 0.95
+ ef = 1.15
+ mjswgs = 0.95
+ k1 = 0.30425
+ k2 = -0.0081283305
+ k3 = -2.5823
+ pcit = -1.00716403e-17
+ em = 20000000.0
+ ppdiblc2 = -3.8737293e-16
+ pclm = 1.1689658
+ pigcd = 2.572
+ cigbacc = 0.245
+ ll = -1.18e-13
+ aigsd = 0.0063633912
+ lw = 0
+ u0 = 0.01164123
+ w0 = 0
+ ua = 3.3584387e-10
+ ub = 1.2266958e-18
+ uc = -5.8379738e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 3.4e-9
+ tcjswg = 0.00128
+ lvoff = -4.2658924e-9
+ phin = 0.15
+ tnoimod = 0
+ lvsat = 8.000000000000001e-6
+ pkt1 = 6.7955166e-15
+ pkt2 = 2.2627554e-16
+ lvth0 = 4.3253579e-9
+ cigbinv = 0.006
+ delta = 0.018814
+ laigc = -1.8017042e-11
+ wvfbsdoff = 0
+ rnoia = 0
+ rnoib = 0
+ lvfbsdoff = 0
+ rbdb = 50
+ pua1 = -2.7108228e-23
+ pkvth0we = 0.0
+ prwb = 0
+ pub1 = 7.1177686e-32
+ prwg = 0
+ puc1 = 8.7727027e-25
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ pketa = 2.0432143e-15
+ version = 4.5
+ ngate = 1.7e+20
+ pute = 1.6065563e-14
+ fprout = 200
+ rdsw = 200
+ ngcon = 1
+ tempmod = 0
+ wpclm = -1.1447315e-8
+ xrcrg1 = 12
+ xrcrg2 = 1
+ vfbsdoff = 0.01
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ aigbacc = 0.012071
+ wtvoff = -1.7507555e-10
+ paramchk = 1
+ rshg = 14.1
+ capmod = 2
+ aigbinv = 0.009974
+ wku0we = 1.5e-11
+ mobmod = 0
+ ijthdfwd = 0.01
+ tvoff = 0.002323434
+ tnom = 25
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ poxedge = 1
+ ijthdrev = 0.01
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = -4.8e-10
+ lpdiblc2 = 4.7505822e-10
+ binunit = 2
+ ppclm = 0
+ wags = 5.6744004e-7
+ wcit = 2.107191e-11
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ voff = -0.12137687
+ acde = 0.5
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ vsat = 91103.982
+ wint = 0
+ vth0 = -0.42406475000000005
+ wkt1 = -2.4180539e-8
+ wkt2 = 4.7880041e-9
+ wmax = 5.426e-7
+ dmcgt = 0
+ aigc = 0.0067599617
+ wmin = 2.726e-7
+ tcjsw = 9.34e-5
+ lkvth0we = 3e-12
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ wua1 = 1.9431072e-17
+ wub1 = -1.3369336e-25
+ wuc1 = -7.3645279e-17
+ acnqsmod = 0
+ bigc = 0.0012521
+ bigsd = 0.0003327
+ wute = -7.6140111e-8
+ wwlc = 0
+ wvoff = 1.674468e-9
+ toxref = 3e-9
+ rbodymod = 0
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ wvsat = 0.0034765009
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ wvth0 = -1.9714099000000003e-9
+ cigc = 0.15259
+ waigc = 1.7749876e-11
+ njtsswg = 6.489
+ lketa = -2.19178e-8
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ ltvoff = -2.3990075e-10
+ xpart = 1
+ ckappad = 0.6
+ wpdiblc2 = 1.1524564e-9
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.0090247504
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ pdiblcb = 0
+ egidl = 0.001
+ pvfbsdoff = 0
+ )

.model pch_fs_29 pmos (
+ level = 54
+ ijthdrev = 0.01
+ ngcon = 1
+ pbswgd = 0.8
+ pbswgs = 0.8
+ wpclm = -1.2079184e-7
+ aigbinv = 0.009974
+ nigc = 2.291
+ igcmod = 1
+ lpdiblc2 = -1.1954251e-9
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ ntox = 1.0
+ pcit = -8.9298391e-18
+ pclm = 1.5407845
+ poxedge = 1
+ phin = 0.15
+ lkvth0we = 3e-12
+ pkt1 = -1.2548200000000001e-15
+ pkt2 = -1.4992738e-15
+ binunit = 2
+ permod = 1
+ tvoff = 0.00085372815
+ acnqsmod = 0
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ rbdb = 50
+ pua1 = 1.9617826e-23
+ prwb = 0
+ pub1 = -3.1346313e-32
+ prwg = 0
+ puc1 = 1.1713402e-23
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ rbodymod = 0
+ voffcv = -0.125
+ wpemod = 1
+ rdsw = 200
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = -4.8e-10
+ ppclm = 2.3071337e-14
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ rshg = 14.1
+ wpdiblc2 = -7.3926191e-10
+ tpbswg = 0.001
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ njtsswg = 6.489
+ ptvoff = -3.132788e-17
+ tnom = 25
+ bigsd = 0.0003327
+ waigsd = 1.9297907e-12
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ wkvth0we = 0.0
+ wvoff = 3.1859801e-10
+ diomod = 1
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.016941733
+ trnqsmod = 0
+ pdiblcb = 0
+ wvsat = 0.0032472346
+ pditsd = 0
+ wvth0 = -7.1269425e-9
+ pditsl = 0
+ cjswgd = 1.9113600000000002e-10
+ pku0we = 0.0
+ cjswgs = 1.9113600000000002e-10
+ waigc = -1.7260908e-11
+ wags = -1.0331048e-6
+ wcit = 1.566053e-11
+ lketa = 7.1935383e-9
+ voff = -0.13201276
+ mjswgd = 0.95
+ mjswgs = 0.95
+ bigbacc = 0.0054401
+ acde = 0.5
+ xpart = 1
+ rgatemod = 0
+ tcjswg = 0.00128
+ vsat = 91523.884
+ wint = 0
+ tnjtsswg = 1
+ vth0 = -0.42162236000000003
+ pvfbsdoff = 0
+ kvth0we = -0.00022
+ egidl = 0.001
+ wkt1 = 1.3972715e-8
+ wkt2 = 1.2965963e-8
+ wmax = 5.426e-7
+ aigc = 0.0067957378
+ wmin = 2.726e-7
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ wua1 = -2.0201942e-16
+ wub1 = 3.5220237e-25
+ wuc1 = -1.2500135e-16
+ bigc = 0.0012521
+ wwlc = 0
+ fprout = 200
+ cdsc = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ a0 = 1.1444157
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ at = 108550.2
+ xtid = 3
+ cf = 8.17e-11
+ xtis = 3
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.025395241
+ k3 = -2.5823
+ em = 20000000.0
+ ll = -1.18e-13
+ lw = 0
+ u0 = 0.0100017592
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ w0 = 0
+ ua = -3.1599722e-11
+ ub = 1.4008434e-18
+ uc = -1.6299488e-10
+ ud = 0
+ cigc = 0.15259
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 3.4e-9
+ pvoff = 7.954647100000001e-17
+ wtvoff = 2.1129256e-10
+ cdscb = 0
+ cdscd = 0
+ pvsat = 4.83709e-11
+ wk2we = 0.0
+ pvth0 = 2.7104823999999996e-16
+ drout = 0.56
+ paigc = 3.4373281e-18
+ nfactor = 1
+ capmod = 2
+ voffl = 0
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ wku0we = 1.5e-11
+ dmdg = 0
+ weta0 = -1.7872176e-8
+ wetab = 1.9534667e-8
+ mobmod = 0
+ ags = 5.9031333
+ lpclm = -7.8453093e-8
+ cjd = 0.001421376
+ cit = 0.00015305446
+ cjs = 0.001421376
+ clc = 1e-7
+ cle = 0.6
+ k2we = 5e-5
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 1.38228675e-8
+ ijthsfwd = 0.01
+ k3b = 2.1176
+ dsub = 0.5
+ cgidl = 1
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ dtox = 3.91e-10
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ nigbacc = 10
+ la0 = -5.7105222e-8
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = -0.0070720921
+ kt1 = -0.27233533
+ kt2 = -0.10755274
+ lk2 = 4.887788899999999e-9
+ eta0 = 0.17962267
+ llc = -1.18e-13
+ lln = 0.7
+ lu0 = -1.9777630000000002e-10
+ etab = -0.19577778
+ mjd = 0.335
+ mjs = 0.335
+ lua = -2.5370884e-17
+ lub = -4.2051244e-26
+ luc = 1.7994313e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ pbswd = 0.9
+ pbsws = 0.9
+ njd = 1.02
+ njs = 1.02
+ pa0 = -3.159814e-15
+ ijthsrev = 0.01
+ nsd = 1e+20
+ pbd = 0.75
+ pat = -4.5415452e-10
+ pbs = 0.75
+ pk2 = -2.0710507e-16
+ pu0 = 4.0684676e-18
+ prt = 0
+ pua = 6.5898257e-24
+ pub = -4.9701536e-33
+ puc = -7.066739e-24
+ pud = 0
+ nigbinv = 2.171
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 2.8369875e-9
+ ub1 = -4.0389099e-18
+ uc1 = 4.2708978e-10
+ tpb = 0.0016
+ wa0 = -1.0988104e-7
+ pdits = 0
+ ute = -1
+ wat = 0.0021523911
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 4.2303646e-9
+ cigsd = 0.013281
+ wlc = 0
+ wln = 1
+ wu0 = -2.2579117e-10
+ xgl = -8.2e-9
+ xgw = 0
+ wua = -3.3516677e-16
+ dvt0w = 0
+ wub = 2.9047692e-25
+ wuc = 6.2972257e-17
+ wud = 0
+ dvt1w = 0
+ dvt2w = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ ppdiblc2 = 1.1779633e-17
+ pk2we = 0.0
+ fnoimod = 1
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ eigbinv = 1.1
+ tnoia = 0
+ peta0 = -1.6e-17
+ wketa = 1.4826965e-8
+ tpbsw = 0.0025
+ cjswd = 5.3856e-11
+ cjsws = 5.3856e-11
+ pkvth0we = 0.0
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ toxref = 3e-9
+ cigbacc = 0.245
+ vfbsdoff = 0.01
+ tnoimod = 0
+ keta = -0.1440919
+ tvfbsdoff = 0.1
+ wtvfbsdoff = 0
+ cigbinv = 0.006
+ ltvoff = 7.0207177e-11
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 1.1137855999999999e-10
+ paramchk = 1
+ scref = 1e-6
+ kt1l = 0
+ pigcd = 2.572
+ aigsd = 0.0063633912
+ ltvfbsdoff = 0
+ version = 4.5
+ lvoff = -2.0217201e-9
+ lint = 9.7879675e-9
+ tempmod = 0
+ lkt1 = -1.5951622e-9
+ lkt2 = 3.021395e-9
+ lku0we = 1.8e-11
+ lmax = 2.1577e-7
+ lvsat = -8.059139999999999e-5
+ lmin = 9e-8
+ epsrox = 3.9
+ lvth0 = 3.8100147e-9
+ lpe0 = 6.44e-8
+ ijthdfwd = 0.01
+ lpeb = 0
+ delta = 0.018814
+ laigc = -2.5565813e-11
+ aigbacc = 0.012071
+ wvfbsdoff = 0
+ rdsmod = 0
+ lvfbsdoff = 0
+ minv = -0.33
+ rnoia = 0
+ rnoib = 0
+ lua1 = -1.8606111e-16
+ lub1 = 2.6756274e-25
+ luc1 = -2.9861377e-17
+ igbmod = 1
+ ndep = 1e+18
+ ptvfbsdoff = 0
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ lwlc = 0
+ pketa = -1.250643e-15
+ ngate = 1.7e+20
+ moin = 5.5538
+ )

.model pch_fs_30 pmos (
+ level = 54
+ ijthdrev = 0.01
+ ngcon = 1
+ pbswgd = 0.8
+ pbswgs = 0.8
+ wpclm = 4.9341412e-7
+ aigbinv = 0.009974
+ nigc = 2.291
+ igcmod = 1
+ lpdiblc2 = 0
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ ntox = 1.0
+ pcit = -6.978865e-18
+ pclm = 0.08631615
+ paigsd = 8.4526218e-25
+ poxedge = 1
+ phin = 0.15
+ lkvth0we = 3e-12
+ pkt1 = -1.7524191000000001e-15
+ pkt2 = 2.1480498e-17
+ binunit = 2
+ permod = 1
+ tvoff = 0.0012365685
+ acnqsmod = 0
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ rbdb = 50
+ pua1 = 4.1792962e-25
+ prwb = 0
+ pub1 = 6.1746384e-33
+ prwg = 0
+ puc1 = 2.9246063e-24
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ rbodymod = 0
+ voffcv = -0.125
+ wpemod = 1
+ rdsw = 200
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = -9.0458832e-9
+ letab = 1.7579973e-8
+ ppclm = -3.4664022e-14
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ rshg = 14.1
+ wpdiblc2 = -6.1394667e-10
+ tpbswg = 0.001
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ njtsswg = 6.489
+ ptvoff = 2.0376593e-17
+ tnom = 25
+ bigsd = 0.0003327
+ waigsd = 1.9297817e-12
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ wkvth0we = 0.0
+ wvoff = -2.8254962e-9
+ diomod = 1
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.0042244444
+ trnqsmod = 0
+ pdiblcb = 0
+ wvsat = 0.017016245
+ pditsd = 0
+ wvth0 = -5.9631861e-9
+ pditsl = 0
+ cjswgd = 1.9113600000000002e-10
+ pku0we = 0.0
+ cjswgs = 1.9113600000000002e-10
+ waigc = 7.1461687e-12
+ wags = -1.0331048e-6
+ wcit = -5.09452e-12
+ lketa = -1.1878561e-8
+ voff = -0.12098873
+ mjswgd = 0.95
+ mjswgs = 0.95
+ bigbacc = 0.0054401
+ acde = 0.5
+ xpart = 1
+ rgatemod = 0
+ tcjswg = 0.00128
+ vsat = 62231.739
+ wint = 0
+ tnjtsswg = 1
+ vth0 = -0.36546471
+ pvfbsdoff = 0
+ kvth0we = -0.00022
+ egidl = 0.001
+ wkt1 = 1.9266322e-8
+ wkt2 = -3.2122744e-9
+ wmax = 5.426e-7
+ aigc = 0.0067006504
+ wmin = 2.726e-7
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ wua1 = 2.2347963e-18
+ wub1 = -4.6956688e-26
+ wuc1 = -3.1503526e-17
+ bigc = 0.0012521
+ wwlc = 0
+ fprout = 200
+ cdsc = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ a0 = 3.9744452
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ at = 69068.642
+ xtid = 3
+ cf = 8.17e-11
+ xtis = 3
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.022825095
+ k3 = -2.5823
+ em = 20000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.0041656963000000005
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ w0 = 0
+ ua = -9.2439852e-11
+ ub = -1.6232125e-18
+ uc = 5.3507127e-11
+ ud = 0
+ cigc = 0.15259
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 3.4e-9
+ pvoff = 3.7509131999999996e-16
+ wtvoff = -3.3875503e-10
+ cdscb = 0
+ cdscd = 0
+ pvsat = -1.2459161e-9
+ wk2we = 0.0
+ pvth0 = 1.6165514e-16
+ drout = 0.56
+ paigc = 1.1430629e-18
+ nfactor = 1
+ capmod = 2
+ voffl = 0
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ wku0we = 1.5e-11
+ dmdg = 0
+ weta0 = -5.5239839e-8
+ wetab = 4.6876459e-8
+ mobmod = 0
+ ags = 5.9031333
+ lpclm = 5.8266931e-8
+ cjd = 0.001421376
+ cit = -0.00018033605
+ cjs = 0.001421376
+ clc = 1e-7
+ cle = 0.6
+ k2we = 5e-5
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 4.0349e-9
+ ijthsfwd = 0.01
+ k3b = 2.1176
+ dsub = 0.5
+ cgidl = 1
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ dtox = 3.91e-10
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ nigbacc = 10
+ la0 = -3.23128e-7
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = -0.0033608257000000002
+ kt1 = -0.32608492
+ kt2 = -0.08284588
+ lk2 = 4.6461952e-9
+ eta0 = 0.27074908
+ llc = 0
+ lln = 1
+ lu0 = 3.5081362e-10
+ etab = -0.38279877
+ mjd = 0.335
+ mjs = 0.335
+ lua = -1.9651912e-17
+ lub = 2.4221001e-25
+ luc = -2.356876e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ pbswd = 0.9
+ pbsws = 0.9
+ njd = 1.02
+ njs = 1.02
+ pa0 = 9.1746422e-14
+ laigsd = -3.0625433e-18
+ ijthsrev = 0.01
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 6.7620954e-11
+ pbs = 0.75
+ pk2 = 2.5170462e-16
+ pu0 = -8.2666616e-17
+ prt = 0
+ pua = 3.032424e-23
+ pub = -9.6166295e-32
+ puc = -2.0363205e-24
+ pud = 0
+ nigbinv = 2.171
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = -2.7998083e-10
+ ub1 = 8.7083504e-19
+ uc1 = 1.8820988e-11
+ tpb = 0.0016
+ wa0 = -1.1195219e-6
+ pdits = 0
+ ute = -1
+ wat = -0.0033984119
+ web = 6628.3
+ wec = -16935.0
+ wk2 = -6.5058945e-10
+ cigsd = 0.013281
+ wlc = 0
+ wln = 1
+ wu0 = 6.9692249e-10
+ xgl = -8.2e-9
+ xgw = 0
+ wua = -5.8766054e-16
+ dvt0w = 0
+ wub = 1.2606486e-24
+ wuc = 9.4571662e-18
+ wud = 0
+ dvt1w = 0
+ dvt2w = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ ppdiblc2 = 0
+ pk2we = 0.0
+ fnoimod = 1
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ eigbinv = 1.1
+ tnoia = 0
+ peta0 = 3.4965603e-15
+ petab = -2.5701285e-15
+ wketa = -3.6489897e-8
+ tpbsw = 0.0025
+ cjswd = 5.3856e-11
+ cjsws = 5.3856e-11
+ pkvth0we = 0.0
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ toxref = 3e-9
+ cigbacc = 0.245
+ vfbsdoff = 0.01
+ tnoimod = 0
+ keta = 0.058802768
+ tvfbsdoff = 0.1
+ wtvfbsdoff = 0
+ cigbinv = 0.006
+ ltvoff = 3.4220189e-11
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 1.4271727e-10
+ paramchk = 1
+ scref = 1e-6
+ kt1l = 0
+ pigcd = 2.572
+ aigsd = 0.0063633912
+ ltvfbsdoff = 0
+ version = 4.5
+ lvoff = -3.0579783e-9
+ lint = 0
+ tempmod = 0
+ lkt1 = 3.4572998999999996e-9
+ lkt2 = 6.989501e-10
+ lku0we = 1.8e-11
+ lmax = 9e-8
+ lvsat = 0.0026728703
+ lmin = 5.4e-8
+ epsrox = 3.9
+ lvth0 = -1.4688048e-9
+ lpe0 = 6.44e-8
+ ijthdfwd = 0.01
+ lpeb = 0
+ delta = 0.018814
+ laigc = -1.6627591e-11
+ aigbacc = 0.012071
+ wvfbsdoff = 0
+ rdsmod = 0
+ lvfbsdoff = 0
+ minv = -0.33
+ rnoia = 0
+ rnoib = 0
+ lua1 = 1.0693391e-16
+ lub1 = -1.9395329e-25
+ luc1 = 8.5158894e-18
+ igbmod = 1
+ ndep = 1e+18
+ ptvfbsdoff = 0
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ lwlc = 0
+ pketa = 3.573142e-15
+ ngate = 1.7e+20
+ moin = 5.5538
+ )

.model pch_fs_31 pmos (
+ level = 54
+ paigc = -3.8652128e-18
+ voff = -0.11425646
+ nigbacc = 10
+ ags = 5.9031333
+ acde = 0.5
+ ppdiblc2 = 0
+ voffl = 0
+ cjd = 0.001421376
+ cit = -0.0023632098
+ cjs = 0.001421376
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ vsat = 205509.49
+ dlc = 4.0349e-9
+ wint = 0
+ k3b = 2.1176
+ vth0 = -0.34541972000000004
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ weta0 = 4.5345198e-8
+ wkt1 = -9.053012e-8
+ wkt2 = -4.5663135e-8
+ wetab = 2.1214781e-8
+ wmax = 5.426e-7
+ aigc = 0.0065523001
+ wmin = 2.726e-7
+ lpclm = -1.6067206e-7
+ permod = 1
+ nigbinv = 2.171
+ la0 = 2.2449695e-9
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = -0.0003052786699999999
+ kt1 = -0.078489325
+ kt2 = 0.051187672
+ lk2 = 5.7431101e-9
+ llc = 0
+ lln = 1
+ cgidl = 1
+ lu0 = -6.4229203e-10
+ mjd = 0.335
+ mjs = 0.335
+ lua = -5.2618623e-17
+ lub = -3.080728e-25
+ luc = -2.0280652e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ wua1 = 2.8402308e-15
+ njs = 1.02
+ wub1 = -3.9062366e-24
+ wuc1 = 2.0276364e-16
+ pa0 = -4.432942e-14
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 1.8264736e-9
+ pbs = 0.75
+ pk2 = -1.1995676e-16
+ pu0 = 2.2577126e-16
+ bigc = 0.0012521
+ prt = 0
+ pua = 1.5923531e-23
+ pub = 9.2000466e-32
+ puc = 3.3504384e-24
+ pud = 0
+ wwlc = 0
+ pkvth0we = 0.0
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = -3.345352e-9
+ ub1 = 3.9080279e-18
+ uc1 = 1.4308247e-10
+ tpb = 0.0016
+ voffcv = -0.125
+ wpemod = 1
+ pbswd = 0.9
+ pbsws = 0.9
+ wa0 = 1.2266134e-6
+ cdsc = 0
+ ute = -1
+ wat = -0.033723458
+ web = 6628.3
+ wec = -16935.0
+ fnoimod = 1
+ wk2 = 5.7573654e-9
+ wlc = 0
+ cgbo = 0
+ wln = 1
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ wu0 = -4.6209719e-9
+ xtid = 3
+ xgl = -8.2e-9
+ xtis = 3
+ xgw = 0
+ wua = -3.3937245e-16
+ wub = -1.9836059e-24
+ wuc = -8.3417988e-17
+ wud = 0
+ eigbinv = 1.1
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ vfbsdoff = 0.01
+ cigc = 0.15259
+ pdits = 0
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ paramchk = 1
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ tpbswg = 0.001
+ cigbacc = 0.245
+ tnoia = 0
+ k2we = 5e-5
+ tnoimod = 0
+ ijthdfwd = 0.01
+ peta0 = -2.3373718e-15
+ dsub = 0.5
+ petab = -1.0817512e-15
+ dtox = 3.91e-10
+ wketa = 7.0696889e-8
+ ptvoff = -1.3332507e-17
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ tpbsw = 0.0025
+ waigsd = 1.9297962e-12
+ cigbinv = 0.006
+ cjswd = 5.3856e-11
+ cjsws = 5.3856e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ eta0 = 0.012687945
+ etab = -0.23454709
+ diomod = 1
+ ijthdrev = 0.01
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.9113600000000002e-10
+ pku0we = 0.0
+ version = 4.5
+ cjswgs = 1.9113600000000002e-10
+ lpdiblc2 = 0
+ tempmod = 0
+ tvfbsdoff = 0.1
+ aigbacc = 0.012071
+ mjswgd = 0.95
+ mjswgs = 0.95
+ scref = 1e-6
+ tcjswg = 0.00128
+ pigcd = 2.572
+ aigsd = 0.0063633912
+ lvoff = -3.4484499e-9
+ lkvth0we = 3e-12
+ aigbinv = 0.009974
+ lvsat = -0.0056372393
+ lvth0 = -2.6314143e-9
+ delta = 0.018814
+ wvfbsdoff = 0
+ laigc = -8.0232722e-12
+ lvfbsdoff = 0
+ rnoia = 0
+ rnoib = 0
+ acnqsmod = 0
+ fprout = 200
+ pketa = -2.6436916e-15
+ ngate = 1.7e+20
+ xrcrg1 = 12
+ xrcrg2 = 1
+ rbodymod = 0
+ ngcon = 1
+ wpclm = -6.9641486e-7
+ poxedge = 1
+ gbmin = 1e-12
+ wtvoff = 2.4243635e-10
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ keta = -0.44725926
+ binunit = 2
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 2.6932394999999997e-10
+ capmod = 2
+ kt1l = 0
+ wku0we = 1.5e-11
+ wpdiblc2 = -6.1394667e-10
+ mobmod = 0
+ lint = 0
+ lkt1 = -1.0903245e-8
+ lkt2 = -7.0749959e-9
+ lmax = 5.4e-8
+ lmin = 4.5e-8
+ a0 = -1.6354335
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 16386.797
+ cf = 8.17e-11
+ lpe0 = 6.44e-8
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.041737421
+ k3 = -2.5823
+ em = 20000000.0
+ lpeb = 0
+ ll = 0
+ lw = 0
+ u0 = 0.021288207
+ w0 = 0
+ tvoff = 0.0019328761
+ ua = 4.7595173e-10
+ ub = 7.8644222e-18
+ uc = 4.7837975e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 3.4e-9
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ minv = -0.33
+ xjbvd = 1
+ xjbvs = 1
+ lua1 = 2.8472544e-16
+ lub1 = -3.7011047e-25
+ lk2we = 0.0
+ luc1 = 1.3087235e-18
+ ndep = 1e+18
+ wkvth0we = 0.0
+ lwlc = 0
+ moin = 5.5538
+ ku0we = -0.0007
+ trnqsmod = 0
+ nigc = 2.291
+ beta0 = 13.32
+ leta0 = 5.9216629e-9
+ letab = 8.9813755e-9
+ ppclm = 3.4346058e-14
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ njtsswg = 6.489
+ ntox = 1.0
+ pcit = -1.8424609999999998e-17
+ pclm = 3.8611263
+ rgatemod = 0
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ tnjtsswg = 1
+ dmcgt = 0
+ ckappad = 0.6
+ phin = 0.15
+ ckappas = 0.6
+ tcjsw = 9.34e-5
+ pdiblc1 = 0
+ pdiblc2 = 0.0042244444
+ pdiblcb = 0
+ pkt1 = 4.6157745000000004e-15
+ pkt2 = 2.4836304e-15
+ bigsd = 0.0003327
+ toxref = 3e-9
+ rbdb = 50
+ pua1 = -1.6418584e-22
+ prwb = 0
+ pub1 = 2.3001287e-31
+ prwg = 0
+ puc1 = -1.0662889e-23
+ wtvfbsdoff = 0
+ bigbacc = 0.0054401
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ wvoff = 3.9335999e-9
+ rdsw = 200
+ wvsat = -0.031328619
+ kvth0we = -0.00022
+ ltvfbsdoff = 0
+ wvth0 = 8.982980999999999e-9
+ waigc = 9.3495749e-11
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ ltvoff = -6.1656569e-12
+ lketa = 1.7473037e-8
+ xpart = 1
+ rshg = 14.1
+ pvfbsdoff = 0
+ egidl = 0.001
+ ptvfbsdoff = 0
+ lku0we = 1.8e-11
+ epsrox = 3.9
+ ijthsfwd = 0.01
+ rdsmod = 0
+ igbmod = 1
+ tnom = 25
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ nfactor = 1
+ pbswgd = 0.8
+ pbswgs = 0.8
+ ijthsrev = 0.01
+ igcmod = 1
+ pvoff = -1.6936247999999996e-17
+ cdscb = 0
+ cdscd = 0
+ wags = -1.0331048e-6
+ pvsat = 1.5580861e-9
+ wk2we = 0.0
+ pvth0 = -7.0522254e-16
+ wcit = 1.9224593e-10
+ drout = 0.56
+ )

.model pch_fs_32 pmos (
+ level = 54
+ tvoff = 0.0050068134
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ voffcv = -0.125
+ wpemod = 1
+ njtsswg = 6.489
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = 2.2314638e-9
+ ckappad = 0.6
+ letab = 1.8240871e-9
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.0042244444
+ pdiblcb = 0
+ keta = -0.10111506
+ ppclm = 1.7398739e-15
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 1.11605e-11
+ kt1l = 0
+ tpbswg = 0.001
+ bigbacc = 0.0054401
+ lint = 0
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ lkt1 = -1.3889032e-8
+ lkt2 = 2.2261728e-10
+ lmax = 4.5e-8
+ kvth0we = -0.00022
+ lmin = 3.6e-8
+ lpe0 = 6.44e-8
+ ijthsfwd = 0.01
+ lpeb = 0
+ ptvoff = 3.2244316e-17
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ waigsd = 1.9257033e-12
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ minv = -0.33
+ bigsd = 0.0003327
+ lua1 = -1.7116539e-16
+ lub1 = 1.8549471e-25
+ luc1 = 2.2025561e-17
+ ndep = 1e+18
+ diomod = 1
+ lwlc = 0
+ wvoff = 1.094003e-8
+ moin = 5.5538
+ ijthsrev = 0.01
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.9113600000000002e-10
+ pku0we = 0.0
+ cjswgs = 1.9113600000000002e-10
+ nigc = 2.291
+ wvsat = -0.018712604
+ wvth0 = 1.3422333e-8
+ waigc = 1.753535e-10
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ mjswgd = 0.95
+ mjswgs = 0.95
+ lketa = 5.1197136e-10
+ tcjswg = 0.00128
+ xpart = 1
+ ntox = 1.0
+ ppdiblc2 = 0
+ pcit = 1.2074904e-16
+ pclm = 0.85281474
+ pvfbsdoff = 0
+ nfactor = 1
+ egidl = 0.001
+ phin = 0.15
+ pkt1 = 2.398466e-15
+ pkt2 = -1.2154904e-16
+ fprout = 200
+ pkvth0we = 0.0
+ rbdb = 50
+ pua1 = 5.9435365e-23
+ prwb = 0
+ pub1 = -6.8901825e-32
+ prwg = 0
+ puc1 = -3.4884574e-24
+ xrcrg1 = 12
+ xrcrg2 = 1
+ nigbacc = 10
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ rdsw = 200
+ wtvoff = -6.8770288e-10
+ vfbsdoff = 0.01
+ pvoff = -3.6025133000000004e-16
+ ags = 5.9031333
+ nigbinv = 2.171
+ cdscb = 0
+ cdscd = 0
+ cjd = 0.001421376
+ cit = 0.0029054321
+ cjs = 0.001421376
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ pvsat = 9.3990127e-10
+ dlc = 4.0349e-9
+ wk2we = 0.0
+ pvth0 = -9.227508000000001e-16
+ k3b = 2.1176
+ dwb = 0
+ drout = 0.56
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ capmod = 2
+ paramchk = 1
+ paigc = -7.8762427e-18
+ wku0we = 1.5e-11
+ rshg = 14.1
+ voffl = 0
+ la0 = -2.1218621e-7
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0.011148083
+ mobmod = 0
+ kt1 = -0.017554887
+ kt2 = -0.09774321
+ lk2 = 4.3772258e-9
+ llc = 0
+ lln = 1
+ lu0 = -2.443917e-10
+ mjd = 0.335
+ mjs = 0.335
+ lua = 4.1444844e-17
+ lub = -1.5666965e-25
+ luc = -1.4956542e-17
+ lud = 0
+ lwc = 0
+ weta0 = 6.5061382e-9
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ wetab = -5.613608e-9
+ njs = 1.02
+ pa0 = 5.0455005e-14
+ fnoimod = 1
+ nsd = 1e+20
+ pbd = 0.75
+ pat = -2.4847929e-9
+ pbs = 0.75
+ pk2 = 3.3742201e-16
+ lpclm = -1.3264792e-8
+ pu0 = 1.5059926e-16
+ eigbinv = 1.1
+ prt = 0
+ pua = 9.2877876e-24
+ pub = 3.2782262e-32
+ puc = 3.1614905e-24
+ pud = 0
+ ijthdfwd = 0.01
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 5.9585425e-9
+ ub1 = -7.4308533e-18
+ uc1 = -2.7971012e-10
+ cgidl = 1
+ tpb = 0.0016
+ wa0 = -7.0776268e-7
+ ute = -1
+ wat = 0.054261574
+ web = 6628.3
+ wec = -16935.0
+ wk2 = -3.5768953e-9
+ wlc = 0
+ wln = 1
+ wu0 = -3.0868494e-9
+ tnom = 25
+ xgl = -8.2e-9
+ xgw = 0
+ wua = -2.0394912e-16
+ wub = -7.7507108e-25
+ wuc = -7.9561907e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ laigsd = -3.6731852e-16
+ pbswd = 0.9
+ pbsws = 0.9
+ ijthdrev = 0.01
+ cigbacc = 0.245
+ lpdiblc2 = 0
+ pdits = 0
+ wags = -1.0331048e-6
+ cigsd = 0.013281
+ tnoimod = 0
+ dvt0w = 0
+ dvt1w = 0
+ wcit = -2.6480326e-9
+ dvt2w = 0
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ a0 = 2.7407131
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = -217355.29
+ cf = 8.17e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.013862232
+ k3 = -2.5823
+ em = 20000000.0
+ voff = -0.14966725
+ ll = 0
+ lw = 0
+ u0 = 0.013167793
+ w0 = 0
+ cigbinv = 0.006
+ acde = 0.5
+ ua = -1.4437109e-9
+ ub = 4.7745619e-18
+ uc = 3.1168444e-10
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 3.4e-9
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ vsat = 182315.32
+ wint = 0
+ vth0 = -0.41707143
+ wkt1 = -4.5278925e-8
+ wkt2 = 7.5037926e-9
+ wtvfbsdoff = 0
+ wmax = 5.426e-7
+ aigc = 0.006152944
+ wmin = 2.726e-7
+ lkvth0we = 3e-12
+ tnoia = 0
+ version = 4.5
+ tempmod = 0
+ peta0 = -4.3425789e-16
+ ltvfbsdoff = 0
+ petab = 2.3283989e-16
+ wketa = 1.3494424e-8
+ wua1 = -1.7234672e-15
+ wub1 = 2.1940634e-24
+ wuc1 = 5.6346661e-17
+ tpbsw = 0.0025
+ acnqsmod = 0
+ toxref = 3e-9
+ bigc = 0.0012521
+ aigbacc = 0.012071
+ cjswd = 5.3856e-11
+ cjsws = 5.3856e-11
+ wwlc = 0
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ rbodymod = 0
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigc = 0.15259
+ aigbinv = 0.009974
+ tvfbsdoff = 0.1
+ ptvfbsdoff = 0
+ ltvoff = -1.5678858e-10
+ scref = 1e-6
+ pigcd = 2.572
+ aigsd = 0.0063633987
+ wpdiblc2 = -6.1394667e-10
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ lku0we = 1.8e-11
+ lvoff = -1.7133213e-9
+ epsrox = 3.9
+ lvsat = -0.0045007251
+ poxedge = 1
+ lvth0 = 8.795196e-10
+ k2we = 5e-5
+ wvfbsdoff = 0
+ rdsmod = 0
+ lvfbsdoff = 0
+ delta = 0.018814
+ dsub = 0.5
+ dtox = 3.91e-10
+ laigc = 1.1545174e-11
+ igbmod = 1
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ binunit = 2
+ rnoia = 0
+ rnoib = 0
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ pbswgd = 0.8
+ wkvth0we = 0.0
+ pbswgs = 0.8
+ eta0 = 0.08799813
+ pketa = 1.5922924e-16
+ etab = -0.088479977
+ ngate = 1.7e+20
+ ngcon = 1
+ igcmod = 1
+ wpclm = -3.0982532e-8
+ trnqsmod = 0
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ paigsd = 2.0055591e-22
+ rgatemod = 0
+ tnjtsswg = 1
+ permod = 1
+ )

.model pch_fs_33 pmos (
+ level = 54
+ version = 4.5
+ pdits = 0
+ cigsd = 0.013281
+ tempmod = 0
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ tpbswg = 0.001
+ rshg = 14.1
+ aigbacc = 0.012071
+ wpdiblc2 = 3.3638075e-10
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ tnoia = 0
+ ptvoff = 0
+ aigbinv = 0.009974
+ peta0 = -1.6e-17
+ waigsd = 1.9846811e-12
+ wketa = -1.9384664e-9
+ tpbsw = 0.0025
+ tnom = 25
+ diomod = 1
+ cjswd = 5.3856e-11
+ cjsws = 5.3856e-11
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ wkvth0we = 0.0
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.9113600000000002e-10
+ pku0we = 0.0
+ cjswgs = 1.9113600000000002e-10
+ trnqsmod = 0
+ tvfbsdoff = 0.1
+ poxedge = 1
+ mjswgd = 0.95
+ wags = 5.1942014e-9
+ mjswgs = 0.95
+ tcjswg = 0.00128
+ binunit = 2
+ scref = 1e-6
+ voff = -0.10372023
+ acde = 0.5
+ pigcd = 2.572
+ aigsd = 0.0063632583
+ rgatemod = 0
+ vsat = 108525.44
+ tnjtsswg = 1
+ wint = 0
+ vth0 = -0.39687116
+ lvoff = 0
+ wkt1 = -3.0503659e-9
+ wkt2 = -7.2833333e-10
+ wmax = 2.726e-7
+ aigc = 0.0068302204
+ wmin = 1.08e-7
+ lvsat = 8.000000000000001e-6
+ lvth0 = -2.4e-10
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ delta = 0.018814
+ wua1 = -5.5326541e-17
+ wub1 = -1.0689498e-25
+ wuc1 = -1.2119467e-17
+ fprout = 200
+ rnoia = 0
+ rnoib = 0
+ bigc = 0.0012521
+ wute = -7.6523556e-8
+ xrcrg1 = 12
+ xrcrg2 = 1
+ wwlc = 0
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ ngate = 1.7e+20
+ ngcon = 1
+ cdsc = 0
+ wpclm = 7.1298978e-9
+ cgbo = 0
+ cgdl = 3.0105e-11
+ wtvoff = -7.3630015e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigc = 0.15259
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ capmod = 2
+ wku0we = 1.5e-11
+ mobmod = 0
+ njtsswg = 6.489
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ k2we = 5e-5
+ ckappad = 0.6
+ ckappas = 0.6
+ ijthsfwd = 0.01
+ pdiblc1 = 0
+ pdiblc2 = 0.0015492917
+ dsub = 0.5
+ pdiblcb = 0
+ dtox = 3.91e-10
+ tvoff = 0.0025423547
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ eta0 = 0.10792519
+ etab = -0.13555556
+ ijthsrev = 0.01
+ ku0we = -0.0007
+ bigbacc = 0.0054401
+ beta0 = 13.32
+ leta0 = -4.8e-10
+ wtvfbsdoff = 0
+ kvth0we = -0.00022
+ ppclm = 0
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ dlcig = 2.5e-9
+ lintnoi = -5e-9
+ bgidl = 1834800000.0
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ ltvfbsdoff = 0
+ ppdiblc2 = 0
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ toxref = 3e-9
+ bigsd = 0.0003327
+ ptvfbsdoff = 0
+ pkvth0we = 0.0
+ wvoff = 1.4142431e-9
+ a0 = 2.5876667
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 72000
+ cf = 8.17e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.015389268
+ k3 = -2.5823
+ em = 20000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.0096471852
+ w0 = 0
+ ua = -1.9215717e-10
+ ub = 1.2747184e-18
+ uc = -1.7585185e-12
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 3.4e-9
+ wvsat = -0.0013318206
+ nfactor = 1
+ wvth0 = -5.3854372e-9
+ vfbsdoff = 0.01
+ waigc = 1.6569661e-12
+ keta = 0.02482765
+ ltvoff = 0
+ jswd = 3.69e-13
+ lketa = 0
+ jsws = 3.69e-13
+ paramchk = 1
+ lcit = 1.6e-11
+ xpart = 1
+ pvfbsdoff = 0
+ kt1l = 0
+ lku0we = 1.8e-11
+ nigbacc = 10
+ egidl = 0.001
+ epsrox = 3.9
+ lint = 6.5375218e-9
+ lkt1 = -4.8e-10
+ lmax = 2.001e-5
+ lmin = 8.9991e-6
+ rdsmod = 0
+ ijthdfwd = 0.01
+ lpe0 = 6.44e-8
+ igbmod = 1
+ lpeb = 0
+ nigbinv = 2.171
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ minv = -0.33
+ pbswgd = 0.8
+ pbswgs = 0.8
+ ndep = 1e+18
+ ags = 0.89683683
+ lwlc = 0
+ igcmod = 1
+ moin = 5.5538
+ ijthdrev = 0.01
+ cjd = 0.001421376
+ cit = 5e-6
+ cjs = 0.001421376
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 1.0572421799999999e-8
+ nigc = 2.291
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ lpdiblc2 = 0
+ fnoimod = 1
+ pvoff = 2e-17
+ eigbinv = 1.1
+ cdscb = 0
+ cdscd = 0
+ la0 = 0
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ jsd = 1.5e-7
+ pvsat = 0
+ jss = 1.5e-7
+ lat = 0.00064
+ kt1 = -0.17197747
+ lk2 = 3.2000000000000003e-10
+ kt2 = -0.050761111
+ wk2we = 0.0
+ pvth0 = -1.2e-16
+ llc = 0
+ lln = 1
+ lu0 = -8e-13
+ drout = 0.56
+ mjd = 0.335
+ mjs = 0.335
+ lub = 0
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 0
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ pk2 = 0
+ pu0 = 0
+ ntox = 1.0
+ voffl = 0
+ prt = 0
+ pub = 0
+ pcit = -8.000000000000001e-19
+ pud = 0
+ pclm = 1.101657
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 9.8162749e-10
+ ub1 = -3.8648101e-20
+ uc1 = 8.1681111e-11
+ tpb = 0.0016
+ weta0 = 1.9163288999999998e-9
+ permod = 1
+ wa0 = 4.8944e-8
+ wetab = 2.9133333e-9
+ ute = -0.81574074
+ phin = 0.15
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 3.9065138e-9
+ lkvth0we = 3e-12
+ lpclm = 0
+ wlc = 0
+ wln = 1
+ wu0 = 5.8460889e-11
+ xgl = -8.2e-9
+ xgw = 0
+ wua = -4.8614483e-17
+ wub = 8.106039e-27
+ wuc = 3.3309111e-18
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ cigbacc = 0.245
+ pkt1 = -4e-17
+ cgidl = 1
+ tnoimod = 0
+ acnqsmod = 0
+ voffcv = -0.125
+ wpemod = 1
+ rbdb = 50
+ prwb = 0
+ prwg = 0
+ rbpb = 50
+ rbpd = 50
+ cigbinv = 0.006
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ pbswd = 0.9
+ rbodymod = 0
+ pbsws = 0.9
+ rdsw = 200
+ )

.model pch_fs_34 pmos (
+ level = 54
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ nfactor = 1
+ ptvoff = -5.393716e-17
+ k2we = 5e-5
+ waigsd = 1.9861139e-12
+ ijthdfwd = 0.01
+ dsub = 0.5
+ dtox = 3.91e-10
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ diomod = 1
+ bigsd = 0.0003327
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.9113600000000002e-10
+ pku0we = 0.0
+ cjswgs = 1.9113600000000002e-10
+ eta0 = 0.10792519
+ wvoff = 1.3100722e-9
+ etab = -0.13555556
+ ijthdrev = 0.01
+ nigbacc = 10
+ wvsat = -0.0013318206
+ wvth0 = -5.481113100000001e-9
+ lpdiblc2 = 6.2970633e-9
+ waigc = 1.4905459e-12
+ mjswgd = 0.95
+ mjswgs = 0.95
+ tcjswg = 0.00128
+ nigbinv = 2.171
+ lketa = -5.5366519e-8
+ pvfbsdoff = 0
+ xpart = 1
+ egidl = 0.001
+ lkvth0we = 3e-12
+ fnoimod = 1
+ ags = 0.84380759
+ eigbinv = 1.1
+ fprout = 200
+ cjd = 0.001421376
+ cit = 5e-6
+ cjs = 0.001421376
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ acnqsmod = 0
+ dlc = 1.0572421799999999e-8
+ xrcrg1 = 12
+ xrcrg2 = 1
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ rbodymod = 0
+ la0 = -3.9401851e-7
+ wtvoff = -6.7630331e-11
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0.00064
+ kt1 = -0.17107141
+ kt2 = -0.050597496
+ lk2 = 5.8519403e-9
+ llc = 0
+ lln = 1
+ lu0 = 9.9598999e-10
+ mjd = 0.335
+ mjs = 0.335
+ lua = -7.2048384e-17
+ lub = 4.3514377e-25
+ luc = 1.4270275e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = -3.1655381e-14
+ pvoff = 9.5649624e-16
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ pk2 = 9.285497e-17
+ keta = 0.030986328
+ pu0 = 3.0504276e-17
+ prt = 0
+ cdscb = 0
+ cdscd = 0
+ pua = 2.7735079e-23
+ pub = -4.2717478e-32
+ puc = 1.20866e-25
+ pud = 0
+ cigbacc = 0.245
+ capmod = 2
+ pvsat = 0
+ rsh = 15.2
+ wk2we = 0.0
+ tcj = 0.000832
+ ua1 = 8.0734953e-10
+ pvth0 = 7.4012639e-16
+ ub1 = 2.6826436e-19
+ uc1 = 8.9789043e-11
+ drout = 0.56
+ lags = 4.7673289e-7
+ wku0we = 1.5e-11
+ tpb = 0.0016
+ wa0 = 5.2465177e-8
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ ute = -0.817454
+ paigc = 1.4961177e-18
+ lcit = 1.6e-11
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 3.8961851e-9
+ tnoimod = 0
+ mobmod = 0
+ wlc = 0
+ wln = 1
+ wu0 = 5.5067755e-11
+ xgl = -8.2e-9
+ xgw = 0
+ kt1l = 0
+ wua = -5.1699586e-17
+ wub = 1.2857705e-26
+ wuc = 3.3174666e-18
+ wud = 0
+ voffl = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ wpdiblc2 = 3.5925269e-10
+ cigbinv = 0.006
+ weta0 = 1.9163288999999998e-9
+ wetab = 2.9133333e-9
+ lint = 6.5375218e-9
+ lpclm = 0
+ lkt1 = -8.6254893e-9
+ lkt2 = -1.4709041e-9
+ lmax = 8.9991e-6
+ lmin = 8.9908e-7
+ lpe0 = 6.44e-8
+ cgidl = 1
+ lpeb = 0
+ version = 4.5
+ tempmod = 0
+ minv = -0.33
+ wtvfbsdoff = 0
+ laigsd = -1.8524358e-14
+ lua1 = 1.5667589e-15
+ lub1 = -2.759143e-24
+ luc1 = -7.2890309e-17
+ ndep = 1e+18
+ wkvth0we = 0.0
+ lute = 1.5402209e-8
+ lwlc = 0
+ pbswd = 0.9
+ pbsws = 0.9
+ moin = 5.5538
+ aigbacc = 0.012071
+ ltvfbsdoff = 0
+ trnqsmod = 0
+ nigc = 2.291
+ pdits = 0
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ noff = 2.2684
+ cigsd = 0.013281
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ aigbinv = 0.009974
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ pags = -1.92428e-14
+ ntox = 1.0
+ pcit = -8.000000000000001e-19
+ rgatemod = 0
+ pclm = 1.101657
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ ptvfbsdoff = 0
+ tnjtsswg = 1
+ phin = 0.15
+ tnoia = 0
+ pkt1 = -2.8522213999999998e-15
+ pkt2 = 2.4239149e-16
+ peta0 = -1.6e-17
+ toxref = 3e-9
+ wketa = -2.0595747e-9
+ poxedge = 1
+ tpbsw = 0.0025
+ cjswd = 5.3856e-11
+ cjsws = 5.3856e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ rbdb = 50
+ pua1 = -1.1776704e-22
+ binunit = 2
+ prwb = 0
+ pub1 = 2.7996299e-31
+ prwg = 0
+ puc1 = 9.811687e-24
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ pute = 1.5923616e-14
+ rdsw = 200
+ tvfbsdoff = 0.1
+ ltvoff = -3.3500511e-10
+ scref = 1e-6
+ pigcd = 2.572
+ rshg = 14.1
+ aigsd = 0.0063632604
+ lku0we = 1.8e-11
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ epsrox = 3.9
+ lvoff = -2.4480721e-8
+ a0 = 2.6314952
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ rdsmod = 0
+ wvfbsdoff = 0
+ at = 72000
+ cf = 8.17e-11
+ lvsat = 8.000000000000001e-6
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.016004612
+ k3 = -2.5823
+ em = 20000000.0
+ lvfbsdoff = 0
+ lvth0 = -1.4106904000000001e-8
+ igbmod = 1
+ ll = 0
+ lw = 0
+ u0 = 0.0095363075
+ w0 = 0
+ ua = -1.8414289e-10
+ ub = 1.2263153e-18
+ uc = -3.3458683e-12
+ ud = 0
+ ijthsfwd = 0.01
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 3.4e-9
+ delta = 0.018814
+ laigc = -5.3027874e-11
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ rnoia = 0
+ rnoib = 0
+ pbswgd = 0.8
+ pbswgs = 0.8
+ tnom = 25
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ igcmod = 1
+ pketa = 1.0887638e-15
+ ngate = 1.7e+20
+ ngcon = 1
+ ijthsrev = 0.01
+ wpclm = 7.1298978e-9
+ njtsswg = 6.489
+ gbmin = 1e-12
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ wags = 7.3346686e-9
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.00084883969
+ pdiblcb = 0
+ paigsd = -1.2880862e-20
+ voff = -0.10099712
+ acde = 0.5
+ ppdiblc2 = -2.0561872e-16
+ vsat = 108525.44
+ wint = 0
+ permod = 1
+ vth0 = -0.39532868000000004
+ wkt1 = -2.7375492e-9
+ wkt2 = -7.5529568e-10
+ wmax = 2.726e-7
+ aigc = 0.0068361189
+ wmin = 1.08e-7
+ bigbacc = 0.0054401
+ tvoff = 0.0025796189
+ kvth0we = -0.00022
+ wua1 = -4.222676e-17
+ wub1 = -1.3803658e-25
+ wuc1 = -1.3210867e-17
+ xjbvd = 1
+ xjbvs = 1
+ voffcv = -0.125
+ wpemod = 1
+ lk2we = 0.0
+ lintnoi = -5e-9
+ bigc = 0.0012521
+ wute = -7.8294814e-8
+ bigbinv = 0.00149
+ pkvth0we = 0.0
+ wwlc = 0
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ cdsc = 0
+ ku0we = -0.0007
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ beta0 = 13.32
+ leta0 = -4.8e-10
+ vfbsdoff = 0.01
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigc = 0.15259
+ ppclm = 0
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ paramchk = 1
+ tpbswg = 0.001
+ )

.model pch_fs_35 pmos (
+ level = 54
+ cjsws = 5.3856e-11
+ cjswgd = 1.9113600000000002e-10
+ pku0we = 0.0
+ cjswgs = 1.9113600000000002e-10
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ ndep = 1e+18
+ lute = -1.0958354e-8
+ lwlc = 0
+ moin = 5.5538
+ ijthsrev = 0.01
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ tvfbsdoff = 0.1
+ nigc = 2.291
+ mjswgd = 0.95
+ mjswgs = 0.95
+ tcjswg = 0.00128
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ scref = 1e-6
+ pags = 1.1742809e-13
+ ppdiblc2 = -6.1367245e-16
+ pigcd = 2.572
+ ntox = 1.0
+ aigsd = 0.0063632396
+ pcit = -8.000000000000001e-19
+ pclm = 1.101657
+ lvoff = -2.4340257e-9
+ phin = 0.15
+ wvfbsdoff = 0
+ njtsswg = 6.489
+ lvfbsdoff = 0
+ lvsat = 8.000000000000001e-6
+ lvth0 = -2.6799405e-10
+ pkt1 = 5.7073332e-15
+ pkt2 = -5.7270183e-16
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ delta = 0.018814
+ fprout = 200
+ laigc = -3.3884553e-11
+ xrcrg1 = 12
+ xrcrg2 = 1
+ ckappad = 0.6
+ ckappas = 0.6
+ rnoia = 0
+ rnoib = 0
+ pdiblc1 = 0
+ pdiblc2 = 0.0027845581
+ pdiblcb = 0
+ pkvth0we = 0.0
+ rbdb = 50
+ pua1 = -9.8048843e-24
+ prwb = 0
+ pub1 = -2.3189739e-32
+ prwg = 0
+ puc1 = -4.5795492e-24
+ pketa = -3.0075994e-15
+ rbpb = 50
+ rbpd = 50
+ ngate = 1.7e+20
+ rbps = 50
+ rbsb = 50
+ wtvoff = -2.2790108e-10
+ pvag = 2.1
+ pute = -9.4649237e-15
+ ngcon = 1
+ wpclm = 7.1298978e-9
+ rdsw = 200
+ vfbsdoff = 0.01
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ bigbacc = 0.0054401
+ capmod = 2
+ wku0we = 1.5e-11
+ kvth0we = -0.00022
+ mobmod = 0
+ paramchk = 1
+ lintnoi = -5e-9
+ rshg = 14.1
+ bigbinv = 0.00149
+ wtvfbsdoff = 0
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ ltvfbsdoff = 0
+ ijthdfwd = 0.01
+ tvoff = 0.0027416725
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ tnom = 25
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ ijthdrev = 0.01
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = -4.8e-10
+ lpdiblc2 = 4.574275e-9
+ ptvfbsdoff = 0
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ nfactor = 1
+ ppclm = 0
+ wags = -1.4622812e-7
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ voff = -0.12576869
+ acde = 0.5
+ vsat = 108525.44
+ wint = 0
+ vth0 = -0.41087802
+ wkt1 = -1.2355026e-8
+ wkt2 = 1.605395e-10
+ dmcgt = 0
+ wmax = 2.726e-7
+ tcjsw = 9.34e-5
+ lkvth0we = 3e-12
+ aigc = 0.0068146096
+ wmin = 1.08e-7
+ nigbacc = 10
+ toxref = 3e-9
+ wua1 = -1.6353255e-16
+ wub1 = 2.0258446e-25
+ wuc1 = 2.9590615e-18
+ acnqsmod = 0
+ bigsd = 0.0003327
+ bigc = 0.0012521
+ wute = -4.9768365e-8
+ nigbinv = 2.171
+ wwlc = 0
+ wvoff = 3.4766421e-9
+ rbodymod = 0
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ wvsat = -0.0013318206
+ xtid = 3
+ xtis = 3
+ wvth0 = -4.7116532000000006e-9
+ ltvoff = -4.7923289e-10
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigc = 0.15259
+ waigc = 2.7104678e-12
+ fnoimod = 1
+ eigbinv = 1.1
+ pvfbsdoff = 0
+ lketa = 4.197898e-9
+ xpart = 1
+ lku0we = 1.8e-11
+ epsrox = 3.9
+ wpdiblc2 = 8.1773971e-10
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ ags = 1.7348065
+ dmdg = 0
+ egidl = 0.001
+ cjd = 0.001421376
+ rdsmod = 0
+ cit = -8.7888889e-5
+ cjs = 0.001421376
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 1.0572421799999999e-8
+ igbmod = 1
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ k2we = 5e-5
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ dsub = 0.5
+ dtox = 3.91e-10
+ pbswgd = 0.8
+ la0 = -1.044589e-6
+ cigbacc = 0.245
+ pbswgs = 0.8
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0.00064
+ kt1 = -0.11040563
+ kt2 = -0.048714998
+ lk2 = 3.4090726e-9
+ llc = 0
+ lln = 1
+ lu0 = -1.8180818e-9
+ mjd = 0.335
+ mjs = 0.335
+ lua = -6.2776752e-16
+ lub = 4.4518935e-25
+ luc = 5.1177769e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ igcmod = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 1.0817056e-13
+ wkvth0we = 0.0
+ nsd = 1e+20
+ pbd = 0.75
+ tnoimod = 0
+ pat = 0
+ pbs = 0.75
+ pk2 = -1.5480351e-16
+ eta0 = 0.10792519
+ etab = -0.13555556
+ pu0 = 1.5955157e-16
+ prt = 0
+ pua = 4.4574845e-23
+ pub = -2.7161351e-32
+ puc = -4.8372521e-24
+ pud = 0
+ rsh = 15.2
+ trnqsmod = 0
+ tcj = 0.000832
+ ua1 = 2.771768e-9
+ ub1 = -3.1924567e-18
+ uc1 = -6.2120134e-12
+ cigbinv = 0.006
+ tpb = 0.0016
+ wa0 = -1.0464262e-7
+ ute = -0.78783539
+ pvoff = -9.7175093e-16
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 4.174453e-9
+ wlc = 0
+ wln = 1
+ wu0 = -8.9929205e-11
+ xgl = -8.2e-9
+ xgw = 0
+ wua = -7.0620672e-17
+ wub = -4.621089e-27
+ wuc = 8.8883858e-18
+ wud = 0
+ cdscb = 0
+ cdscd = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ pvsat = 0
+ a0 = 3.3624733
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ wk2we = 0.0
+ pvth0 = 5.5307120000000006e-17
+ at = 72000
+ cf = 8.17e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.013259817
+ k3 = -2.5823
+ em = 20000000.0
+ drout = 0.56
+ version = 4.5
+ ll = 0
+ lw = 0
+ u0 = 0.012698186
+ w0 = 0
+ ua = 4.4026063e-10
+ ub = 1.2150282e-18
+ uc = -4.4814963e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ paigc = 4.1038726e-19
+ xw = 3.4e-9
+ tempmod = 0
+ voffl = 0
+ rgatemod = 0
+ permod = 1
+ tnjtsswg = 1
+ weta0 = 1.9163288999999998e-9
+ wetab = 2.9133333e-9
+ aigbacc = 0.012071
+ lpclm = 0
+ cgidl = 1
+ voffcv = -0.125
+ wpemod = 1
+ aigbinv = 0.009974
+ pbswd = 0.9
+ pbsws = 0.9
+ keta = -0.035939983
+ pdits = 0
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ lags = -3.1625612e-7
+ tpbswg = 0.001
+ poxedge = 1
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 9.8671111e-11
+ kt1l = 0
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ binunit = 2
+ lint = 6.5375218e-9
+ ptvoff = 8.8703803e-17
+ lkt1 = -6.2618035e-8
+ lkt2 = -3.1463267e-9
+ tnoia = 0
+ lmax = 8.9908e-7
+ waigsd = 1.9716411e-12
+ lmin = 4.4908e-7
+ ijthsfwd = 0.01
+ peta0 = -1.6e-17
+ lpe0 = 6.44e-8
+ lpeb = 0
+ wketa = 2.5430806e-9
+ diomod = 1
+ tpbsw = 0.0025
+ minv = -0.33
+ lua1 = -1.8157361e-16
+ lub1 = 3.2089876e-25
+ luc1 = 1.2550631e-17
+ pditsd = 0
+ cjswd = 5.3856e-11
+ pditsl = 0
+ )

.model pch_fs_36 pmos (
+ level = 54
+ ags = 0.79842724
+ pvfbsdoff = 0
+ wcit = 5.8162887e-11
+ lketa = -1.0850486e-8
+ cigbacc = 0.245
+ cjd = 0.001421376
+ cit = -0.00049977211
+ cjs = 0.001421376
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ voff = -0.11894985
+ xpart = 1
+ dlc = 1.38228675e-8
+ k3b = 2.1176
+ acde = 0.5
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ rgatemod = 0
+ tnjtsswg = 1
+ vsat = 108525.44
+ tnoimod = 0
+ wint = 0
+ vth0 = -0.41750626
+ egidl = 0.001
+ wkt1 = 8.365112e-10
+ wkt2 = -1.4765978e-9
+ la0 = -3.2362015e-7
+ wmax = 2.726e-7
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0.00064
+ aigc = 0.0068096243
+ wmin = 1.08e-7
+ kt1 = -0.25321364
+ kt2 = -0.04359324
+ lk2 = -2.273089999999996e-11
+ llc = -1.18e-13
+ lln = 0.7
+ cigbinv = 0.006
+ lu0 = -4.5139607999999997e-10
+ mjd = 0.335
+ mjs = 0.335
+ lua = -1.7021816e-16
+ lub = 1.0550853e-25
+ luc = -1.2975077e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ fprout = 200
+ njs = 1.02
+ pa0 = -3.1370244e-14
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ pk2 = 1.4083403e-16
+ xrcrg1 = 12
+ xrcrg2 = 1
+ pu0 = -1.3937081e-17
+ prt = 0
+ pua = 4.7117679e-24
+ pub = -8.7289665e-33
+ puc = -3.0945045e-25
+ pud = 0
+ wua1 = -2.3000717e-16
+ wub1 = 1.2114667e-25
+ wuc1 = -1.9684753e-17
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 2.6350858e-9
+ ub1 = -2.2549964e-18
+ uc1 = 3.1191962e-11
+ bigc = 0.0012521
+ wute = -1.1762912e-7
+ version = 4.5
+ tpb = 0.0016
+ wa0 = 2.1249557e-7
+ wwlc = 0
+ ute = -0.71022675
+ wtvoff = -1.1036076e-10
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 3.5025496e-9
+ tempmod = 0
+ wlc = 0
+ wln = 1
+ wu0 = 3.0436319e-10
+ xgl = -8.2e-9
+ xgw = 0
+ wua = 1.9977231e-17
+ wub = -4.6512873e-26
+ wuc = -1.4020724e-18
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ wtvfbsdoff = 0
+ aigbacc = 0.012071
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigc = 0.15259
+ pvoff = 1.15942711e-16
+ capmod = 2
+ cdscb = 0
+ cdscd = 0
+ wku0we = 1.5e-11
+ pvsat = 0
+ wk2we = 0.0
+ pvth0 = -3.5393785e-16
+ ltvfbsdoff = 0
+ drout = 0.56
+ mobmod = 0
+ paigc = -1.759214e-19
+ aigbinv = 0.009974
+ voffl = 0
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ weta0 = 1.9163288999999998e-9
+ wetab = 2.9133333e-9
+ lpclm = 0
+ k2we = 5e-5
+ ijthsfwd = 0.01
+ cgidl = 1
+ dsub = 0.5
+ ptvfbsdoff = 0
+ dtox = 3.91e-10
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ poxedge = 1
+ eta0 = 0.10792519
+ pbswd = 0.9
+ etab = -0.13555556
+ pbsws = 0.9
+ ijthsrev = 0.01
+ binunit = 2
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ pdits = 0
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ ppdiblc2 = 9.2177422e-17
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ tnoia = 0
+ toxref = 3e-9
+ peta0 = -1.6e-17
+ wketa = -1.9938172e-9
+ tpbsw = 0.0025
+ cjswd = 5.3856e-11
+ cjsws = 5.3856e-11
+ pkvth0we = 0.0
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ tvfbsdoff = 0.1
+ ltvoff = -1.9203223e-10
+ vfbsdoff = 0.01
+ njtsswg = 6.489
+ keta = -0.0017391106
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ lags = 9.5750741e-8
+ lku0we = 1.8e-11
+ paramchk = 1
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ scref = 1e-6
+ ckappad = 0.6
+ ckappas = 0.6
+ lcit = 2.7989972999999997e-10
+ pdiblc1 = 0
+ pdiblc2 = 0.016049816
+ epsrox = 3.9
+ pdiblcb = 0
+ pigcd = 2.572
+ kt1l = 0
+ aigsd = 0.0063632396
+ rdsmod = 0
+ lvoff = -5.4343156e-9
+ wvfbsdoff = 0
+ lint = 9.7879675e-9
+ igbmod = 1
+ lvfbsdoff = 0
+ lkt1 = 2.1786599999999996e-10
+ lkt2 = -5.3999005e-9
+ lvsat = 8.000000000000001e-6
+ lmax = 4.4908e-7
+ lvth0 = 2.6484329e-9
+ lmin = 2.1577e-7
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ ijthdfwd = 0.01
+ lpe0 = 6.44e-8
+ delta = 0.018814
+ bigbacc = 0.0054401
+ lpeb = 0
+ pbswgd = 0.8
+ laigc = -3.1691048e-11
+ pbswgs = 0.8
+ rnoia = 0
+ rnoib = 0
+ minv = -0.33
+ igcmod = 1
+ lua1 = -1.2143343e-16
+ lub1 = -9.158653e-26
+ luc1 = -3.907118e-18
+ kvth0we = -0.00022
+ ndep = 1e+18
+ lute = -4.5106156e-8
+ pketa = -1.0113644e-15
+ ngate = 1.7e+20
+ lwlc = 0
+ lintnoi = -5e-9
+ moin = 5.5538
+ ijthdrev = 0.01
+ ngcon = 1
+ bigbinv = 0.00149
+ wpclm = 7.1298978e-9
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ nigc = 2.291
+ lpdiblc2 = -1.262443e-9
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ pags = 5.2660461e-14
+ permod = 1
+ ntox = 1.0
+ pcit = -2.639167e-17
+ pclm = 1.101657
+ phin = 0.15
+ lkvth0we = 3e-12
+ pkt1 = -9.70475e-17
+ pkt2 = 1.4763857e-16
+ voffcv = -0.125
+ wpemod = 1
+ tvoff = 0.0020889601
+ nfactor = 1
+ xjbvd = 1
+ acnqsmod = 0
+ xjbvs = 1
+ lk2we = 0.0
+ a0 = 1.7239078
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ rbdb = 50
+ pua1 = 1.9443948e-23
+ prwb = 0
+ pub1 = 1.2643651e-32
+ prwg = 0
+ at = 72000
+ puc1 = 5.3837292e-24
+ cf = 8.17e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.0054602636
+ k3 = -2.5823
+ em = 20000000.0
+ rbpb = 50
+ rbpd = 50
+ ll = -1.18e-13
+ lw = 0
+ rbps = 50
+ u0 = 0.009592082
+ rbsb = 50
+ pvag = 2.1
+ w0 = 0
+ rbodymod = 0
+ ua = -5.9962427e-10
+ ub = 1.98703e-18
+ uc = 1.0098696e-10
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ pute = 2.0393808e-14
+ xw = 3.4e-9
+ rdsw = 200
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = -4.8e-10
+ nigbacc = 10
+ ppclm = 0
+ tpbswg = 0.001
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ rshg = 14.1
+ nigbinv = 2.171
+ wpdiblc2 = -7.8646151e-10
+ ptvoff = 3.6984079e-17
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ waigsd = 1.9716411e-12
+ diomod = 1
+ fnoimod = 1
+ pditsd = 0
+ pditsl = 0
+ bigsd = 0.0003327
+ cjswgd = 1.9113600000000002e-10
+ pku0we = 0.0
+ tnom = 25
+ cjswgs = 1.9113600000000002e-10
+ eigbinv = 1.1
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ wkvth0we = 0.0
+ wvoff = 1.0046111e-9
+ trnqsmod = 0
+ wvsat = -0.0013318206
+ mjswgd = 0.95
+ wvth0 = -3.781551e-9
+ mjswgs = 0.95
+ tcjswg = 0.00128
+ waigc = 4.0429874e-12
+ wags = 9.7102189e-10
+ )

.model pch_fs_37 pmos (
+ level = 54
+ fprout = 200
+ lvth0 = 5.2874905e-9
+ xrcrg1 = 12
+ xrcrg2 = 1
+ delta = 0.018814
+ wtvfbsdoff = 0
+ laigc = -4.357169e-12
+ rnoia = 0
+ rnoib = 0
+ acnqsmod = 0
+ wtvoff = 1.2048366e-10
+ ltvfbsdoff = 0
+ pketa = 4.1278959e-16
+ ngate = 1.7e+20
+ rbodymod = 0
+ ngcon = 1
+ wpclm = 6.8691006e-8
+ capmod = 2
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ wku0we = 1.5e-11
+ keta = -0.058692164
+ mobmod = 0
+ nfactor = 1
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 4.1291477e-11
+ ptvfbsdoff = 0
+ kt1l = 0
+ wpdiblc2 = -7.28246e-10
+ lint = 9.7879675e-9
+ lkt1 = -5.1570694e-9
+ lkt2 = -3.7791597e-9
+ lmax = 2.1577e-7
+ lmin = 9e-8
+ lpe0 = 6.44e-8
+ nigbacc = 10
+ lpeb = 0
+ tvoff = 0.0011827459
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ minv = -0.33
+ lua1 = -2.1218464e-16
+ lub1 = 2.7818737e-25
+ luc1 = 2.2554944e-17
+ ndep = 1e+18
+ wkvth0we = 0.0
+ lute = 1.5508066e-9
+ lwlc = 0
+ moin = 5.5538
+ nigbinv = 2.171
+ ku0we = -0.0007
+ trnqsmod = 0
+ beta0 = 13.32
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ nigc = 2.291
+ leta0 = -4.8e-10
+ ppclm = -1.2989269e-14
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ fnoimod = 1
+ eigbinv = 1.1
+ ntox = 1.0
+ rgatemod = 0
+ pcit = 1.0414196e-17
+ pclm = 0.85425247
+ tnjtsswg = 1
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ phin = 0.15
+ toxref = 3e-9
+ pkt1 = -2.717336e-16
+ pkt2 = 3.7767926e-16
+ bigsd = 0.0003327
+ cigbacc = 0.245
+ rbdb = 50
+ pua1 = 2.6827919e-23
+ prwb = 0
+ pub1 = -3.4278711e-32
+ prwg = 0
+ puc1 = -2.7535024e-24
+ wvoff = 8.5374562e-10
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ pute = -4.2802262e-16
+ ltvoff = -8.1627e-13
+ rdsw = 200
+ tnoimod = 0
+ wvsat = -0.00089129698
+ ags = 1.2522222
+ wvth0 = -4.810948000000001e-9
+ cjd = 0.001421376
+ cit = 0.00063107268
+ cjs = 0.001421376
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 1.38228675e-8
+ waigc = 1.4660694e-11
+ k3b = 2.1176
+ cigbinv = 0.006
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ pvfbsdoff = 0
+ lku0we = 1.8e-11
+ lketa = 1.1666086e-9
+ epsrox = 3.9
+ la0 = 6.219346e-9
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = -0.0069043287
+ xpart = 1
+ kt1 = -0.22773883
+ kt2 = -0.051274476
+ lk2 = 3.9911471e-9
+ llc = -1.18e-13
+ lln = 0.7
+ lu0 = -1.6394862000000002e-10
+ mjd = 0.335
+ version = 4.5
+ mjs = 0.335
+ lua = 1.3101868e-17
+ lub = -8.7271368e-26
+ luc = -1.2812174e-17
+ lud = 0
+ rshg = 14.1
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = -2.0637395e-14
+ rdsmod = 0
+ nsd = 1e+20
+ pbd = 0.75
+ tempmod = 0
+ pat = -5.0045721e-10
+ pbs = 0.75
+ pk2 = 4.0368065e-17
+ egidl = 0.001
+ igbmod = 1
+ pu0 = -5.2679707e-18
+ prt = 0
+ pua = -4.0286539e-24
+ pub = 7.5106005e-33
+ puc = 1.4358513e-24
+ pud = 0
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 3.0651863e-9
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ ub1 = -4.0074881e-18
+ uc1 = -9.4220652e-11
+ tpb = 0.0016
+ aigbacc = 0.012071
+ wa0 = 1.6162969e-7
+ pbswgd = 0.8
+ pbswgs = 0.8
+ ute = -0.93134979
+ ijthsfwd = 0.01
+ wat = 0.0023718351
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 3.9786916e-9
+ wlc = 0
+ wln = 1
+ wu0 = 2.6327735e-10
+ xgl = -8.2e-9
+ xgw = 0
+ wua = 6.1401032e-17
+ wub = -1.2347765e-25
+ wuc = -9.6736445e-18
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ igcmod = 1
+ tnom = 25
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ aigbinv = 0.009974
+ ijthsrev = 0.01
+ pvoff = 1.4777532e-16
+ cdscb = 0
+ cdscd = 0
+ pvsat = -9.2948987e-11
+ wags = 2.5054667e-7
+ wk2we = 0.0
+ pvth0 = -1.3673509200000002e-16
+ drout = 0.56
+ wcit = -1.162725e-10
+ paigc = -2.4162575e-18
+ permod = 1
+ voff = -0.1339517
+ acde = 0.5
+ ppdiblc2 = 7.9894307e-17
+ voffl = 0
+ poxedge = 1
+ vsat = 106518.57
+ wint = 0
+ vth0 = -0.43001365
+ weta0 = 1.9163288999999998e-9
+ wetab = 2.9133333e-9
+ wkt1 = 1.664079e-9
+ wkt2 = -2.566838e-9
+ wmax = 2.726e-7
+ lpclm = 5.2201277e-8
+ binunit = 2
+ aigc = 0.0066800799
+ wmin = 1.08e-7
+ voffcv = -0.125
+ wpemod = 1
+ cgidl = 1
+ wua1 = -2.6500229e-16
+ wub1 = 3.4352994e-25
+ wuc1 = 1.8880326e-17
+ bigc = 0.0012521
+ wute = -1.8947457e-8
+ pkvth0we = 0.0
+ wwlc = 0
+ pbswd = 0.9
+ pbsws = 0.9
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ vfbsdoff = 0.01
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigc = 0.15259
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ pdits = 0
+ tpbswg = 0.001
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ paramchk = 1
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ ptvoff = -1.1725409e-17
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ a0 = 0.16068118
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ waigsd = 1.9716411e-12
+ at = 107755.11
+ cf = 8.17e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.024483382
+ k3 = -2.5823
+ em = 20000000.0
+ ll = -1.18e-13
+ lw = 0
+ u0 = 0.0082297718
+ tnoia = 0
+ w0 = 0
+ ua = -1.4684396e-9
+ ub = 2.9006788e-18
+ uc = 1.0021491e-10
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 3.4e-9
+ diomod = 1
+ k2we = 5e-5
+ ijthdfwd = 0.01
+ peta0 = -1.6e-17
+ njtsswg = 6.489
+ dsub = 0.5
+ dtox = 3.91e-10
+ wketa = -8.743362e-9
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.9113600000000002e-10
+ pku0we = 0.0
+ cjswgs = 1.9113600000000002e-10
+ tpbsw = 0.0025
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ cjswd = 5.3856e-11
+ cjsws = 5.3856e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.01690182
+ eta0 = 0.10792519
+ pdiblcb = 0
+ etab = -0.13555556
+ tvfbsdoff = 0.1
+ ijthdrev = 0.01
+ mjswgd = 0.95
+ mjswgs = 0.95
+ lpdiblc2 = -1.4422174e-9
+ tcjswg = 0.00128
+ bigbacc = 0.0054401
+ scref = 1e-6
+ pigcd = 2.572
+ aigsd = 0.0063632396
+ kvth0we = -0.00022
+ wvfbsdoff = 0
+ lvoff = -2.268926e-9
+ lintnoi = -5e-9
+ lvfbsdoff = 0
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ lkvth0we = 3e-12
+ lvsat = 0.00043143718999999996
+ )

.model pch_fs_38 pmos (
+ level = 54
+ poxedge = 1
+ ptvfbsdoff = 0
+ rdsw = 200
+ capmod = 2
+ vfbsdoff = 0.01
+ wku0we = 1.5e-11
+ pvoff = -1.2373467e-16
+ binunit = 2
+ cdscb = 0
+ cdscd = 0
+ mobmod = 0
+ pvsat = 1.729604e-10
+ wk2we = 0.0
+ pvth0 = -6.3236866e-17
+ drout = 0.56
+ paramchk = 1
+ paigc = -1.1563004e-18
+ voffl = 0
+ rshg = 14.1
+ weta0 = 1.2733501000000001e-8
+ wetab = 4.1458967e-9
+ lpclm = -1.0127779e-7
+ ijthdfwd = 0.01
+ jtsswgd = 1.75e-7
+ cgidl = 1
+ jtsswgs = 1.75e-7
+ tnom = 25
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ pbswd = 0.9
+ pbsws = 0.9
+ ijthdrev = 0.01
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ lpdiblc2 = -1.4113545e-11
+ pdits = 0
+ cigsd = 0.013281
+ wags = 2.5054667e-7
+ dvt0w = 0
+ dvt1w = 0
+ njtsswg = 6.489
+ dvt2w = 0
+ wcit = 7.0487744e-11
+ xtsswgd = 0.32
+ voff = -0.14478455
+ xtsswgs = 0.32
+ acde = 0.5
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ ckappad = 0.6
+ ckappas = 0.6
+ vsat = 137363.5
+ wint = 0
+ pdiblc1 = 0
+ pdiblc2 = 0.0017092259
+ vth0 = -0.36680653
+ pdiblcb = 0
+ wkt1 = -1.350742e-8
+ wkt2 = 1.8825744e-9
+ toxref = 3e-9
+ wmax = 2.726e-7
+ lkvth0we = 3e-12
+ aigc = 0.0067219883
+ wmin = 1.08e-7
+ tnoia = 0
+ peta0 = -1.0328142000000001e-15
+ petab = -1.1586096e-16
+ wketa = -6.6698086e-9
+ wua1 = 1.6631395e-16
+ wub1 = -2.121384e-25
+ wuc1 = 2.5860689e-17
+ tpbsw = 0.0025
+ acnqsmod = 0
+ bigbacc = 0.0054401
+ cjswd = 5.3856e-11
+ bigc = 0.0012521
+ cjsws = 5.3856e-11
+ wute = -6.1363432e-8
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ wwlc = 0
+ tvfbsdoff = 0.1
+ ltvoff = 3.7319947e-11
+ rbodymod = 0
+ kvth0we = -0.00022
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ lintnoi = -5e-9
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ bigbinv = 0.00149
+ cigc = 0.15259
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ lku0we = 1.8e-11
+ epsrox = 3.9
+ scref = 1e-6
+ pigcd = 2.572
+ aigsd = 0.0063632396
+ rdsmod = 0
+ wpdiblc2 = 8.0253658e-11
+ igbmod = 1
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ lvoff = -1.2506377e-9
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ lvsat = -0.0024679865
+ pbswgd = 0.8
+ pbswgs = 0.8
+ lvth0 = -6.539787e-10
+ k2we = 5e-5
+ delta = 0.018814
+ laigc = -8.2965642e-12
+ dsub = 0.5
+ igcmod = 1
+ dtox = 3.91e-10
+ rnoia = 0
+ rnoib = 0
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ nfactor = 1
+ wkvth0we = 0.0
+ pketa = 2.1787556e-16
+ ngate = 1.7e+20
+ eta0 = 0.024468866
+ etab = -0.22797789
+ ngcon = 1
+ wpclm = -1.6917696e-7
+ trnqsmod = 0
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ nigbacc = 10
+ permod = 1
+ rgatemod = 0
+ tnjtsswg = 1
+ nigbinv = 2.171
+ voffcv = -0.125
+ wpemod = 1
+ tvoff = 0.00077704148
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ fnoimod = 1
+ eigbinv = 1.1
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = 7.364893999999999e-9
+ letab = 8.6876992e-9
+ tpbswg = 0.001
+ ppclm = 9.3703198e-15
+ keta = -0.049241031
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 1.4330569e-10
+ kt1l = 0
+ ptvoff = 1.952106e-17
+ cigbacc = 0.245
+ waigsd = 1.9716411e-12
+ dmcgt = 0
+ lint = 0
+ tcjsw = 9.34e-5
+ tnoimod = 0
+ lkt1 = -7.0746074e-9
+ lkt2 = 9.2375447e-10
+ diomod = 1
+ lmax = 9e-8
+ lmin = 5.4e-8
+ ijthsfwd = 0.01
+ lpe0 = 6.44e-8
+ pditsd = 0
+ pditsl = 0
+ lpeb = 0
+ cigbinv = 0.006
+ cjswgd = 1.9113600000000002e-10
+ pku0we = 0.0
+ cjswgs = 1.9113600000000002e-10
+ bigsd = 0.0003327
+ minv = -0.33
+ ags = 1.2522222
+ lua1 = 1.5814311e-16
+ lub1 = -2.3663254e-25
+ luc1 = 3.1466117e-17
+ cjd = 0.001421376
+ cit = -0.00045418481
+ cjs = 0.001421376
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ ndep = 1e+18
+ bvs = 8.2
+ lute = -1.2895214e-8
+ dlc = 4.0349e-9
+ wvoff = 3.7421498e-9
+ k3b = 2.1176
+ lwlc = 0
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ version = 4.5
+ moin = 5.5538
+ mjswgd = 0.95
+ mjswgs = 0.95
+ ijthsrev = 0.01
+ tempmod = 0
+ wvsat = -0.0037201203
+ nigc = 2.291
+ tcjswg = 0.00128
+ wvth0 = -5.592844000000001e-9
+ la0 = 3.4503642e-8
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = -0.0074128059
+ kt1 = -0.20733948
+ kt2 = -0.10130548
+ lk2 = 5.867862999999999e-9
+ waigc = 1.256895e-12
+ llc = 0
+ lln = 1
+ a0 = -0.1402156
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ lu0 = 4.500914e-11
+ mjd = 0.335
+ mjs = 0.335
+ lua = 1.1003971e-16
+ lub = -1.3258131e-25
+ luc = -1.072064e-17
+ at = 113164.44
+ lud = 0
+ cf = 8.17e-11
+ lwc = 0
+ pvfbsdoff = 0
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.044448444
+ k3 = -2.5823
+ lwl = 0
+ lwn = 1
+ em = 20000000.0
+ aigbacc = 0.012071
+ njd = 1.02
+ njs = 1.02
+ ll = 0
+ noff = 2.2684
+ pa0 = -6.959911e-15
+ lw = 0
+ u0 = 0.006006816900000001
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ w0 = 0
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 1.1859675e-9
+ ua = -2.4996932e-9
+ ub = 3.3826995e-18
+ uc = 7.7964547e-11
+ ud = 0
+ pbs = 0.75
+ pk2 = -8.547569e-17
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 3.4e-9
+ pu0 = 1.7354187e-18
+ prt = 0
+ lketa = 2.7820203e-10
+ pua = -5.4706466e-24
+ pub = 7.2761107e-33
+ puc = 2.7207836e-25
+ pud = 0
+ wtvfbsdoff = 0
+ xpart = 1
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = -8.7447052e-10
+ ub1 = 1.4693195e-18
+ uc1 = -1.8902037e-10
+ ppdiblc2 = 3.8953385e-18
+ ntox = 1.0
+ tpb = 0.0016
+ pcit = -7.1412667e-18
+ pclm = 2.4870084
+ wa0 = 1.612455e-8
+ ute = -0.77766872
+ wat = -0.015568853
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 5.3174549e-9
+ aigbinv = 0.009974
+ wlc = 0
+ egidl = 0.001
+ wln = 1
+ wu0 = 1.8877321e-10
+ xgl = -8.2e-9
+ xgw = 0
+ wua = 7.6741379e-17
+ wub = -1.2098307e-25
+ wuc = 2.7069183e-18
+ wud = 0
+ wwc = 0
+ ltvfbsdoff = 0
+ wwl = 0
+ wwn = 1
+ phin = 0.15
+ fprout = 200
+ xrcrg1 = 12
+ xrcrg2 = 1
+ pkt1 = 1.1543873e-15
+ pkt2 = -4.056551e-17
+ wtvoff = -2.1192558e-10
+ pkvth0we = 0.0
+ rbdb = 50
+ pua1 = -1.3715808e-23
+ prwb = 0
+ pub1 = 1.7954113e-32
+ prwg = 0
+ puc1 = -3.4096566e-24
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ pute = 3.5590791e-15
+ )

.model pch_fs_39 pmos (
+ level = 54
+ fnoimod = 1
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ eigbinv = 1.1
+ k2we = 5e-5
+ ijthsfwd = 0.01
+ tvoff = 0.00092289205
+ dsub = 0.5
+ dtox = 3.91e-10
+ xjbvd = 1
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ xjbvs = 1
+ lk2we = 0.0
+ eta0 = 0.19463541
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ etab = -0.16706384
+ ijthsrev = 0.01
+ cigbacc = 0.245
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = -2.5047657e-9
+ letab = 5.1546845e-9
+ tnoimod = 0
+ ppclm = 7.8094068e-15
+ dlcig = 2.5e-9
+ cigbinv = 0.006
+ bgidl = 1834800000.0
+ ppdiblc2 = 0
+ toxref = 3e-9
+ version = 4.5
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ tempmod = 0
+ ags = 1.2522222
+ cjd = 0.001421376
+ cit = -0.0026753087
+ cjs = 0.001421376
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 4.0349e-9
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ aigbacc = 0.012071
+ bigsd = 0.0003327
+ pkvth0we = 0.0
+ la0 = -1.4904033e-7
+ ltvoff = 2.8860613e-11
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0.010012509
+ kt1 = -0.53950997
+ kt2 = -0.12590838
+ lk2 = 4.5365993e-9
+ wvoff = 1.4341134e-10
+ llc = 0
+ lln = 1
+ lu0 = 4.1571089e-10
+ mjd = 0.335
+ mjs = 0.335
+ lua = 7.9060667e-17
+ lub = -2.7964918e-26
+ luc = 5.5424848e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = -2.574678e-15
+ nsd = 1e+20
+ pbd = 0.75
+ pat = -1.0212358e-9
+ wvsat = -0.0027183681
+ pbs = 0.75
+ pk2 = 2.1304022e-16
+ aigbinv = 0.009974
+ wvth0 = -4.342128e-9
+ pu0 = -6.6237547e-17
+ vfbsdoff = 0.01
+ prt = 0
+ pua = -2.0419953e-23
+ pub = 1.469069e-32
+ puc = 1.2609666e-24
+ pud = 0
+ waigc = 6.0357037e-12
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 8.3453493e-9
+ ub1 = -1.1410668e-17
+ pvfbsdoff = 0
+ uc1 = 1.6197295e-9
+ keta = -0.31465021
+ lku0we = 1.8e-11
+ tpb = 0.0016
+ wa0 = -5.9482929e-8
+ epsrox = 3.9
+ ute = -1
+ wat = 0.022486376
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 1.7062889e-10
+ wlc = 0
+ wln = 1
+ wu0 = 1.3607209e-9
+ xgl = -8.2e-9
+ xgw = 0
+ wua = 3.3448805e-16
+ wub = -2.4882066e-25
+ wuc = -1.434288e-17
+ wud = 0
+ lketa = 1.5671934e-8
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ paramchk = 1
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 2.7213086e-10
+ xpart = 1
+ rdsmod = 0
+ kt1l = 0
+ igbmod = 1
+ egidl = 0.001
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ lint = 0
+ poxedge = 1
+ pbswgd = 0.8
+ pbswgs = 0.8
+ lkt1 = 1.2191281e-8
+ lkt2 = 2.350723e-9
+ lmax = 5.4e-8
+ lmin = 4.5e-8
+ ijthdfwd = 0.01
+ igcmod = 1
+ binunit = 2
+ lpe0 = 6.44e-8
+ lpeb = 0
+ minv = -0.33
+ lua1 = -3.7660644e-16
+ lub1 = 5.1040674e-25
+ luc1 = -7.3441373e-17
+ ndep = 1e+18
+ lwlc = 0
+ ijthdrev = 0.01
+ moin = 5.5538
+ nigc = 2.291
+ lpdiblc2 = 0
+ pvoff = 8.4992158e-17
+ cdscb = 0
+ cdscd = 0
+ pvsat = 1.1485877e-10
+ noff = 2.2684
+ wk2we = 0.0
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ pvth0 = -1.35778397e-16
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ permod = 1
+ drout = 0.56
+ paigc = -1.4334713e-18
+ voffl = 0
+ ntox = 1.0
+ pcit = -1.9199318e-17
+ pclm = 1.8533357
+ weta0 = -4.8723037e-9
+ wetab = 2.5894049e-9
+ lpclm = -6.4524768e-8
+ lkvth0we = 3e-12
+ phin = 0.15
+ voffcv = -0.125
+ wpemod = 1
+ pkt1 = -1.7583146000000001e-15
+ pkt2 = -1.1786798e-16
+ cgidl = 1
+ acnqsmod = 0
+ njtsswg = 6.489
+ rbdb = 50
+ pua1 = 1.8341764e-23
+ prwb = 0
+ pub1 = -1.3009877e-32
+ prwg = 0
+ puc1 = 9.9681375e-24
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ pbswd = 0.9
+ rbpb = 50
+ rbpd = 50
+ pbsws = 0.9
+ rbps = 50
+ rbodymod = 0
+ rbsb = 50
+ pvag = 2.1
+ ckappad = 0.6
+ ckappas = 0.6
+ rdsw = 200
+ pdiblc1 = 0
+ pdiblc2 = 0.0014658889
+ pdiblcb = 0
+ tpbswg = 0.001
+ pdits = 0
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ bigbacc = 0.0054401
+ ptvoff = -2.2999757e-17
+ pk2we = 0.0
+ wpdiblc2 = 1.4741467e-10
+ rshg = 14.1
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ waigsd = 1.9716411e-12
+ kvth0we = -0.00022
+ diomod = 1
+ tnoia = 0
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ pditsd = 0
+ pditsl = 0
+ vtsswgd = 1.1
+ peta0 = -1.1677509400000002e-17
+ vtsswgs = 1.1
+ cjswgd = 1.9113600000000002e-10
+ pku0we = 0.0
+ cjswgs = 1.9113600000000002e-10
+ petab = -2.558443e-17
+ wketa = 3.409679e-8
+ tpbsw = 0.0025
+ tnom = 25
+ cjswd = 5.3856e-11
+ cjsws = 5.3856e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ tvfbsdoff = 0.1
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ wkvth0we = 0.0
+ mjswgd = 0.95
+ mjswgs = 0.95
+ wtvfbsdoff = 0
+ tcjswg = 0.00128
+ trnqsmod = 0
+ ltvfbsdoff = 0
+ wags = 2.5054667e-7
+ wcit = 2.7838518e-10
+ scref = 1e-6
+ voff = -0.1005239
+ pigcd = 2.572
+ acde = 0.5
+ aigsd = 0.0063632396
+ nfactor = 1
+ rgatemod = 0
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ tnjtsswg = 1
+ vsat = 101849.16
+ wint = 0
+ lvoff = -3.8177557e-9
+ vth0 = -0.29714034
+ fprout = 200
+ wkt1 = 3.6711578e-8
+ wkt2 = 3.2153756e-9
+ wmax = 2.726e-7
+ xrcrg1 = 12
+ xrcrg2 = 1
+ aigc = 0.0068691843
+ wmin = 1.08e-7
+ lvsat = -0.00040815496000000005
+ lvth0 = -4.6946177e-9
+ ptvfbsdoff = 0
+ delta = 0.018814
+ laigc = -1.683393e-11
+ wtvoff = 5.2119196e-10
+ wua1 = -3.864028e-16
+ wub1 = 3.2172349e-25
+ wuc1 = -2.0479093e-16
+ rnoia = 0
+ rnoib = 0
+ a0 = 3.0243356
+ a1 = 0
+ a2 = 1
+ nigbacc = 10
+ b0 = 0
+ b1 = 0
+ at = -187272.02
+ cf = 8.17e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.021495622
+ k3 = -2.5823
+ em = 20000000.0
+ bigc = 0.0012521
+ ll = 0
+ lw = 0
+ u0 = -0.00038459259
+ w0 = 0
+ wwlc = 0
+ ua = -1.9655718e-9
+ ub = 1.5789686e-18
+ uc = -2.0243416e-10
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 3.4e-9
+ pketa = -2.1465872e-15
+ ngate = 1.7e+20
+ ngcon = 1
+ capmod = 2
+ wpclm = -1.4226467e-7
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ wku0we = 1.5e-11
+ xtid = 3
+ xtis = 3
+ gbmin = 1e-12
+ nigbinv = 2.171
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigc = 0.15259
+ jswgd = 3.69e-13
+ mobmod = 0
+ jswgs = 3.69e-13
+ )

.model pch_fs_40 pmos (
+ level = 54
+ fnoimod = 1
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ eigbinv = 1.1
+ laigsd = 6.1219753e-16
+ k2we = 5e-5
+ ijthsfwd = 0.01
+ tvoff = -0.00058332606
+ dsub = 0.5
+ dtox = 3.91e-10
+ xjbvd = 1
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ xjbvs = 1
+ lk2we = 0.0
+ eta0 = 0.11700471
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ etab = -0.15063456
+ ijthsrev = 0.01
+ cigbacc = 0.245
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = 1.2991389e-9
+ letab = 4.3496496e-9
+ tnoimod = 0
+ ppclm = -3.5647768e-15
+ dlcig = 2.5e-9
+ cigbinv = 0.006
+ bgidl = 1834800000.0
+ ppdiblc2 = 0
+ toxref = 3e-9
+ version = 4.5
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ tempmod = 0
+ ags = 1.2522222
+ cjd = 0.001421376
+ cit = -0.0077632099
+ cjs = 0.001421376
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 4.0349e-9
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ aigbacc = 0.012071
+ bigsd = 0.0003327
+ pkvth0we = 0.0
+ la0 = -3.4726683e-8
+ ltvoff = 1.026653e-10
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0.0023511307
+ kt1 = -0.31430817
+ kt2 = -0.12562663
+ lk2 = 6.6041473e-9
+ wvoff = 3.3909703e-9
+ llc = 0
+ lln = 1
+ lu0 = 5.2561728e-10
+ mjd = 0.335
+ mjs = 0.335
+ lua = 9.0470184e-17
+ lub = -1.3836274e-26
+ luc = 2.7216576e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 1.4761752e-15
+ nsd = 1e+20
+ pbd = 0.75
+ pat = -5.6834015e-11
+ wvsat = -0.010288162
+ pbs = 0.75
+ pk2 = -2.7720832e-16
+ aigbinv = 0.009974
+ wvth0 = -2.0296264100000005e-9
+ pu0 = -6.1923224e-17
+ vfbsdoff = 0.01
+ prt = 0
+ pua = -4.2432063e-24
+ pub = -6.6397485e-33
+ puc = -1.7176927e-24
+ pud = 0
+ waigc = -4.0606639e-11
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 2.1566906e-9
+ ub1 = -3.7269546e-18
+ pvfbsdoff = 0
+ uc1 = -1.7258848e-10
+ keta = 0.15497942
+ lku0we = 1.8e-11
+ tpb = 0.0016
+ wa0 = -1.421534e-7
+ epsrox = 3.9
+ ute = -1
+ wat = 0.002804707
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 1.0175701e-8
+ wlc = 0
+ wln = 1
+ wu0 = 1.2726735e-9
+ xgl = -8.2e-9
+ xgw = 0
+ wua = 4.3503521e-18
+ wub = 1.8649442e-25
+ wuc = 4.6446086e-17
+ wud = 0
+ lketa = -7.3399177e-9
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ paramchk = 1
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 5.2143803e-10
+ xpart = 1
+ rdsmod = 0
+ kt1l = 0
+ igbmod = 1
+ egidl = 0.001
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ lint = 0
+ poxedge = 1
+ pbswgd = 0.8
+ pbswgs = 0.8
+ lkt1 = 1.1563929e-9
+ lkt2 = 2.3369169e-9
+ lmax = 4.5e-8
+ lmin = 3.6e-8
+ ijthdfwd = 0.01
+ igcmod = 1
+ binunit = 2
+ lpe0 = 6.44e-8
+ lpeb = 0
+ minv = -0.33
+ lua1 = -7.3362164e-17
+ lub1 = 1.3390478e-25
+ luc1 = 1.4382206e-17
+ ndep = 1e+18
+ lwlc = 0
+ ijthdrev = 0.01
+ moin = 5.5538
+ nigc = 2.291
+ paigsd = -6.9790518e-23
+ lpdiblc2 = 0
+ pvoff = -7.4138231e-17
+ cdscb = 0
+ cdscd = 0
+ pvsat = 4.8577866e-10
+ noff = 2.2684
+ wk2we = 0.0
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ pvth0 = -2.4909097e-16
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ permod = 1
+ drout = 0.56
+ paigc = 8.520035e-19
+ voffl = 0
+ ntox = 1.0
+ pcit = -2.0087561999999998e-17
+ pclm = 0.41497396
+ weta0 = -1.499677e-9
+ wetab = 1.1541057e-8
+ lpclm = 5.9549575e-9
+ lkvth0we = 3e-12
+ phin = 0.15
+ voffcv = -0.125
+ wpemod = 1
+ pkt1 = -1.7540714e-15
+ pkt2 = -7.0509572e-16
+ cgidl = 1
+ acnqsmod = 0
+ njtsswg = 6.489
+ rbdb = 50
+ pua1 = 3.2441676e-23
+ prwb = 0
+ pub1 = -5.4663004e-32
+ prwg = 0
+ puc1 = -1.3788915e-24
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ pbswd = 0.9
+ rbpb = 50
+ rbpd = 50
+ pbsws = 0.9
+ rbps = 50
+ rbodymod = 0
+ rbsb = 50
+ pvag = 2.1
+ ckappad = 0.6
+ ckappas = 0.6
+ rdsw = 200
+ pdiblc1 = 0
+ pdiblc2 = 0.0014658889
+ pdiblcb = 0
+ tpbswg = 0.001
+ pdits = 0
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ bigbacc = 0.0054401
+ ptvoff = -3.9364956e-17
+ pk2we = 0.0
+ wpdiblc2 = 1.4741467e-10
+ rshg = 14.1
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ waigsd = 1.9730654e-12
+ kvth0we = -0.00022
+ diomod = 1
+ tnoia = 0
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ pditsd = 0
+ pditsl = 0
+ vtsswgd = 1.1
+ peta0 = -1.7693622e-16
+ vtsswgs = 1.1
+ cjswgd = 1.9113600000000002e-10
+ pku0we = 0.0
+ cjswgs = 1.9113600000000002e-10
+ petab = -4.6421536e-16
+ wketa = -5.7187654e-8
+ tpbsw = 0.0025
+ tnom = 25
+ cjswd = 5.3856e-11
+ cjsws = 5.3856e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ tvfbsdoff = 0.1
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ wkvth0we = 0.0
+ mjswgd = 0.95
+ mjswgs = 0.95
+ wtvfbsdoff = 0
+ tcjswg = 0.00128
+ trnqsmod = 0
+ ltvfbsdoff = 0
+ wags = 2.5054667e-7
+ wcit = 2.9651259e-10
+ scref = 1e-6
+ voff = -0.12231559
+ pigcd = 2.572
+ acde = 0.5
+ aigsd = 0.0063632271
+ nfactor = 1
+ rgatemod = 0
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ tnjtsswg = 1
+ vsat = 151791.98
+ wint = 0
+ lvoff = -2.7499629e-9
+ vth0 = -0.36108607000000004
+ fprout = 200
+ wkt1 = 3.6624982e-8
+ wkt2 = 1.5199615e-8
+ wmax = 2.726e-7
+ xrcrg1 = 12
+ xrcrg2 = 1
+ aigc = 0.0069354083
+ wmin = 1.08e-7
+ lvsat = -0.0028553534
+ lvth0 = -1.5612769e-9
+ ptvfbsdoff = 0
+ delta = 0.018814
+ laigc = -2.0078906e-11
+ wtvoff = 8.5517561e-10
+ wua1 = -6.7415611e-16
+ wub1 = 1.1717873e-24
+ wuc1 = 2.6781086e-17
+ rnoia = 0
+ rnoib = 0
+ a0 = 0.69140412
+ a1 = 0
+ a2 = 1
+ nigbacc = 10
+ b0 = 0
+ b1 = 0
+ at = -30917.36
+ cf = 8.17e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.06369048
+ k3 = -2.5823
+ em = 20000000.0
+ bigc = 0.0012521
+ ll = 0
+ lw = 0
+ u0 = -0.0026275802999999997
+ w0 = 0
+ wwlc = 0
+ ua = -2.1984191e-9
+ ub = 1.2906289e-18
+ uc = -1.4486626e-10
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 3.4e-9
+ pketa = 2.3263506e-15
+ ngate = 1.7e+20
+ ngcon = 1
+ capmod = 2
+ wpclm = 8.9861524e-8
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ wku0we = 1.5e-11
+ xtid = 3
+ xtis = 3
+ gbmin = 1e-12
+ nigbinv = 2.171
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigc = 0.15259
+ jswgd = 3.69e-13
+ mobmod = 0
+ jswgs = 3.69e-13
+ )

.model pch_sf_1 pmos (
+ level = 54
+ ppclm = 0
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ bigbacc = 0.0054401
+ wpdiblc2 = 0
+ tnom = 25
+ kvth0we = -0.00022
+ tvfbsdoff = 0.1
+ dmcgt = 0
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ tcjsw = 9.34e-5
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ toxref = 3e-9
+ bigsd = 0.0003327
+ wkvth0we = 0.0
+ wvoff = 0
+ trnqsmod = 0
+ voff = -0.11110337
+ acde = 0.5
+ wvsat = 0
+ wvfbsdoff = 0
+ wvth0 = 2.1600000000000004e-9
+ lvfbsdoff = 0
+ vsat = 120000
+ wint = 0
+ vth0 = -0.36113526999999995
+ ltvoff = 0
+ wmax = 0.00090001
+ aigc = 0.0068307507
+ wmin = 8.9974e-6
+ a0 = 2.531
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 72000
+ cf = 8.17e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.00077592763
+ k3 = -2.5823
+ em = 20000000.0
+ lketa = 0
+ ll = 0
+ lw = 0
+ u0 = 0.009715
+ w0 = 0
+ rgatemod = 0
+ ua = 1.297e-10
+ ub = 1.182572e-18
+ uc = 2.014e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xpart = 1
+ xw = 8.600000000000001e-9
+ nfactor = 1
+ tnjtsswg = 1
+ lku0we = 1.8e-11
+ bigc = 0.0012521
+ egidl = 0.001
+ wwlc = 0
+ epsrox = 3.9
+ cdsc = 0
+ rdsmod = 0
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ igbmod = 1
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigc = 0.15259
+ nigbacc = 10
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ pbswgd = 0.8
+ pbswgs = 0.8
+ igcmod = 1
+ nigbinv = 2.171
+ pvoff = -2e-17
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ cdscb = 0
+ cdscd = 0
+ pvsat = 0
+ wk2we = 0.0
+ pvth0 = 1.2e-16
+ drout = 0.56
+ k2we = 5e-5
+ dsub = 0.5
+ dtox = 3.91e-10
+ voffl = 0
+ fnoimod = 1
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ eigbinv = 1.1
+ weta0 = 2.2400000000000003e-10
+ permod = 1
+ lpclm = 0
+ eta0 = 0.1672
+ etab = -0.23
+ ijthsfwd = 0.01
+ cgidl = 1
+ voffcv = -0.125
+ wpemod = 1
+ ijthsrev = 0.01
+ pbswd = 0.9
+ pbsws = 0.9
+ cigbacc = 0.245
+ tnoimod = 0
+ pdits = 0
+ cigsd = 0.013281
+ cigbinv = 0.006
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ ppdiblc2 = 0
+ tpbswg = 0.001
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ version = 4.5
+ tempmod = 0
+ tnoia = 0
+ peta0 = 1.6e-17
+ ptvoff = 0
+ aigbacc = 0.012071
+ tpbsw = 0.0025
+ pkvth0we = 0.0
+ pvfbsdoff = 0
+ keta = -0.042350111
+ cjswd = 4.8144e-11
+ cjsws = 4.8144e-11
+ diomod = 1
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ pditsd = 0
+ pditsl = 0
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ cjswgd = 1.7086399999999997e-10
+ pku0we = 0.0
+ cjswgs = 1.7086399999999997e-10
+ lcit = -1.6e-11
+ aigbinv = 0.009974
+ vfbsdoff = 0.01
+ wtvfbsdoff = 0
+ kt1l = 0
+ lint = 6.5375218e-9
+ ltvfbsdoff = 0
+ mjswgd = 0.95
+ mjswgs = 0.95
+ lkt1 = 4.8e-10
+ paramchk = 1
+ lmax = 2.001e-5
+ lmin = 8.9991e-6
+ tcjswg = 0.00128
+ scref = 1e-6
+ lpe0 = 6.44e-8
+ lpeb = 0
+ pigcd = 2.572
+ aigsd = 0.0063636
+ minv = -0.33
+ lvoff = 0
+ poxedge = 1
+ ndep = 1e+18
+ lwlc = 0
+ ijthdfwd = 0.01
+ lvsat = -8.000000000000001e-6
+ moin = 5.5538
+ lvth0 = 2.4e-10
+ binunit = 2
+ ptvfbsdoff = 0
+ nigc = 2.291
+ delta = 0.018814
+ rnoia = 0
+ rnoib = 0
+ fprout = 200
+ noff = 2.2684
+ ags = 0.8379228
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ ijthdrev = 0.01
+ ngate = 1.7e+20
+ cjd = 0.001270624
+ cit = 5e-6
+ cjs = 0.001270624
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 1.0572421799999999e-8
+ ngcon = 1
+ k3b = 2.1176
+ wpclm = 0
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ lpdiblc2 = 0
+ ntox = 1.0
+ wtvoff = 0
+ pcit = 8.000000000000001e-19
+ pclm = 1.484
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ la0 = 0
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = -0.00064
+ kt1 = -0.17107633
+ lk2 = -3.2000000000000003e-10
+ kt2 = -0.04747
+ jtsswgd = 1.75e-7
+ phin = 0.15
+ llc = 0
+ jtsswgs = 1.75e-7
+ lln = 1
+ lu0 = 8e-13
+ mjd = 0.335
+ mjs = 0.335
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 0
+ capmod = 2
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ pk2 = 0
+ pkt1 = 4e-17
+ pu0 = 0
+ prt = 0
+ wku0we = 1.5e-11
+ pud = 0
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 1.1969344e-9
+ ub1 = -1.3666143e-18
+ uc1 = 6.873e-11
+ mobmod = 0
+ tpb = 0.0016
+ wa0 = 0
+ lkvth0we = 3e-12
+ ute = -1
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 0
+ wlc = 0
+ wln = 1
+ rbdb = 50
+ prwb = 0
+ wu0 = 0
+ prwg = 0
+ xgl = -8.2e-9
+ xgw = 0
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ rdsw = 200
+ tvoff = 0.0026155642
+ acnqsmod = 0
+ njtsswg = 6.489
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ xtsswgd = 0.32
+ rbodymod = 0
+ xtsswgs = 0.32
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.0026729629
+ ku0we = -0.0007
+ pdiblcb = 0
+ beta0 = 13.32
+ rshg = 14.1
+ leta0 = 4.8e-10
+ )

.model pch_sf_2 pmos (
+ level = 54
+ aigbinv = 0.009974
+ eta0 = 0.1672
+ tnoia = 0
+ etab = -0.23
+ ijthdfwd = 0.01
+ peta0 = 1.6e-17
+ toxref = 3e-9
+ pvfbsdoff = 0
+ tpbsw = 0.0025
+ cjswd = 4.8144e-11
+ cjsws = 4.8144e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ ijthdrev = 0.01
+ lpdiblc2 = 7.1311563e-9
+ poxedge = 1
+ ltvoff = -4.7585658e-10
+ binunit = 2
+ scref = 1e-6
+ pigcd = 2.572
+ aigsd = 0.0063636
+ lku0we = 1.8e-11
+ epsrox = 3.9
+ lkvth0we = 3e-12
+ lvoff = -8.0044387e-9
+ lvsat = -8.000000000000001e-6
+ rdsmod = 0
+ lvth0 = -4.8867661e-9
+ ags = 0.80385259
+ igbmod = 1
+ delta = 0.018814
+ laigc = -4.8397409e-11
+ cjd = 0.001270624
+ cit = 5e-6
+ cjs = 0.001270624
+ clc = 1e-7
+ cle = 0.6
+ acnqsmod = 0
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 1.0572421799999999e-8
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ k3b = 2.1176
+ rnoia = 0
+ rnoib = 0
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ keta = -0.040853613
+ pbswgd = 0.8
+ pbswgs = 0.8
+ rbodymod = 0
+ a0 = 2.5747309
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 72000
+ lags = 3.062912e-7
+ ngate = 1.7e+20
+ cf = 8.17e-11
+ igcmod = 1
+ la0 = -3.9314047e-7
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.0012551498
+ k3 = -2.5823
+ em = 20000000.0
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = -0.00064
+ ll = 0
+ lw = 0
+ kt1 = -0.16652617
+ kt2 = -0.046491549
+ lk2 = 3.988207500000001e-9
+ u0 = 0.0097148901
+ ngcon = 1
+ w0 = 0
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ ua = 1.4083134e-10
+ ub = 1.1675774e-18
+ uc = 1.8373185e-11
+ ud = 0
+ llc = 0
+ wpclm = 0
+ lln = 1
+ lcit = -1.6e-11
+ wl = 0
+ wr = 1
+ lu0 = 1.78779012e-12
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ mjd = 0.335
+ mjs = 0.335
+ lua = -1.0007073e-16
+ lub = 1.3480174e-25
+ luc = 1.5883665e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ kt1l = 0
+ njs = 1.02
+ pa0 = 0
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ pk2 = 0
+ gbmin = 1e-12
+ pu0 = 0
+ jswgd = 3.69e-13
+ prt = 0
+ jswgs = 3.69e-13
+ pud = 0
+ lint = 6.5375218e-9
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 1.1817684e-9
+ ub1 = -1.3634053e-18
+ uc1 = 6.7786161e-11
+ tpb = 0.0016
+ lkt1 = -4.0426013e-8
+ lkt2 = -8.7962711e-9
+ wa0 = 0
+ lmax = 8.9991e-6
+ ute = -1
+ lmin = 8.9908e-7
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 0
+ wlc = 0
+ wln = 1
+ wu0 = 0
+ xgl = -8.2e-9
+ xgw = 0
+ njtsswg = 6.489
+ lpe0 = 6.44e-8
+ wud = 0
+ wpdiblc2 = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ lpeb = 0
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ minv = -0.33
+ lua1 = 1.3634229e-16
+ lub1 = -2.8849398e-26
+ luc1 = 8.4851172e-18
+ permod = 1
+ ckappad = 0.6
+ ckappas = 0.6
+ ndep = 1e+18
+ pdiblc1 = 0
+ pdiblc2 = 0.0018797309
+ pdiblcb = 0
+ lwlc = 0
+ moin = 5.5538
+ nigc = 2.291
+ tvoff = 0.002668496
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ wkvth0we = 0.0
+ voffcv = -0.125
+ wpemod = 1
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ bigbacc = 0.0054401
+ trnqsmod = 0
+ ku0we = -0.0007
+ beta0 = 13.32
+ kvth0we = -0.00022
+ ntox = 1.0
+ pcit = 8.000000000000001e-19
+ pclm = 1.484
+ leta0 = 4.8e-10
+ lintnoi = -5e-9
+ ppclm = 0
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ phin = 0.15
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ pkt1 = 4e-17
+ rgatemod = 0
+ tpbswg = 0.001
+ tnjtsswg = 1
+ tvfbsdoff = 0.1
+ dmcgt = 0
+ rbdb = 50
+ tcjsw = 9.34e-5
+ prwb = 0
+ prwg = 0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ ptvoff = 0
+ wtvfbsdoff = 0
+ rdsw = 200
+ bigsd = 0.0003327
+ diomod = 1
+ ltvfbsdoff = 0
+ pditsd = 0
+ pditsl = 0
+ nfactor = 1
+ wvoff = 0
+ cjswgd = 1.7086399999999997e-10
+ pku0we = 0.0
+ cjswgs = 1.7086399999999997e-10
+ wvfbsdoff = 0
+ wvsat = 0
+ lvfbsdoff = 0
+ wvth0 = 2.1600000000000004e-9
+ rshg = 14.1
+ mjswgd = 0.95
+ mjswgs = 0.95
+ tcjswg = 0.00128
+ lketa = -1.3453518e-8
+ ptvfbsdoff = 0
+ nigbacc = 10
+ xpart = 1
+ tnom = 25
+ egidl = 0.001
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ ijthsfwd = 0.01
+ nigbinv = 2.171
+ fprout = 200
+ xrcrg1 = 12
+ xrcrg2 = 1
+ ijthsrev = 0.01
+ fnoimod = 1
+ voff = -0.110213
+ wtvoff = 0
+ acde = 0.5
+ eigbinv = 1.1
+ pvoff = -2e-17
+ vsat = 120000
+ wint = 0
+ vth0 = -0.36056499999999997
+ cdscb = 0
+ cdscd = 0
+ wmax = 0.00090001
+ pvsat = 0
+ aigc = 0.0068361342
+ wmin = 8.9974e-6
+ wk2we = 0.0
+ capmod = 2
+ pvth0 = 1.2e-16
+ drout = 0.56
+ wku0we = 1.5e-11
+ ppdiblc2 = 0
+ mobmod = 0
+ voffl = 0
+ bigc = 0.0012521
+ weta0 = 2.2400000000000003e-10
+ cigbacc = 0.245
+ wwlc = 0
+ lpclm = 0
+ cdsc = 0
+ tnoimod = 0
+ cgbo = 0
+ cgidl = 1
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigc = 0.15259
+ pkvth0we = 0.0
+ cigbinv = 0.006
+ pbswd = 0.9
+ pbsws = 0.9
+ vfbsdoff = 0.01
+ version = 4.5
+ tempmod = 0
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ pdits = 0
+ cigsd = 0.013281
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ dvt0w = 0
+ paramchk = 1
+ dvt1w = 0
+ dvt2w = 0
+ aigbacc = 0.012071
+ k2we = 5e-5
+ dsub = 0.5
+ dtox = 3.91e-10
+ pk2we = 0.0
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ )

.model pch_sf_3 pmos (
+ level = 54
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ nigbacc = 10
+ ijthsrev = 0.01
+ wvoff = 0
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ wvsat = 0
+ ntox = 1.0
+ wvth0 = 2.1600000000000004e-9
+ pcit = 8.000000000000001e-19
+ pclm = 1.484
+ ltvoff = -2.3123852e-10
+ nigbinv = 2.171
+ phin = 0.15
+ lketa = -1.5940244e-8
+ pkt1 = 4e-17
+ ppdiblc2 = 0
+ xpart = 1
+ lku0we = 1.8e-11
+ epsrox = 3.9
+ egidl = 0.001
+ rbdb = 50
+ fnoimod = 1
+ prwb = 0
+ prwg = 0
+ rdsmod = 0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ eigbinv = 1.1
+ igbmod = 1
+ rdsw = 200
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ pbswgd = 0.8
+ pbswgs = 0.8
+ pkvth0we = 0.0
+ igcmod = 1
+ vfbsdoff = 0.01
+ rshg = 14.1
+ cigbacc = 0.245
+ pvoff = -2e-17
+ cdscb = 0
+ cdscd = 0
+ pvsat = 0
+ tnoimod = 0
+ wk2we = 0.0
+ pvth0 = 1.2e-16
+ paramchk = 1
+ drout = 0.56
+ cigbinv = 0.006
+ voffl = 0
+ permod = 1
+ tnom = 25
+ weta0 = 2.2400000000000003e-10
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ a0 = 2.8917556
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ lpclm = 0
+ at = 72000
+ cf = 8.17e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = 0.0040664684
+ k3 = -2.5823
+ em = 20000000.0
+ ijthdfwd = 0.01
+ version = 4.5
+ ll = 0
+ lw = 0
+ u0 = 0.009946756
+ w0 = 0
+ ua = 1.1413788e-10
+ ub = 1.1978347e-18
+ uc = 4.3035111e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ tempmod = 0
+ cgidl = 1
+ voffcv = -0.125
+ wpemod = 1
+ aigbacc = 0.012071
+ ijthdrev = 0.01
+ pbswd = 0.9
+ pbsws = 0.9
+ voff = -0.10886793
+ lpdiblc2 = 1.7469722e-9
+ acde = 0.5
+ vsat = 120000
+ aigbinv = 0.009974
+ wint = 0
+ vth0 = -0.36318963
+ pdits = 0
+ cigsd = 0.013281
+ wmax = 0.00090001
+ aigc = 0.00683106
+ wmin = 8.9974e-6
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ wtvfbsdoff = 0
+ tpbswg = 0.001
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ ltvfbsdoff = 0
+ lkvth0we = 3e-12
+ bigc = 0.0012521
+ wwlc = 0
+ tnoia = 0
+ ptvoff = 0
+ poxedge = 1
+ cdsc = 0
+ peta0 = 1.6e-17
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ acnqsmod = 0
+ pvfbsdoff = 0
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigc = 0.15259
+ binunit = 2
+ diomod = 1
+ tpbsw = 0.0025
+ cjswd = 4.8144e-11
+ cjsws = 4.8144e-11
+ mjswd = 0.01
+ pditsd = 0
+ mjsws = 0.01
+ pditsl = 0
+ rbodymod = 0
+ agidl = 3.2166e-9
+ cjswgd = 1.7086399999999997e-10
+ pku0we = 0.0
+ cjswgs = 1.7086399999999997e-10
+ ptvfbsdoff = 0
+ dmcg = 3.1e-8
+ mjswgd = 0.95
+ dmci = 3.1e-8
+ dmdg = 0
+ mjswgs = 0.95
+ tcjswg = 0.00128
+ k2we = 5e-5
+ jtsswgd = 1.75e-7
+ scref = 1e-6
+ jtsswgs = 1.75e-7
+ wpdiblc2 = 0
+ dsub = 0.5
+ pigcd = 2.572
+ dtox = 3.91e-10
+ aigsd = 0.0063635603
+ ags = 0.82774541
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ lvoff = -9.201547e-9
+ cjd = 0.001270624
+ cit = -8.7888889e-5
+ cjs = 0.001270624
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 1.0572421799999999e-8
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ eta0 = 0.1672
+ etab = -0.23
+ lvsat = -8.000000000000001e-6
+ lvth0 = -2.5508401e-9
+ delta = 0.018814
+ laigc = -4.3881382e-11
+ la0 = -6.7529244e-7
+ fprout = 200
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = -0.00064
+ kt1 = -0.19559142
+ kt2 = -0.048919444
+ lk2 = -7.480327200000001e-10
+ llc = 0
+ lln = 1
+ lu0 = -2.0457243999999998e-10
+ rnoia = 0
+ rnoib = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ mjd = 0.335
+ mjs = 0.335
+ lua = -7.6313554e-17
+ lub = 1.0787275e-25
+ luc = -6.0654489e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ wkvth0we = 0.0
+ njs = 1.02
+ pa0 = 0
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ pk2 = 0
+ njtsswg = 6.489
+ pu0 = 0
+ prt = 0
+ pud = 0
+ ngate = 1.7e+20
+ trnqsmod = 0
+ wtvoff = 0
+ ngcon = 1
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 1.2804108e-9
+ ub1 = -1.1625424e-18
+ uc1 = 4.6637333e-11
+ wpclm = 0
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ tpb = 0.0016
+ wa0 = 0
+ ute = -1
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 0
+ ckappad = 0.6
+ ckappas = 0.6
+ gbmin = 1e-12
+ wlc = 0
+ wln = 1
+ wu0 = 0
+ xgl = -8.2e-9
+ xgw = 0
+ pdiblc1 = 0
+ pdiblc2 = 0.0079293759
+ wud = 0
+ jswgd = 3.69e-13
+ wwc = 0
+ jswgs = 3.69e-13
+ wwl = 0
+ wwn = 1
+ pdiblcb = 0
+ capmod = 2
+ wku0we = 1.5e-11
+ rgatemod = 0
+ mobmod = 0
+ tnjtsswg = 1
+ bigbacc = 0.0054401
+ kvth0we = -0.00022
+ lintnoi = -5e-9
+ tvoff = 0.0023936443
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ laigsd = 3.5374533e-14
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ keta = -0.03805954
+ lags = 2.8502658e-7
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 6.6671111e-11
+ ku0we = -0.0007
+ beta0 = 13.32
+ kt1l = 0
+ leta0 = 4.8e-10
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ ppclm = 0
+ lint = 6.5375218e-9
+ lkt1 = -1.4557938999999999e-8
+ lkt2 = -6.6354444e-9
+ dlcig = 2.5e-9
+ lmax = 8.9908e-7
+ bgidl = 1834800000.0
+ lmin = 4.4908e-7
+ lpe0 = 6.44e-8
+ lpeb = 0
+ tvfbsdoff = 0.1
+ minv = -0.33
+ lua1 = 4.8550568e-17
+ nfactor = 1
+ lub1 = -2.0761736e-25
+ luc1 = 2.7307573e-17
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ ndep = 1e+18
+ lwlc = 0
+ ijthsfwd = 0.01
+ moin = 5.5538
+ nigc = 2.291
+ toxref = 3e-9
+ bigsd = 0.0003327
+ )

.model pch_sf_4 pmos (
+ level = 54
+ aigc = 0.0067884199
+ wmin = 8.9974e-6
+ cjd = 0.001270624
+ cit = -0.00054497817
+ cjs = 0.001270624
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 1.38228675e-8
+ scref = 1e-6
+ k3b = 2.1176
+ rgatemod = 0
+ lku0we = 1.8e-11
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ pigcd = 2.572
+ tnjtsswg = 1
+ epsrox = 3.9
+ aigsd = 0.0063636407
+ njtsswg = 6.489
+ lvoff = -3.8830249e-9
+ bigc = 0.0012521
+ la0 = -4.3379389e-8
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = -0.00064
+ rdsmod = 0
+ kt1 = -0.2000222
+ kt2 = -0.054670852
+ lk2 = 1.0430220999999998e-9
+ wwlc = 0
+ llc = -1.18e-13
+ xtsswgd = 0.32
+ lln = 0.7
+ xtsswgs = 0.32
+ lu0 = -4.824545e-10
+ igbmod = 1
+ mjd = 0.335
+ mjs = 0.335
+ lua = -1.5477844e-16
+ lub = 5.0676856e-26
+ luc = -5.2541764e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ lvsat = -8.000000000000001e-6
+ njd = 1.02
+ njs = 1.02
+ pa0 = 0
+ lvth0 = 4.5804654e-9
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ ckappad = 0.6
+ pk2 = 0
+ ckappas = 0.6
+ cdsc = 0
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ pu0 = 0
+ pdiblc1 = 0
+ pdiblc2 = 0.013802718
+ delta = 0.018814
+ cgbo = 0
+ prt = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ pud = 0
+ pdiblcb = 0
+ xtid = 3
+ xtis = 3
+ laigc = -2.5119727e-11
+ pbswgd = 0.8
+ pbswgs = 0.8
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ rsh = 15.2
+ tcj = 0.000832
+ cigc = 0.15259
+ ua1 = 1.2553592e-9
+ ub1 = -1.2671808e-18
+ uc1 = 1.0455371e-10
+ rnoia = 0
+ rnoib = 0
+ tpb = 0.0016
+ wa0 = 0
+ igcmod = 1
+ ute = -1
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 0
+ wlc = 0
+ wln = 1
+ wu0 = 0
+ xgl = -8.2e-9
+ xgw = 0
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ ngate = 1.7e+20
+ ngcon = 1
+ wpclm = 0
+ bigbacc = 0.0054401
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ kvth0we = -0.00022
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ k2we = 5e-5
+ vtsswgs = 1.1
+ dsub = 0.5
+ dtox = 3.91e-10
+ permod = 1
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ eta0 = 0.1672
+ ijthsfwd = 0.01
+ etab = -0.23
+ tvoff = 0.002134918
+ voffcv = -0.125
+ wpemod = 1
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ ijthsrev = 0.01
+ wtvfbsdoff = 0
+ ku0we = -0.0007
+ beta0 = 13.32
+ nfactor = 1
+ leta0 = 4.8e-10
+ ltvfbsdoff = 0
+ ppclm = 0
+ a0 = 1.4555895
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 72000
+ cf = 8.17e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -4.1106394e-6
+ k3 = -2.5823
+ em = 20000000.0
+ ll = -1.18e-13
+ dlcig = 2.5e-9
+ lw = 0
+ u0 = 0.010578305999999999
+ w0 = 0
+ tpbswg = 0.001
+ ua = 2.9246716e-10
+ ub = 1.3278253e-18
+ uc = 4.119131e-11
+ ud = 0
+ bgidl = 1834800000.0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ ppdiblc2 = 0
+ tvfbsdoff = 0.1
+ nigbacc = 10
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ ptvoff = 0
+ ptvfbsdoff = 0
+ diomod = 1
+ nigbinv = 2.171
+ pkvth0we = 0.0
+ bigsd = 0.0003327
+ keta = -0.029364427
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.7086399999999997e-10
+ pku0we = 0.0
+ cjswgs = 1.7086399999999997e-10
+ wvoff = 0
+ lags = 5.4107004e-7
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 2.6779039e-10
+ vfbsdoff = 0.01
+ wvsat = 0
+ kt1l = 0
+ wvth0 = 2.1600000000000004e-9
+ mjswgd = 0.95
+ mjswgs = 0.95
+ fnoimod = 1
+ eigbinv = 1.1
+ tcjswg = 0.00128
+ lint = 9.7879675e-9
+ lkt1 = -1.2608393e-8
+ lkt2 = -4.1048253e-9
+ paramchk = 1
+ lmax = 4.4908e-7
+ lmin = 2.1577e-7
+ lketa = -1.9766093e-8
+ lpe0 = 6.44e-8
+ xpart = 1
+ lpeb = 0
+ minv = -0.33
+ lua1 = 5.9573279e-17
+ lub1 = -1.6157647e-25
+ egidl = 0.001
+ luc1 = 1.8243668e-18
+ ndep = 1e+18
+ lwlc = 0
+ ijthdfwd = 0.01
+ moin = 5.5538
+ cigbacc = 0.245
+ fprout = 200
+ nigc = 2.291
+ xrcrg1 = 12
+ xrcrg2 = 1
+ tnoimod = 0
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ ijthdrev = 0.01
+ cigbinv = 0.006
+ wtvoff = 0
+ lpdiblc2 = -8.3729822e-10
+ ntox = 1.0
+ pcit = 8.000000000000001e-19
+ pclm = 1.484
+ pvoff = -2e-17
+ capmod = 2
+ version = 4.5
+ cdscb = 0
+ cdscd = 0
+ pvsat = 0
+ phin = 0.15
+ wku0we = 1.5e-11
+ tempmod = 0
+ wk2we = 0.0
+ pvth0 = 1.2e-16
+ drout = 0.56
+ mobmod = 0
+ pkt1 = 4e-17
+ voffl = 0
+ aigbacc = 0.012071
+ lkvth0we = 3e-12
+ weta0 = 2.2400000000000003e-10
+ rbdb = 50
+ prwb = 0
+ prwg = 0
+ lpclm = 0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ rdsw = 200
+ aigbinv = 0.009974
+ cgidl = 1
+ acnqsmod = 0
+ rbodymod = 0
+ pbswd = 0.9
+ pbsws = 0.9
+ rshg = 14.1
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ pdits = 0
+ poxedge = 1
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ binunit = 2
+ wpdiblc2 = 0
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ tnom = 25
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ tnoia = 0
+ toxref = 3e-9
+ peta0 = 1.6e-17
+ pvfbsdoff = 0
+ tpbsw = 0.0025
+ wkvth0we = 0.0
+ cjswd = 4.8144e-11
+ cjsws = 4.8144e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ trnqsmod = 0
+ voff = -0.12095548
+ acde = 0.5
+ ltvoff = -1.1739897e-10
+ vsat = 120000
+ wint = 0
+ vth0 = -0.37939714999999996
+ wmax = 0.00090001
+ ags = 0.24582847
+ )

.model pch_sf_5 pmos (
+ level = 54
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ pbswgd = 0.8
+ pbswgs = 0.8
+ acnqsmod = 0
+ version = 4.5
+ tempmod = 0
+ igcmod = 1
+ keta = -0.12863898
+ rbodymod = 0
+ lags = 3.2185083e-8
+ aigbacc = 0.012071
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 5.994557300000001e-11
+ kt1l = 0
+ pvoff = -2e-17
+ cdscb = 0
+ cdscd = 0
+ lint = 9.7879675e-9
+ pvsat = 0.0
+ wk2we = 0.0
+ pvth0 = 1.2e-16
+ aigbinv = 0.009974
+ lkt1 = -4.2609966e-9
+ lkt2 = -5.2805906e-10
+ drout = 0.56
+ lmax = 2.1577e-7
+ lmin = 9e-8
+ wpdiblc2 = 0
+ lpe0 = 6.44e-8
+ permod = 1
+ lpeb = 0
+ voffl = 0
+ minv = -0.33
+ lua1 = -1.5051887e-16
+ lub1 = 1.742578e-25
+ luc1 = 7.2216103e-18
+ weta0 = 2.2400000000000003e-10
+ ndep = 1e+18
+ lpclm = -1.4239795e-8
+ wtvfbsdoff = 0
+ lwlc = 0
+ moin = 5.5538
+ cgidl = 1
+ voffcv = -0.125
+ wpemod = 1
+ nigc = 2.291
+ ltvfbsdoff = 0
+ poxedge = 1
+ wkvth0we = 0.0
+ noff = 2.2684
+ binunit = 2
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ pbswd = 0.9
+ pbsws = 0.9
+ trnqsmod = 0
+ ntox = 1.0
+ pcit = 8.000000000000001e-19
+ pclm = 1.5514872
+ pdits = 0
+ cigsd = 0.013281
+ phin = 0.15
+ tpbswg = 0.001
+ ptvfbsdoff = 0
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ pkt1 = 4e-17
+ rgatemod = 0
+ tnjtsswg = 1
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ ptvoff = 0
+ rbdb = 50
+ prwb = 0
+ prwg = 0
+ tnoia = 0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ pvfbsdoff = 0
+ rdsw = 200
+ peta0 = 1.6e-17
+ diomod = 1
+ tpbsw = 0.0025
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.7086399999999997e-10
+ pku0we = 0.0
+ cjswgs = 1.7086399999999997e-10
+ cjswd = 4.8144e-11
+ a0 = 1.4508547
+ a1 = 0
+ a2 = 1
+ cjsws = 4.8144e-11
+ b0 = 0
+ b1 = 0
+ mjswd = 0.01
+ at = 72000
+ cf = 8.17e-11
+ mjsws = 0.01
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.013949949
+ k3 = -2.5823
+ agidl = 3.2166e-9
+ em = 20000000.0
+ ll = -1.18e-13
+ lw = 0
+ u0 = 0.0091621197
+ w0 = 0
+ ua = -3.1871506e-10
+ ub = 1.6925299e-18
+ uc = 2.1642376e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ ags = 2.6576055
+ njtsswg = 6.489
+ mjswgd = 0.95
+ mjswgs = 0.95
+ cjd = 0.001270624
+ cit = 0.00044006838
+ cjs = 0.001270624
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ rshg = 14.1
+ bvs = 8.2
+ dlc = 1.38228675e-8
+ xtsswgd = 0.32
+ k3b = 2.1176
+ xtsswgs = 0.32
+ tcjswg = 0.00128
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.016932267
+ pdiblcb = 0
+ la0 = -4.2380342e-8
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = -0.00064
+ kt1 = -0.23958332
+ kt2 = -0.07162235
+ lk2 = 3.9855939000000005e-9
+ scref = 1e-6
+ llc = -1.18e-13
+ lln = 0.7
+ lu0 = -1.8363925e-10
+ mjd = 0.335
+ mjs = 0.335
+ lua = -2.581899e-17
+ lub = -2.6275812e-26
+ luc = -1.1293514e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ pigcd = 2.572
+ njd = 1.02
+ njs = 1.02
+ aigsd = 0.0063636407
+ pa0 = 0
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ pk2 = 0
+ pu0 = 0
+ prt = 0
+ pud = 0
+ tnom = 25
+ lvoff = -1.3382853e-9
+ rsh = 15.2
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ tcj = 0.000832
+ ua1 = 2.2510566e-9
+ ub1 = -2.8588123e-18
+ uc1 = 7.8974359e-11
+ bigbacc = 0.0054401
+ tpb = 0.0016
+ lvsat = 0.00083960684
+ ijthsfwd = 0.01
+ wa0 = 0
+ ute = -1
+ lvth0 = 5.4177832e-9
+ web = 6628.3
+ wec = -16935.0
+ fprout = 200
+ wk2 = 0
+ wlc = 0
+ wln = 1
+ wu0 = 0
+ xgl = -8.2e-9
+ xgw = 0
+ delta = 0.018814
+ wud = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ laigc = -2.0986759e-11
+ kvth0we = -0.00022
+ rnoia = 0
+ rnoib = 0
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ wtvoff = 0
+ vtsswgs = 1.1
+ ijthsrev = 0.01
+ ngate = 1.7e+20
+ wcit = 0.0
+ ngcon = 1
+ wpclm = 0
+ voff = -0.13301586
+ acde = 0.5
+ gbmin = 1e-12
+ capmod = 2
+ vsat = 115982.91
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ wint = 0
+ vth0 = -0.38336548
+ wku0we = 1.5e-11
+ wmax = 0.00090001
+ aigc = 0.0067688324
+ wmin = 8.9974e-6
+ mobmod = 0
+ ppdiblc2 = 0
+ bigc = 0.0012521
+ wwlc = 0
+ nfactor = 1
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ tvoff = 0.0018930751
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigc = 0.15259
+ xjbvd = 1
+ xjbvs = 1
+ pkvth0we = 0.0
+ lk2we = 0.0
+ vfbsdoff = 0.01
+ ku0we = -0.0007
+ nigbacc = 10
+ beta0 = 13.32
+ leta0 = 4.8e-10
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ ppclm = 0
+ paramchk = 1
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ nigbinv = 2.171
+ k2we = 5e-5
+ tvfbsdoff = 0.1
+ dsub = 0.5
+ dtox = 3.91e-10
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ eta0 = 0.1672
+ ijthdfwd = 0.01
+ etab = -0.23
+ toxref = 3e-9
+ fnoimod = 1
+ eigbinv = 1.1
+ bigsd = 0.0003327
+ ijthdrev = 0.01
+ wvfbsdoff = 0
+ wvoff = 0
+ lvfbsdoff = 0
+ ltvoff = -6.6370123e-11
+ lpdiblc2 = -1.4976331e-9
+ wvsat = 0.0
+ wvth0 = 2.1600000000000004e-9
+ cigbacc = 0.245
+ lku0we = 1.8e-11
+ lketa = 1.1808374e-9
+ tnoimod = 0
+ epsrox = 3.9
+ xpart = 1
+ rdsmod = 0
+ cigbinv = 0.006
+ egidl = 0.001
+ lkvth0we = 3e-12
+ igbmod = 1
+ )

.model pch_sf_6 pmos (
+ level = 54
+ wpclm = 0
+ vfbsdoff = 0.01
+ rshg = 14.1
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ nfactor = 1
+ wtvfbsdoff = 0
+ paramchk = 1
+ permod = 1
+ ltvfbsdoff = 0
+ tnom = 25
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ nigbacc = 10
+ ijthdfwd = 0.01
+ voffcv = -0.125
+ wpemod = 1
+ tvoff = 0.00091084129
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ nigbinv = 2.171
+ ptvfbsdoff = 0
+ ijthdrev = 0.01
+ wcit = 0.0
+ ku0we = -0.0007
+ lpdiblc2 = 0
+ voff = -0.11896044
+ beta0 = 13.32
+ acde = 0.5
+ leta0 = -6.341465e-10
+ letab = 2.0255694e-8
+ vsat = 185878.73
+ wint = 0
+ vth0 = -0.31330292
+ ppclm = 0
+ tpbswg = 0.001
+ wmax = 0.00090001
+ fnoimod = 1
+ aigc = 0.0067067782
+ wmin = 8.9974e-6
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ eigbinv = 1.1
+ tvfbsdoff = 0.1
+ ptvoff = 0
+ lkvth0we = 3e-12
+ bigc = 0.0012521
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ wwlc = 0
+ diomod = 1
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ acnqsmod = 0
+ pditsd = 0
+ pditsl = 0
+ cgsl = 3.0105e-11
+ cjswgd = 1.7086399999999997e-10
+ pku0we = 0.0
+ cgso = 2.6482e-11
+ cigbacc = 0.245
+ cjswgs = 1.7086399999999997e-10
+ cigc = 0.15259
+ bigsd = 0.0003327
+ rbodymod = 0
+ wvfbsdoff = 0
+ tnoimod = 0
+ lvfbsdoff = 0
+ wvoff = 0
+ mjswgd = 0.95
+ mjswgs = 0.95
+ wvsat = 0.0
+ cigbinv = 0.006
+ wvth0 = 2.1600000000000004e-9
+ tcjswg = 0.00128
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ version = 4.5
+ lketa = 8.4925319e-9
+ k2we = 5e-5
+ tempmod = 0
+ wpdiblc2 = 0
+ xpart = 1
+ dsub = 0.5
+ dtox = 3.91e-10
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ egidl = 0.001
+ a0 = 3.4166667
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 140456.11
+ cf = 8.17e-11
+ aigbacc = 0.012071
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.010241786
+ k3 = -2.5823
+ em = 20000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.0051538889
+ w0 = 0
+ ua = -1.1682959e-9
+ ub = 1.3034444e-18
+ uc = -8.7638e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ fprout = 200
+ eta0 = 0.17905262
+ etab = -0.44548611
+ xrcrg1 = 12
+ xrcrg2 = 1
+ aigbinv = 0.009974
+ wkvth0we = 0.0
+ wtvoff = 0
+ trnqsmod = 0
+ capmod = 2
+ pvoff = -2e-17
+ wku0we = 1.5e-11
+ cdscb = 0
+ cdscd = 0
+ mobmod = 0
+ pvsat = 0.0
+ wk2we = 0.0
+ pvth0 = 1.2e-16
+ drout = 0.56
+ poxedge = 1
+ rgatemod = 0
+ voffl = 0
+ tnjtsswg = 1
+ binunit = 2
+ weta0 = 2.2400000000000003e-10
+ lpclm = -9.8438889e-8
+ cgidl = 1
+ keta = -0.20642296
+ pbswd = 0.9
+ pbsws = 0.9
+ lags = -2.8753242e-8
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ lcit = 1.6951944e-10
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ kt1l = 0
+ pdits = 0
+ cigsd = 0.013281
+ lint = 0
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ lkt1 = -7.5119e-10
+ lkt2 = 1.5220167e-10
+ lmax = 9e-8
+ lmin = 5.4e-8
+ lpe0 = 6.44e-8
+ lpeb = 0
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ minv = -0.33
+ lua1 = -7.3062676e-18
+ lub1 = 1.0038041e-26
+ luc1 = 7.6176556e-18
+ ndep = 1e+18
+ toxref = 3e-9
+ njtsswg = 6.489
+ tnoia = 0
+ ijthsfwd = 0.01
+ lwlc = 0
+ pvfbsdoff = 0
+ moin = 5.5538
+ xtsswgd = 0.32
+ peta0 = 1.6e-17
+ xtsswgs = 0.32
+ nigc = 2.291
+ ckappad = 0.6
+ ckappas = 0.6
+ tpbsw = 0.0025
+ ags = 3.3058856
+ pdiblc1 = 0
+ pdiblc2 = 0.001
+ pdiblcb = 0
+ cjswd = 4.8144e-11
+ cjd = 0.001270624
+ cjsws = 4.8144e-11
+ cit = -0.00072561111
+ cjs = 0.001270624
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ dlc = 4.0349e-9
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ k3b = 2.1176
+ ijthsrev = 0.01
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ ltvoff = 2.5959859e-11
+ la0 = -2.2716667e-7
+ ntox = 1.0
+ pcit = 8.000000000000001e-19
+ jsd = 1.5e-7
+ pclm = 2.4472222
+ jss = 1.5e-7
+ lat = -0.0070748744
+ kt1 = -0.27692169
+ kt2 = -0.078859167
+ lk2 = 3.6370265999999995e-9
+ llc = 0
+ lln = 1
+ lu0 = 1.9313444000000001e-10
+ mjd = 0.335
+ bigbacc = 0.0054401
+ mjs = 0.335
+ lua = 5.4041604e-17
+ lub = 1.0298222e-26
+ luc = 9.143004e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 0
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ pk2 = 0
+ phin = 0.15
+ pu0 = 0
+ lku0we = 1.8e-11
+ prt = 0
+ pub = 0.0
+ pud = 0
+ kvth0we = -0.00022
+ epsrox = 3.9
+ ppdiblc2 = 0
+ rsh = 15.2
+ scref = 1e-6
+ pkt1 = 4e-17
+ tcj = 0.000832
+ ua1 = 7.2751825e-10
+ ub1 = -1.1117937e-18
+ uc1 = 7.4761111e-11
+ tpb = 0.0016
+ pigcd = 2.572
+ lintnoi = -5e-9
+ wa0 = 0
+ aigsd = 0.0063636407
+ ute = -1
+ web = 6628.3
+ wec = -16935.0
+ bigbinv = 0.00149
+ wk2 = 0
+ rdsmod = 0
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ wlc = 0
+ wln = 1
+ wu0 = 0
+ xgl = -8.2e-9
+ xgw = 0
+ wub = 0.0
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ igbmod = 1
+ lvoff = -2.6594942e-9
+ rbdb = 50
+ prwb = 0
+ prwg = 0
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ rbpb = 50
+ rbpd = 50
+ lvsat = -0.0057306009000000005
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ lvth0 = -1.168097e-9
+ pbswgd = 0.8
+ pbswgs = 0.8
+ rdsw = 200
+ delta = 0.018814
+ laigc = -1.5153664e-11
+ igcmod = 1
+ rnoia = 0
+ rnoib = 0
+ pkvth0we = 0.0
+ ngate = 1.7e+20
+ ngcon = 1
+ )

.model pch_sf_7 pmos (
+ level = 54
+ voffl = 0
+ dsub = 0.5
+ dtox = 3.91e-10
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ weta0 = 2.2400000000000003e-10
+ ptvfbsdoff = 0
+ lpclm = -4.4240467e-8
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ eta0 = 0.18948293
+ ijthsfwd = 0.01
+ voffcv = -0.125
+ wpemod = 1
+ etab = -0.27185615
+ cgidl = 1
+ ijthsrev = 0.01
+ pbswd = 0.9
+ pbsws = 0.9
+ njtsswg = 6.489
+ tpbswg = 0.001
+ pdits = 0
+ cigsd = 0.013281
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ ppdiblc2 = 0
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.001
+ pdiblcb = 0
+ pk2we = 0.0
+ ptvoff = 0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ ags = 2.81014
+ pvfbsdoff = 0
+ tnoia = 0
+ diomod = 1
+ cjd = 0.001270624
+ cit = -0.0030912222
+ cjs = 0.001270624
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 4.0349e-9
+ peta0 = 1.6e-17
+ k3b = 2.1176
+ pditsd = 0
+ pditsl = 0
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ bigbacc = 0.0054401
+ dwj = 0
+ cjswgd = 1.7086399999999997e-10
+ pku0we = 0.0
+ cjswgs = 1.7086399999999997e-10
+ tpbsw = 0.0025
+ pkvth0we = 0.0
+ keta = 0.048888889
+ cjswd = 4.8144e-11
+ kvth0we = -0.00022
+ cjsws = 4.8144e-11
+ la0 = -1.5788889e-7
+ jsd = 1.5e-7
+ mjswd = 0.01
+ jss = 1.5e-7
+ lat = 0.0036261578
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ kt1 = -0.090229195
+ kt2 = -0.087042222
+ lk2 = 4.0153879e-9
+ llc = 0
+ lln = 1
+ lu0 = -7.1828889e-11
+ mjd = 0.335
+ mjs = 0.335
+ lua = -4.5270917e-17
+ lub = -1.9748742e-26
+ luc = -2.161341e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ lintnoi = -5e-9
+ njd = 1.02
+ mjswgd = 0.95
+ njs = 1.02
+ mjswgs = 0.95
+ pa0 = 0
+ bigbinv = 0.00149
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ jswd = 3.69e-13
+ vtsswgd = 1.1
+ pk2 = 0
+ jsws = 3.69e-13
+ vtsswgs = 1.1
+ vfbsdoff = 0.01
+ lcit = 3.0672489e-10
+ pu0 = 0
+ tcjswg = 0.00128
+ prt = 0
+ pub = 0.0
+ pud = 0
+ kt1l = 0
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 1.0031266e-9
+ ub1 = -2.5489021e-18
+ uc1 = 1.9738889e-10
+ tpb = 0.0016
+ wa0 = 0
+ ute = -1
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 0
+ lint = 0
+ wlc = 0
+ wln = 1
+ wu0 = 0
+ xgl = -8.2e-9
+ xgw = 0
+ paramchk = 1
+ wub = 0.0
+ wud = 0
+ wwc = 0
+ lkt1 = -1.1579355e-8
+ lkt2 = 6.2681889e-10
+ wwl = 0
+ wwn = 1
+ lmax = 5.4e-8
+ lmin = 4.5e-8
+ scref = 1e-6
+ lpe0 = 6.44e-8
+ lpeb = 0
+ pigcd = 2.572
+ aigsd = 0.0063636407
+ minv = -0.33
+ lvoff = -4.1866651e-9
+ lua1 = -2.3291554e-17
+ lub1 = 9.339033e-26
+ luc1 = 5.0524444e-19
+ fprout = 200
+ ndep = 1e+18
+ lvsat = -0.00014810428
+ ijthdfwd = 0.01
+ xrcrg1 = 12
+ xrcrg2 = 1
+ lwlc = 0
+ lvth0 = -2.0766339e-9
+ moin = 5.5538
+ delta = 0.018814
+ laigc = -9.9932362e-12
+ nigc = 2.291
+ nfactor = 1
+ rnoia = 0
+ rnoib = 0
+ wtvoff = 0
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ ijthdrev = 0.01
+ ngate = 1.7e+20
+ ngcon = 1
+ wpclm = 0
+ lpdiblc2 = 0
+ capmod = 2
+ ntox = 1.0
+ pcit = 8.000000000000001e-19
+ wku0we = 1.5e-11
+ pclm = 1.5127667
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ nigbacc = 10
+ a0 = 2.2222222
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = -44044.444
+ mobmod = 0
+ cf = 8.17e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.016765256
+ k3 = -2.5823
+ em = 20000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.0097222222
+ w0 = 0
+ ua = 5.4398899e-10
+ ub = 1.8214956e-18
+ uc = 4.42645e-10
+ ud = 0
+ phin = 0.15
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ pkt1 = 4e-17
+ nigbinv = 2.171
+ lkvth0we = 3e-12
+ rbdb = 50
+ prwb = 0
+ prwg = 0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ rdsw = 200
+ tvoff = 0.0051729841
+ acnqsmod = 0
+ fnoimod = 1
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ eigbinv = 1.1
+ rbodymod = 0
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = -1.2391043e-9
+ rshg = 14.1
+ letab = 1.0185157e-8
+ ppclm = 0
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ tvfbsdoff = 0.1
+ cigbacc = 0.245
+ wpdiblc2 = 0
+ tnoimod = 0
+ tnom = 25
+ dmcgt = 0
+ toxref = 3e-9
+ tcjsw = 9.34e-5
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ cigbinv = 0.006
+ bigsd = 0.0003327
+ wkvth0we = 0.0
+ version = 4.5
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ tempmod = 0
+ ltvoff = -2.2124443e-10
+ wvoff = 0
+ wcit = 0.0
+ trnqsmod = 0
+ voff = -0.092629909
+ wvsat = 0.0
+ acde = 0.5
+ wvth0 = 2.1600000000000004e-9
+ aigbacc = 0.012071
+ vsat = 89628.791
+ wint = 0
+ vth0 = -0.29763849
+ lku0we = 1.8e-11
+ wmax = 0.00090001
+ aigc = 0.0066178053
+ wmin = 8.9974e-6
+ epsrox = 3.9
+ lketa = -6.3155556e-9
+ rgatemod = 0
+ xpart = 1
+ aigbinv = 0.009974
+ tnjtsswg = 1
+ rdsmod = 0
+ igbmod = 1
+ egidl = 0.001
+ bigc = 0.0012521
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ wwlc = 0
+ pbswgd = 0.8
+ pbswgs = 0.8
+ cdsc = 0
+ cgbo = 0
+ igcmod = 1
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigc = 0.15259
+ wtvfbsdoff = 0
+ poxedge = 1
+ binunit = 2
+ ltvfbsdoff = 0
+ pvoff = -2e-17
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ cdscb = 0
+ cdscd = 0
+ pvsat = 0.0
+ wk2we = 0.0
+ pvth0 = 1.2e-16
+ drout = 0.56
+ permod = 1
+ k2we = 5e-5
+ )

.model pch_sf_8 pmos (
+ level = 54
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ wkvth0we = 0.0
+ cigbacc = 0.245
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ trnqsmod = 0
+ ku0we = -0.0007
+ tnoimod = 0
+ beta0 = 13.32
+ leta0 = 2.6123128e-9
+ ntox = 1.0
+ letab = 3.9337702e-9
+ pcit = 8.000000000000001e-19
+ pclm = 1.0208333
+ tpbswg = 0.001
+ cigbinv = 0.006
+ ppclm = 0
+ phin = 0.15
+ dlcig = 2.5e-9
+ tvfbsdoff = 0.1
+ bgidl = 1834800000.0
+ pkt1 = 4e-17
+ rgatemod = 0
+ ptvoff = 0
+ tnjtsswg = 1
+ version = 4.5
+ tempmod = 0
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ diomod = 1
+ rbdb = 50
+ prwb = 0
+ prwg = 0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ aigbacc = 0.012071
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.7086399999999997e-10
+ pku0we = 0.0
+ cjswgs = 1.7086399999999997e-10
+ rdsw = 200
+ bigsd = 0.0003327
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ mjswgd = 0.95
+ mjswgs = 0.95
+ wvoff = 0
+ aigbinv = 0.009974
+ tcjswg = 0.00128
+ wvsat = 0.0
+ wvth0 = 2.1600000000000004e-9
+ rshg = 14.1
+ lketa = 8.0381778e-9
+ xpart = 1
+ poxedge = 1
+ egidl = 0.001
+ tnom = 25
+ fprout = 200
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ xrcrg1 = 12
+ xrcrg2 = 1
+ binunit = 2
+ ijthsfwd = 0.01
+ wtvoff = 0
+ ijthsrev = 0.01
+ wcit = 0.0
+ capmod = 2
+ voff = -0.10032114
+ wku0we = 1.5e-11
+ acde = 0.5
+ pvoff = -2e-17
+ mobmod = 0
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ vsat = 122520.32
+ wint = 0
+ vth0 = -0.34438557
+ cdscb = 0
+ cdscd = 0
+ wkt1 = 0.0
+ pvsat = 0.0
+ wmax = 0.00090001
+ wk2we = 0.0
+ pvth0 = 1.2e-16
+ aigc = 0.0065563017
+ wmin = 8.9974e-6
+ drout = 0.56
+ ppdiblc2 = 0
+ voffl = 0
+ weta0 = 2.2400000000000003e-10
+ wetab = 0
+ bigc = 0.0012521
+ wwlc = 0
+ lpclm = -2.0135733e-8
+ laigsd = -2.1777787e-18
+ cdsc = 0
+ cgidl = 1
+ njtsswg = 6.489
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigc = 0.15259
+ a0 = -0.19555556
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ xtsswgd = 0.32
+ pkvth0we = 0.0
+ xtsswgs = 0.32
+ at = 76220.0
+ cf = 8.17e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.012217534
+ k3 = -2.5823
+ em = 20000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.0052177778
+ w0 = 0
+ ua = -1.1794951e-9
+ ub = 1.5005044e-18
+ uc = 5.0701667e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.001
+ pbswd = 0.9
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ pbsws = 0.9
+ pdiblcb = 0
+ vfbsdoff = 0.01
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ pdits = 0
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ paramchk = 1
+ bigbacc = 0.0054401
+ k2we = 5e-5
+ ags = 1.0774289
+ dsub = 0.5
+ kvth0we = -0.00022
+ dtox = 3.91e-10
+ cjd = 0.001270624
+ cit = -0.00097166667
+ pk2we = 0.0
+ cjs = 0.001270624
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ dlc = 4.0349e-9
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ k3b = 2.1176
+ toxref = 3e-9
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ pvfbsdoff = 0
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ tnoia = 0
+ ijthdfwd = 0.01
+ eta0 = 0.11088258
+ etab = -0.14427684
+ la0 = -3.9417778e-8
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = -0.0022668000000000002
+ kt1 = -0.30391077
+ kt2 = -0.08425
+ lk2 = 3.7925495e-9
+ peta0 = 1.6e-17
+ llc = 0
+ lln = 1
+ lu0 = 1.4888889e-10
+ petab = 0
+ mjd = 0.335
+ mjs = 0.335
+ lua = 3.9179804e-17
+ lub = -4.0201778e-27
+ luc = -2.4081867e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 0
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0.0
+ pbs = 0.75
+ tpbsw = 0.0025
+ pk2 = 0
+ pu0 = 0
+ prt = 0
+ pub = 0.0
+ pud = 0
+ cjswd = 4.8144e-11
+ cjsws = 4.8144e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ ltvoff = -2.4936809e-11
+ agidl = 3.2166e-9
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 1.4917512e-9
+ ub1 = -1.5908843e-18
+ uc1 = 1.6325556e-10
+ ijthdrev = 0.01
+ tpb = 0.0016
+ wa0 = 0
+ ute = -1
+ wat = 0.0
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 0
+ wlc = 0
+ wln = 1
+ lpdiblc2 = 0
+ wu0 = 0
+ xgl = -8.2e-9
+ xgw = 0
+ wub = 0.0
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ lku0we = 1.8e-11
+ epsrox = 3.9
+ nfactor = 1
+ scref = 1e-6
+ rdsmod = 0
+ pigcd = 2.572
+ aigsd = 0.0063636407
+ igbmod = 1
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ wtvfbsdoff = 0
+ lvoff = -3.8097951e-9
+ lkvth0we = 3e-12
+ pbswgd = 0.8
+ pbswgs = 0.8
+ lvsat = -0.0017597894
+ lvth0 = 2.13972942e-10
+ igcmod = 1
+ ltvfbsdoff = 0
+ delta = 0.018814
+ nigbacc = 10
+ laigc = -6.97956e-12
+ acnqsmod = 0
+ rnoia = 0
+ rnoib = 0
+ keta = -0.24404444
+ rbodymod = 0
+ ngate = 1.7e+20
+ lags = 8.4902844e-8
+ ngcon = 1
+ nigbinv = 2.171
+ wpclm = 0
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 2.0286667e-10
+ kt1l = 0
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ ptvfbsdoff = 0
+ lint = 0
+ permod = 1
+ lkt1 = -1.1089574e-9
+ lkt2 = 4.9e-10
+ lmax = 4.5e-8
+ lmin = 3.6e-8
+ fnoimod = 1
+ wpdiblc2 = 0
+ lpe0 = 6.44e-8
+ lpeb = 0
+ eigbinv = 1.1
+ minv = -0.33
+ lua1 = -4.7234158e-17
+ lub1 = 4.6447457e-26
+ luc1 = 2.1777778e-18
+ voffcv = -0.125
+ wpemod = 1
+ ndep = 1e+18
+ lwlc = 0
+ moin = 5.5538
+ tvoff = 0.0011667062
+ nigc = 2.291
+ )

.model pch_sf_9 pmos (
+ level = 54
+ vtsswgs = 1.1
+ ags = 0.82538676
+ vsat = 121084.96
+ wint = 0
+ vth0 = -0.36147733
+ pdits = 0
+ cjd = 0.001270624
+ cit = 5e-6
+ cjs = 0.001270624
+ clc = 1e-7
+ cle = 0.6
+ cigsd = 0.013281
+ bvd = 8.2
+ bvs = 8.2
+ wkt1 = -1.0361455e-8
+ wkt2 = -3.8769913e-9
+ dlc = 1.0572421799999999e-8
+ wmax = 8.9974e-6
+ dvt0w = 0
+ k3b = 2.1176
+ dvt1w = 0
+ aigc = 0.0068303602
+ dvt2w = 0
+ wmin = 8.974e-7
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ ptvoff = 0
+ waigsd = 1.9139418e-12
+ la0 = 0
+ pk2we = 0.0
+ jsd = 1.5e-7
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ jss = 1.5e-7
+ lat = -0.00064
+ wua1 = -3.2799159e-16
+ kt1 = -0.16992583
+ lk2 = -3.2000000000000003e-10
+ kt2 = -0.04703951
+ wub1 = 5.9231251e-25
+ wuc1 = -8.7396626e-17
+ llc = 0
+ lln = 1
+ lu0 = 8e-13
+ mjd = 0.335
+ mjs = 0.335
+ lkvth0we = 3e-12
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ diomod = 1
+ pvfbsdoff = 0
+ njd = 1.02
+ bigc = 0.0012521
+ njs = 1.02
+ wute = -7.8572347e-8
+ pa0 = 0
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ wwlc = 0
+ pk2 = 0
+ tnoia = 0
+ pu0 = 0
+ pditsd = 0
+ pditsl = 0
+ prt = 0
+ pud = 0
+ cjswgd = 1.7086399999999997e-10
+ pku0we = 0.0
+ cjswgs = 1.7086399999999997e-10
+ rsh = 15.2
+ tcj = 0.000832
+ peta0 = 1.6e-17
+ cdsc = 0
+ ua1 = 1.2333536e-9
+ ub1 = -1.432383e-18
+ uc1 = 7.8434267e-11
+ cgbo = 0
+ tpb = 0.0016
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ acnqsmod = 0
+ xtid = 3
+ xtis = 3
+ wketa = 2.2362589e-8
+ wa0 = 3.3745816e-7
+ ute = -0.99127556
+ web = 6628.3
+ wec = -16935.0
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ wk2 = -2.287053e-9
+ tpbsw = 0.0025
+ cigc = 0.15259
+ wlc = 0
+ wln = 1
+ wu0 = -8.6631049e-11
+ xgl = -8.2e-9
+ xgw = 0
+ wua = -1.124189e-16
+ wub = -6.7100784e-26
+ wuc = -2.319496e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ cjswd = 4.8144e-11
+ nfactor = 1
+ cjsws = 4.8144e-11
+ mjswd = 0.01
+ mjswgd = 0.95
+ mjsws = 0.01
+ mjswgs = 0.95
+ agidl = 3.2166e-9
+ rbodymod = 0
+ tcjswg = 0.00128
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ nigbacc = 10
+ scref = 1e-6
+ k2we = 5e-5
+ wpdiblc2 = 3.6469361e-10
+ pigcd = 2.572
+ dsub = 0.5
+ aigsd = 0.0063633875
+ dtox = 3.91e-10
+ fprout = 200
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ lvoff = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ nigbinv = 2.171
+ lvsat = -8.000000000000001e-6
+ eta0 = 0.16744607
+ etab = -0.23671111
+ lvth0 = 2.4e-10
+ delta = 0.018814
+ wtvoff = -9.8925647e-11
+ rnoia = 0
+ rnoib = 0
+ wkvth0we = 0.0
+ fnoimod = 1
+ ngate = 1.7e+20
+ capmod = 2
+ trnqsmod = 0
+ eigbinv = 1.1
+ ngcon = 1
+ wpclm = -3.01194e-7
+ wku0we = 1.5e-11
+ mobmod = 0
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ rgatemod = 0
+ tnjtsswg = 1
+ cigbacc = 0.245
+ tnoimod = 0
+ tvoff = 0.0026265487
+ cigbinv = 0.006
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ keta = -0.044833188
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ version = 4.5
+ jswd = 3.69e-13
+ ku0we = -0.0007
+ jsws = 3.69e-13
+ lcit = -1.6e-11
+ tempmod = 0
+ beta0 = 13.32
+ leta0 = 4.8e-10
+ kt1l = 0
+ ppclm = 0
+ aigbacc = 0.012071
+ lint = 6.5375218e-9
+ tvfbsdoff = 0.1
+ dlcig = 2.5e-9
+ lkt1 = 4.8e-10
+ bgidl = 1834800000.0
+ lmax = 2.001e-5
+ lmin = 8.9991e-6
+ lpe0 = 6.44e-8
+ lpeb = 0
+ a0 = 2.4935296
+ a1 = 0
+ a2 = 1
+ toxref = 3e-9
+ b0 = 0
+ b1 = 0
+ at = 72000
+ cf = 8.17e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.00052197993
+ k3 = -2.5823
+ em = 20000000.0
+ aigbinv = 0.009974
+ minv = -0.33
+ ll = 0
+ lw = 0
+ u0 = 0.009724619299999999
+ w0 = 0
+ ua = 1.4218267e-10
+ ub = 1.1900227e-18
+ uc = 2.2715501e-11
+ ud = 0
+ dmcgt = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ tcjsw = 9.34e-5
+ ndep = 1e+18
+ ijthsfwd = 0.01
+ lwlc = 0
+ moin = 5.5538
+ nigc = 2.291
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ bigsd = 0.0003327
+ ltvoff = 0
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ ijthsrev = 0.01
+ wvoff = 5.5905393e-9
+ poxedge = 1
+ wvsat = -0.0097711764
+ wvth0 = 5.240586000000001e-9
+ ntox = 1.0
+ pcit = 8.000000000000001e-19
+ pclm = 1.5174437
+ binunit = 2
+ lku0we = 1.8e-11
+ wtvfbsdoff = 0
+ waigc = 3.5172206e-12
+ epsrox = 3.9
+ phin = 0.15
+ lketa = 0
+ rdsmod = 0
+ ltvfbsdoff = 0
+ ppdiblc2 = 0
+ pkt1 = 4e-17
+ xpart = 1
+ igbmod = 1
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ egidl = 0.001
+ pbswgd = 0.8
+ pbswgs = 0.8
+ rbdb = 50
+ prwb = 0
+ prwg = 0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ igcmod = 1
+ rbsb = 50
+ pvag = 2.1
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ rdsw = 200
+ ptvfbsdoff = 0
+ pkvth0we = 0.0
+ vfbsdoff = 0.01
+ rshg = 14.1
+ pvoff = -2e-17
+ cdscb = 0
+ cdscd = 0
+ permod = 1
+ pvsat = 0
+ wk2we = 0.0
+ pvth0 = 1.2e-16
+ paramchk = 1
+ njtsswg = 6.489
+ drout = 0.56
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ voffl = 0
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.0026324684
+ weta0 = -1.9921431e-9
+ tnom = 25
+ pdiblcb = 0
+ wetab = 6.0440267e-8
+ voffcv = -0.125
+ wpemod = 1
+ lpclm = 0
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ ijthdfwd = 0.01
+ cgidl = 1
+ bigbacc = 0.0054401
+ wags = 1.128996e-7
+ ijthdrev = 0.01
+ pbswd = 0.9
+ pbsws = 0.9
+ kvth0we = -0.00022
+ lpdiblc2 = 0
+ voff = -0.11172412
+ tpbswg = 0.001
+ acde = 0.5
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ )

.model pch_sf_10 pmos (
+ level = 54
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ lags = 3.1017116e-7
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = -1.6e-11
+ nfactor = 1
+ kt1l = 0
+ paramchk = 1
+ scref = 1e-6
+ pigcd = 2.572
+ aigsd = 0.0063633879
+ lint = 6.5375218e-9
+ lkt1 = -4.1427451999999996e-8
+ lkt2 = -8.3161855e-9
+ lmax = 8.9991e-6
+ lvoff = -7.1040424e-9
+ lmin = 8.9908e-7
+ lpe0 = 6.44e-8
+ lpeb = 0
+ lvsat = -8.000000000000001e-6
+ lvth0 = -4.2417588e-9
+ ijthdfwd = 0.01
+ toxref = 3e-9
+ nigbacc = 10
+ minv = -0.33
+ delta = 0.018814
+ lua1 = 2.9697696e-17
+ lub1 = 1.2607181e-25
+ luc1 = -4.744495e-18
+ laigc = -4.752933e-11
+ wtvfbsdoff = 0
+ ndep = 1e+18
+ rnoia = 0
+ rnoib = 0
+ lute = -8.6179201e-9
+ lwlc = 0
+ tvfbsdoff = 0.1
+ moin = 5.5538
+ ltvfbsdoff = 0
+ pketa = -2.2807538e-14
+ nigc = 2.291
+ ngate = 1.7e+20
+ ijthdrev = 0.01
+ nigbinv = 2.171
+ ngcon = 1
+ wpclm = -3.01194e-7
+ lpdiblc2 = 7.3300428e-9
+ ltvoff = -4.2514859e-10
+ gbmin = 1e-12
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ pags = -3.4942959e-14
+ ntox = 1.0
+ pcit = 8.000000000000001e-19
+ pclm = 1.5174437
+ fnoimod = 1
+ wvfbsdoff = 0
+ lku0we = 1.8e-11
+ ptvfbsdoff = 0
+ eigbinv = 1.1
+ lvfbsdoff = 0
+ epsrox = 3.9
+ phin = 0.15
+ lkvth0we = 3e-12
+ pkt1 = 9.058958600000001e-15
+ pkt2 = -4.3236504e-15
+ rdsmod = 0
+ igbmod = 1
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ tvoff = 0.0026738399
+ pbswgd = 0.8
+ acnqsmod = 0
+ pbswgs = 0.8
+ rbdb = 50
+ pua1 = 9.6044121e-22
+ prwb = 0
+ pub1 = -1.3952204e-30
+ prwg = 0
+ puc1 = 1.1914589e-22
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ pute = 7.7612988e-14
+ igcmod = 1
+ cigbacc = 0.245
+ rdsw = 200
+ rbodymod = 0
+ tnoimod = 0
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = 4.8e-10
+ cigbinv = 0.006
+ ppclm = 0
+ paigsd = 3.3403436e-20
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ rshg = 14.1
+ version = 4.5
+ wpdiblc2 = 5.6393415e-10
+ permod = 1
+ tempmod = 0
+ ags = 0.79088496
+ dmcgt = 0
+ cjd = 0.001270624
+ cit = 5e-6
+ cjs = 0.001270624
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ tcjsw = 9.34e-5
+ dlc = 1.0572421799999999e-8
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ aigbacc = 0.012071
+ tnom = 25
+ la0 = -3.6651331e-7
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ jsd = 1.5e-7
+ voffcv = -0.125
+ wpemod = 1
+ jss = 1.5e-7
+ lat = -0.00064
+ kt1 = -0.16526426
+ kt2 = -0.046114462
+ lk2 = 4.1845048e-9
+ llc = 0
+ lln = 1
+ bigsd = 0.0003327
+ lu0 = -1.1864212e-10
+ mjd = 0.335
+ mjs = 0.335
+ lua = -1.1601528e-16
+ lub = 1.1870612e-25
+ luc = 1.7407612e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = -2.3980423e-13
+ wkvth0we = 0.0
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ pk2 = -1.7678537e-15
+ aigbinv = 0.009974
+ wvoff = 6.4925381e-9
+ pu0 = 1.0845918e-15
+ prt = 0
+ pua = 1.4359661e-22
+ pub = 1.4495718e-31
+ puc = -1.3724663e-23
+ pud = 0
+ trnqsmod = 0
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 1.2300502e-9
+ ub1 = -1.4464065e-18
+ uc1 = 7.8962019e-11
+ wvsat = -0.0097711764
+ tpb = 0.0016
+ wvth0 = 5.8867412e-9
+ wa0 = 3.6413271e-7
+ ute = -0.99031694
+ wags = 1.1678647e-7
+ web = 6628.3
+ wec = -16935.0
+ wk2 = -2.0904063e-9
+ wlc = 0
+ wln = 1
+ wu0 = -2.0727529e-10
+ xgl = -8.2e-9
+ waigc = 4.3868453e-12
+ xgw = 0
+ wua = -1.2839182e-16
+ wub = -8.3225053e-26
+ wuc = -2.1668301e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ voff = -0.11093391
+ acde = 0.5
+ tpbswg = 0.001
+ lketa = -1.0921036e-8
+ vsat = 121084.96
+ wint = 0
+ xpart = 1
+ vth0 = -0.3609788
+ rgatemod = 0
+ wkt1 = -1.1364676e-8
+ wkt2 = -3.3960513e-9
+ poxedge = 1
+ wmax = 8.9974e-6
+ tnjtsswg = 1
+ aigc = 0.0068356471
+ wmin = 8.974e-7
+ egidl = 0.001
+ binunit = 2
+ ptvoff = -4.5667618e-16
+ waigsd = 1.9102262e-12
+ wua1 = -4.3482598e-16
+ wub1 = 7.4750944e-25
+ wuc1 = -1.0064978e-16
+ bigc = 0.0012521
+ wute = -8.7205605e-8
+ diomod = 1
+ wwlc = 0
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.7086399999999997e-10
+ pku0we = 0.0
+ cjswgs = 1.7086399999999997e-10
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigc = 0.15259
+ pvoff = -8.1289692e-15
+ jtsswgd = 1.75e-7
+ pvfbsdoff = 0
+ mjswgd = 0.95
+ jtsswgs = 1.75e-7
+ mjswgs = 0.95
+ cdscb = 0
+ cdscd = 0
+ tcjswg = 0.00128
+ pvsat = 0
+ wk2we = 0.0
+ pvth0 = -5.6889351e-15
+ drout = 0.56
+ paigc = -7.8179264e-18
+ a0 = 2.5342986
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 72000
+ cf = 8.17e-11
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.0010230372
+ k3 = -2.5823
+ em = 20000000.0
+ voffl = 0
+ ll = 0
+ lw = 0
+ u0 = 0.0097379054
+ w0 = 0
+ ua = 1.5508759e-10
+ ub = 1.1768184e-18
+ uc = 2.077917e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ weta0 = -1.9921431e-9
+ wetab = 6.0440267e-8
+ k2we = 5e-5
+ lpclm = 0
+ dsub = 0.5
+ dtox = 3.91e-10
+ ijthsfwd = 0.01
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ njtsswg = 6.489
+ cgidl = 1
+ fprout = 200
+ xrcrg1 = 12
+ xrcrg2 = 1
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ eta0 = 0.16744607
+ etab = -0.23671111
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.0018171133
+ pdiblcb = 0
+ pbswd = 0.9
+ wtvoff = -4.8127407e-11
+ pbsws = 0.9
+ ijthsrev = 0.01
+ pdits = 0
+ capmod = 2
+ cigsd = 0.013281
+ wku0we = 1.5e-11
+ bigbacc = 0.0054401
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ mobmod = 0
+ ppdiblc2 = -1.7911725e-15
+ kvth0we = -0.00022
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ tnoia = 0
+ peta0 = 1.6e-17
+ wketa = 2.4899578e-8
+ laigsd = -3.7090202e-15
+ tpbsw = 0.0025
+ pkvth0we = 0.0
+ cjswd = 4.8144e-11
+ cjsws = 4.8144e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ keta = -0.04361839
+ vfbsdoff = 0.01
+ )

.model pch_sf_11 pmos (
+ level = 54
+ egidl = 0.001
+ ltvfbsdoff = 0
+ toxref = 3e-9
+ ijthsfwd = 0.01
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ tnom = 25
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ ijthsrev = 0.01
+ ptvfbsdoff = 0
+ ltvoff = -2.603747e-10
+ pvfbsdoff = 0
+ wags = -5.7105665e-9
+ pvoff = 6.031093399999999e-15
+ cdscb = 0
+ cdscd = 0
+ pvsat = 0
+ wk2we = 0.0
+ voff = -0.10782222
+ njtsswg = 6.489
+ pvth0 = 3.3663808e-15
+ drout = 0.56
+ acde = 0.5
+ paigc = 1.0166993e-17
+ lku0we = 1.8e-11
+ xtsswgd = 0.32
+ vsat = 121084.96
+ xtsswgs = 0.32
+ wint = 0
+ ppdiblc2 = 8.932051e-16
+ vth0 = -0.36247368999999996
+ epsrox = 3.9
+ voffl = 0
+ wkt1 = 3.9882501e-9
+ wkt2 = -1.3862366e-8
+ ckappad = 0.6
+ wmax = 8.9974e-6
+ ckappas = 0.6
+ aigc = 0.0068328167
+ wmin = 8.974e-7
+ pdiblc1 = 0
+ pdiblc2 = 0.0082016634
+ pdiblcb = 0
+ weta0 = -1.9921431e-9
+ rdsmod = 0
+ wetab = 6.0440267e-8
+ igbmod = 1
+ lpclm = 0
+ wua1 = 1.0350058e-15
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ wub1 = -1.41997e-24
+ wuc1 = 5.1522417e-17
+ cgidl = 1
+ pbswgd = 0.8
+ bigc = 0.0012521
+ pbswgs = 0.8
+ wwlc = 0
+ bigbacc = 0.0054401
+ igcmod = 1
+ pkvth0we = 0.0
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ pbswd = 0.9
+ pbsws = 0.9
+ kvth0we = -0.00022
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigc = 0.15259
+ vfbsdoff = 0.01
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ pdits = 0
+ cigsd = 0.013281
+ paigsd = -3.7089273e-20
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ paramchk = 1
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ permod = 1
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ k2we = 5e-5
+ tnoia = 0
+ dsub = 0.5
+ dtox = 3.91e-10
+ ijthdfwd = 0.01
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ peta0 = 1.6e-17
+ voffcv = -0.125
+ wpemod = 1
+ wketa = -2.3248862e-8
+ tpbsw = 0.0025
+ eta0 = 0.16744607
+ nfactor = 1
+ etab = -0.23671111
+ cjswd = 4.8144e-11
+ cjsws = 4.8144e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ ijthdrev = 0.01
+ lpdiblc2 = 1.6477933e-9
+ nigbacc = 10
+ tpbswg = 0.001
+ scref = 1e-6
+ pigcd = 2.572
+ aigsd = 0.0063633394
+ lvoff = -9.8734428e-9
+ nigbinv = 2.171
+ ptvoff = 2.6240046e-16
+ lkvth0we = 3e-12
+ waigsd = 1.9894315e-12
+ lvsat = -8.000000000000001e-6
+ lvth0 = -2.9113088e-9
+ delta = 0.018814
+ diomod = 1
+ laigc = -4.5010295e-11
+ acnqsmod = 0
+ rnoia = 0
+ rnoib = 0
+ tvfbsdoff = 0.1
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.7086399999999997e-10
+ pku0we = 0.0
+ cjswgs = 1.7086399999999997e-10
+ fnoimod = 1
+ pketa = 2.0044574e-14
+ rbodymod = 0
+ ngate = 1.7e+20
+ eigbinv = 1.1
+ ngcon = 1
+ wpclm = -3.01194e-7
+ keta = -0.035478054
+ mjswgd = 0.95
+ mjswgs = 0.95
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ tcjswg = 0.00128
+ lags = 2.7680102e-7
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 6.6671111e-11
+ kt1l = 0
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ wpdiblc2 = -2.4522204e-9
+ lint = 6.5375218e-9
+ cigbacc = 0.245
+ lkt1 = -1.4042155e-8
+ lkt2 = -7.1896716e-9
+ lmax = 8.9908e-7
+ lmin = 4.4908e-7
+ tnoimod = 0
+ lpe0 = 6.44e-8
+ lpeb = 0
+ fprout = 200
+ minv = -0.33
+ cigbinv = 0.006
+ lua1 = 8.7159171e-17
+ lub1 = -2.6689299e-25
+ luc1 = 2.9116076e-17
+ tvoff = 0.0024887007
+ xrcrg1 = 12
+ xrcrg2 = 1
+ ndep = 1e+18
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ lwlc = 0
+ moin = 5.5538
+ wkvth0we = 0.0
+ wtvoff = -8.5607868e-10
+ nigc = 2.291
+ version = 4.5
+ a0 = 2.8862723
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ trnqsmod = 0
+ at = 72000
+ cf = 8.17e-11
+ tempmod = 0
+ ef = 1.15
+ ku0we = -0.0007
+ k1 = 0.30425
+ k2 = 0.0046668319
+ k3 = -2.5823
+ em = 20000000.0
+ ll = 0
+ lw = 0
+ beta0 = 13.32
+ u0 = 0.0097244338
+ w0 = 0
+ ua = 8.4190146e-11
+ ub = 1.1838278e-18
+ uc = 4.9200634e-11
+ ud = 0
+ leta0 = 4.8e-10
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ capmod = 2
+ ppclm = 0
+ aigbacc = 0.012071
+ wku0we = 1.5e-11
+ pags = 7.4079401e-14
+ ags = 0.8283795
+ dlcig = 2.5e-9
+ mobmod = 0
+ bgidl = 1834800000.0
+ ntox = 1.0
+ pcit = 8.000000000000001e-19
+ pclm = 1.5174437
+ cjd = 0.001270624
+ cit = -8.7888889e-5
+ cjs = 0.001270624
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 1.0572421799999999e-8
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ rgatemod = 0
+ tnjtsswg = 1
+ phin = 0.15
+ aigbinv = 0.009974
+ dmcgt = 0
+ la0 = -6.797699e-7
+ pkt1 = -4.6051461e-15
+ jsd = 1.5e-7
+ pkt2 = 4.9913693e-15
+ tcjsw = 9.34e-5
+ jss = 1.5e-7
+ lat = -0.00064
+ kt1 = -0.19603426
+ kt2 = -0.047380208
+ lk2 = -8.794787e-10
+ llc = 0
+ lln = 1
+ lu0 = -1.0665246e-10
+ mjd = 0.335
+ mjs = 0.335
+ lua = -5.2916554e-17
+ lub = 1.1246778e-25
+ luc = -7.8874906e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 4.0323955e-14
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ pk2 = 1.1838025e-15
+ pu0 = -8.8186737e-16
+ laigsd = 3.9492818e-14
+ prt = 0
+ pua = -2.1071339e-22
+ pub = -4.1382897e-32
+ puc = 1.6409308e-23
+ pud = 0
+ rbdb = 50
+ pua1 = -3.4770908e-22
+ prwb = 0
+ pub1 = 5.3383631e-31
+ prwg = 0
+ rsh = 15.2
+ puc1 = -1.6287371e-23
+ tcj = 0.000832
+ ua1 = 1.1654868e-9
+ ub1 = -1.004873e-18
+ uc1 = 4.0916434e-11
+ bigsd = 0.0003327
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ tpb = 0.0016
+ wa0 = 4.9381936e-8
+ ute = -1
+ web = 6628.3
+ wec = -16935.0
+ wk2 = -5.406874e-9
+ rdsw = 200
+ wlc = 0
+ wln = 1
+ wu0 = 2.0022293e-9
+ xgl = -8.2e-9
+ wvoff = -9.4176445e-9
+ xgw = 0
+ wua = 2.6970929e-16
+ wub = 1.2614582e-25
+ wuc = -5.5526695e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ poxedge = 1
+ wvsat = -0.0097711764
+ wvth0 = -4.2877711e-9
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ binunit = 2
+ waigc = -1.5820929e-11
+ rshg = 14.1
+ lketa = -1.8165935e-8
+ xpart = 1
+ wtvfbsdoff = 0
+ )

.model pch_sf_12 pmos (
+ level = 54
+ wkvth0we = 0.0
+ pketa = 2.9922765e-15
+ ngate = 1.7e+20
+ ngcon = 1
+ cigbacc = 0.245
+ ltvoff = -1.0992228e-10
+ wpclm = -3.01194e-7
+ trnqsmod = 0
+ gbmin = 1e-12
+ tnoimod = 0
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ cigbinv = 0.006
+ lku0we = 1.8e-11
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ epsrox = 3.9
+ rgatemod = 0
+ tnjtsswg = 1
+ rdsmod = 0
+ version = 4.5
+ igbmod = 1
+ tempmod = 0
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ pbswgd = 0.8
+ pbswgs = 0.8
+ tvoff = 0.0021467634
+ aigbacc = 0.012071
+ igcmod = 1
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ ku0we = -0.0007
+ ags = 0.29253015
+ aigbinv = 0.009974
+ beta0 = 13.32
+ keta = -0.031086208
+ leta0 = 4.8e-10
+ cjd = 0.001270624
+ cit = -0.00056559017
+ cjs = 0.001270624
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 1.38228675e-8
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ lags = 5.1257474e-7
+ ppclm = 0
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 2.7685967e-10
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ kt1l = 0
+ la0 = -1.4357692e-8
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = -0.00064
+ kt1 = -0.19916819
+ kt2 = -0.054700402
+ lk2 = 1.105099e-9
+ permod = 1
+ llc = -1.18e-13
+ lln = 0.7
+ lu0 = -4.7996045e-10
+ mjd = 0.335
+ mjs = 0.335
+ lua = -1.6078561e-16
+ lub = 5.7693033e-26
+ luc = -4.8483261e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ lint = 9.7879675e-9
+ pa0 = -2.613694e-13
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ pk2 = -5.5906497e-16
+ lkt1 = -1.2663224e-8
+ lkt2 = -3.9687861e-9
+ pu0 = -2.2461433e-17
+ lmax = 4.4908e-7
+ prt = 0
+ pua = 5.4100623e-23
+ pub = -6.3187687e-32
+ puc = -3.6550877e-24
+ pud = 0
+ dmcgt = 0
+ lmin = 2.1577e-7
+ poxedge = 1
+ tcjsw = 9.34e-5
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 1.2176874e-9
+ ub1 = -1.2376668e-18
+ lpe0 = 6.44e-8
+ uc1 = 1.0272662e-10
+ lpeb = 0
+ tpb = 0.0016
+ wa0 = 7.3504866e-7
+ ijthsfwd = 0.01
+ ute = -1
+ web = 6628.3
+ wec = -16935.0
+ wk2 = -1.4458115e-9
+ binunit = 2
+ voffcv = -0.125
+ wpemod = 1
+ wlc = 0
+ wln = 1
+ minv = -0.33
+ wu0 = 4.9034036e-11
+ xgl = -8.2e-9
+ xgw = 0
+ lua1 = 6.4190903e-17
+ lub1 = -1.6446372e-25
+ wua = -3.3214073e-16
+ wub = 1.7570216e-25
+ wuc = -9.9257962e-18
+ wud = 0
+ luc1 = 1.9195943e-18
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ ndep = 1e+18
+ bigsd = 0.0003327
+ lwlc = 0
+ moin = 5.5538
+ wvoff = 6.3544834e-9
+ nigc = 2.291
+ ijthsrev = 0.01
+ wvsat = -0.0097711764
+ wvth0 = 2.5712703900000002e-9
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ waigc = 4.9938134e-12
+ tpbswg = 0.001
+ jtsswgd = 1.75e-7
+ pags = 2.5662868e-13
+ jtsswgs = 1.75e-7
+ ntox = 1.0
+ pcit = -8.087793800000001e-17
+ lketa = -2.0098347e-8
+ pclm = 1.5174437
+ xpart = 1
+ ppdiblc2 = -1.9289508e-16
+ phin = 0.15
+ ptvoff = -6.733506e-17
+ egidl = 0.001
+ waigsd = 1.9051377e-12
+ pkt1 = 5.3381460999999995e-16
+ pkt2 = -1.2251691e-15
+ diomod = 1
+ pditsd = 0
+ pditsl = 0
+ rbdb = 50
+ cjswgd = 1.7086399999999997e-10
+ pku0we = 0.0
+ pua1 = -4.1586322e-23
+ prwb = 0
+ pub1 = 2.600258e-32
+ prwg = 0
+ cjswgs = 1.7086399999999997e-10
+ puc1 = -8.5761835e-25
+ njtsswg = 6.489
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ pkvth0we = 0.0
+ rdsw = 200
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ ckappad = 0.6
+ ckappas = 0.6
+ mjswgd = 0.95
+ mjswgs = 0.95
+ pdiblc1 = 0
+ pdiblc2 = 0.01380092
+ pvfbsdoff = 0
+ pdiblcb = 0
+ vfbsdoff = 0.01
+ pvoff = -9.086429e-16
+ tcjswg = 0.00128
+ cdscb = 0
+ cdscd = 0
+ pvsat = 0
+ wk2we = 0.0
+ pvth0 = 3.4840255000000004e-16
+ drout = 0.56
+ paramchk = 1
+ rshg = 14.1
+ paigc = 1.0085061e-18
+ bigbacc = 0.0054401
+ voffl = 0
+ weta0 = -1.9921431e-9
+ kvth0we = -0.00022
+ wetab = 6.0440267e-8
+ lpclm = 0
+ lintnoi = -5e-9
+ fprout = 200
+ ijthdfwd = 0.01
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ xrcrg1 = 12
+ xrcrg2 = 1
+ cgidl = 1
+ tnom = 25
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ wtvoff = -1.0667978e-10
+ pbswd = 0.9
+ pbsws = 0.9
+ ijthdrev = 0.01
+ lpdiblc2 = -8.1587971e-10
+ capmod = 2
+ wags = -4.2059528e-7
+ wku0we = 1.5e-11
+ wcit = 1.8563168e-10
+ pdits = 0
+ cigsd = 0.013281
+ mobmod = 0
+ voff = -0.12166106
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ acde = 0.5
+ vsat = 121084.96
+ wint = 0
+ vth0 = -0.37944280999999996
+ nfactor = 1
+ pk2we = 0.0
+ wkt1 = -7.6912059e-9
+ wkt2 = 2.6613072e-10
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ wmax = 8.9974e-6
+ aigc = 0.0067878654
+ wmin = 8.974e-7
+ lkvth0we = 3e-12
+ tnoia = 0
+ a0 = 1.3739719
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 72000
+ wua1 = 3.3927227e-16
+ cf = 8.17e-11
+ wub1 = -2.6580249e-25
+ wuc1 = 1.6454797e-17
+ ef = 1.15
+ k1 = 0.30425
+ k2 = 0.00015642806
+ k3 = -2.5823
+ em = 20000000.0
+ peta0 = 1.6e-17
+ ll = -1.18e-13
+ lw = 0
+ u0 = 0.010572861
+ w0 = 0
+ ua = 3.293471e-10
+ ub = 1.3083159e-18
+ uc = 4.2293442e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ bigc = 0.0012521
+ xw = 8.600000000000001e-9
+ wketa = 1.5506359e-8
+ wwlc = 0
+ acnqsmod = 0
+ tpbsw = 0.0025
+ nigbacc = 10
+ cjswd = 4.8144e-11
+ cjsws = 4.8144e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ cdsc = 0
+ cgbo = 0
+ rbodymod = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigc = 0.15259
+ wtvfbsdoff = 0
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ nigbinv = 2.171
+ ltvfbsdoff = 0
+ scref = 1e-6
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ pigcd = 2.572
+ wpdiblc2 = 1.6189099e-11
+ aigsd = 0.0063634291
+ fnoimod = 1
+ lvoff = -3.7843526e-9
+ eigbinv = 1.1
+ k2we = 5e-5
+ toxref = 3e-9
+ lvsat = -8.000000000000001e-6
+ dsub = 0.5
+ dtox = 3.91e-10
+ lvth0 = 4.5551043e-9
+ ptvfbsdoff = 0
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ delta = 0.018814
+ laigc = -2.5231709e-11
+ tvfbsdoff = 0.1
+ rnoia = 0
+ rnoib = 0
+ eta0 = 0.16744607
+ etab = -0.23671111
+ )

.model pch_sf_13 pmos (
+ level = 54
+ pags = 7.0037917e-14
+ lku0we = 1.8e-11
+ pvth0 = -6.0768891e-16
+ drout = 0.56
+ epsrox = 3.9
+ ntox = 1.0
+ pcit = 3.2050046000000003e-17
+ pclm = 1.5924795
+ paigc = -7.3857349e-19
+ voffl = 0
+ rdsmod = 0
+ phin = 0.15
+ igbmod = 1
+ weta0 = -1.9921431e-9
+ wetab = 6.0440267e-8
+ lkvth0we = 3e-12
+ pkt1 = 3.2071967e-16
+ pkt2 = -8.6151083e-16
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ lpclm = -1.5832542e-8
+ pbswgd = 0.8
+ pbswgs = 0.8
+ cgidl = 1
+ igcmod = 1
+ acnqsmod = 0
+ rbdb = 50
+ pua1 = -5.7774504e-23
+ prwb = 0
+ pub1 = 1.0356474e-31
+ prwg = 0
+ puc1 = 6.0450908e-24
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ rdsw = 200
+ rbodymod = 0
+ pbswd = 0.9
+ pbsws = 0.9
+ nfactor = 1
+ pdits = 0
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ permod = 1
+ rshg = 14.1
+ nigbacc = 10
+ wpdiblc2 = -2.9527442e-9
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ tnoia = 0
+ voffcv = -0.125
+ wpemod = 1
+ nigbinv = 2.171
+ peta0 = 1.6e-17
+ tnom = 25
+ wketa = 2.8638443e-8
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ tpbsw = 0.0025
+ cjswd = 4.8144e-11
+ cjsws = 4.8144e-11
+ mjswd = 0.01
+ wkvth0we = 0.0
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ trnqsmod = 0
+ fnoimod = 1
+ eigbinv = 1.1
+ wags = 4.6372111e-7
+ tpbswg = 0.001
+ wcit = -3.4957204e-10
+ voff = -0.13366619
+ acde = 0.5
+ scref = 1e-6
+ vsat = 116618.55
+ wint = 0
+ vth0 = -0.38391428
+ rgatemod = 0
+ pigcd = 2.572
+ aigsd = 0.0063634291
+ wkt1 = -6.6812774e-9
+ wkt2 = -1.4573681e-9
+ tnjtsswg = 1
+ ptvoff = -1.8786066e-17
+ wmax = 8.9974e-6
+ aigc = 0.0067673585
+ wmin = 8.974e-7
+ lvoff = -1.2512704e-9
+ waigsd = 1.9051377e-12
+ cigbacc = 0.245
+ lvsat = 0.00093441323
+ diomod = 1
+ lvth0 = 5.4985836e-9
+ wua1 = 4.1599351e-16
+ wub1 = -6.3339564e-25
+ wuc1 = -1.6259465e-17
+ tnoimod = 0
+ delta = 0.018814
+ laigc = -2.090475e-11
+ pditsd = 0
+ pditsl = 0
+ tvfbsdoff = 0.1
+ bigc = 0.0012521
+ cjswgd = 1.7086399999999997e-10
+ pku0we = 0.0
+ cjswgs = 1.7086399999999997e-10
+ wwlc = 0
+ rnoia = 0
+ rnoib = 0
+ cigbinv = 0.006
+ cdsc = 0
+ pketa = 2.2140676e-16
+ ngate = 1.7e+20
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ ngcon = 1
+ mjswgd = 0.95
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ mjswgs = 0.95
+ wpclm = -3.6917638e-7
+ cigc = 0.15259
+ tcjswg = 0.00128
+ version = 4.5
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ tempmod = 0
+ jswgs = 3.69e-13
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ aigbacc = 0.012071
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ k2we = 5e-5
+ fprout = 200
+ aigbinv = 0.009974
+ dsub = 0.5
+ dtox = 3.91e-10
+ xrcrg1 = 12
+ xrcrg2 = 1
+ ijthsfwd = 0.01
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ tvoff = 0.0019304691
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ ags = 2.6061153
+ wtvoff = -3.3676979e-10
+ eta0 = 0.16744607
+ etab = -0.23671111
+ cjd = 0.001270624
+ cit = 0.00047888384
+ cjs = 0.001270624
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 1.38228675e-8
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ ijthsrev = 0.01
+ ku0we = -0.0007
+ beta0 = 13.32
+ capmod = 2
+ leta0 = 4.8e-10
+ la0 = -4.2186937e-8
+ poxedge = 1
+ wku0we = 1.5e-11
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = -0.00035178856000000005
+ kt1 = -0.23884145
+ kt2 = -0.071460529
+ lk2 = 4.0088295e-9
+ llc = -1.18e-13
+ lln = 0.7
+ lu0 = -1.8371508999999998e-10
+ mjd = 0.335
+ ppclm = 1.4344283e-14
+ mjs = 0.335
+ lua = -2.3141614e-17
+ lub = -3.0092793e-26
+ luc = -1.1168748e-18
+ lud = 0
+ lwc = 0
+ mobmod = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = -1.7418058e-15
+ nsd = 1e+20
+ binunit = 2
+ pbd = 0.75
+ pat = -2.5956322e-9
+ pbs = 0.75
+ pk2 = -2.0925962e-16
+ dlcig = 2.5e-9
+ pu0 = 6.8306111e-19
+ bgidl = 1834800000.0
+ prt = 0
+ pua = -2.4112447e-23
+ pub = 3.4375734e-32
+ puc = -1.1236355e-25
+ pud = 0
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 2.2048659e-9
+ ub1 = -2.7884819e-18
+ ppdiblc2 = 4.3354985e-16
+ uc1 = 8.0779763e-11
+ tpb = 0.0016
+ wa0 = -4.9541389e-7
+ ute = -1
+ wat = 0.012301575
+ web = 6628.3
+ wec = -16935.0
+ wk2 = -3.1036812e-9
+ wlc = 0
+ wln = 1
+ wu0 = -6.065551e-11
+ xgl = -8.2e-9
+ xgw = 0
+ wua = 3.8537331e-17
+ wub = -2.8668372e-25
+ wuc = -2.6715958e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ wtvfbsdoff = 0
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ bigsd = 0.0003327
+ ltvfbsdoff = 0
+ pkvth0we = 0.0
+ wvoff = 5.8569161e-9
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ wvsat = -0.0057246059
+ vfbsdoff = 0.01
+ keta = -0.13181891
+ wvth0 = 7.1025095e-9
+ waigc = 1.3273811e-11
+ lags = 2.4408277e-8
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 5.6475659e-11
+ a0 = 1.505864
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ kt1l = 0
+ ptvfbsdoff = 0
+ at = 70634.069
+ paramchk = 1
+ cf = 8.17e-11
+ lketa = 1.156253e-9
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.013605325
+ k3 = -2.5823
+ em = 20000000.0
+ ll = -1.18e-13
+ lw = 0
+ u0 = 0.0091688547
+ w0 = 0
+ xpart = 1
+ ua = -3.2299413e-10
+ ub = 1.7243624e-18
+ uc = 2.4608838e-11
+ ud = 0
+ njtsswg = 6.489
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ lint = 9.7879675e-9
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ lkt1 = -4.2921669e-9
+ lkt2 = -4.3239941e-10
+ egidl = 0.001
+ lmax = 2.1577e-7
+ lmin = 9e-8
+ toxref = 3e-9
+ ckappad = 0.6
+ ckappas = 0.6
+ lpe0 = 6.44e-8
+ pdiblc1 = 0
+ pdiblc2 = 0.017260131
+ lpeb = 0
+ pdiblcb = 0
+ ijthdfwd = 0.01
+ minv = -0.33
+ lua1 = -1.4410376e-16
+ lub1 = 1.6275827e-25
+ luc1 = 6.550381e-18
+ ndep = 1e+18
+ lwlc = 0
+ moin = 5.5538
+ bigbacc = 0.0054401
+ nigc = 2.291
+ ltvoff = -6.4284173e-11
+ ijthdrev = 0.01
+ pvfbsdoff = 0
+ lpdiblc2 = -1.5457732e-9
+ kvth0we = -0.00022
+ pvoff = -8.036562e-16
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ cdscb = 0
+ cdscd = 0
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ pvsat = -8.5382639e-10
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ wk2we = 0.0
+ )

.model pch_sf_14 pmos (
+ level = 54
+ cjd = 0.001270624
+ poxedge = 1
+ cit = -0.00080588346
+ wua1 = -1.4703955e-15
+ cjs = 0.001270624
+ clc = 1e-7
+ cle = 0.6
+ wub1 = 2.631826e-24
+ bvd = 8.2
+ wuc1 = 2.762344e-16
+ bvs = 8.2
+ igcmod = 1
+ dlc = 4.0349e-9
+ k3b = 2.1176
+ tvoff = 0.0011122833
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ bigc = 0.0012521
+ wwlc = 0
+ xjbvd = 1
+ binunit = 2
+ xjbvs = 1
+ lk2we = 0.0
+ pkvth0we = 0.0
+ la0 = -2.3326483e-7
+ jsd = 1.5e-7
+ cdsc = 0
+ jss = 1.5e-7
+ lat = -0.0071902638999999996
+ kt1 = -0.2764195
+ kt2 = -0.075556865
+ lk2 = 3.5609156999999996e-9
+ llc = 0
+ cgbo = 0
+ lln = 1
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ lu0 = 2.0724492000000002e-10
+ xtid = 3
+ xtis = 3
+ mjd = 0.335
+ mjs = 0.335
+ lua = 5.4621428e-17
+ lub = 1.4388057e-26
+ luc = 1.0238844e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ cgsl = 3.0105e-11
+ njs = 1.02
+ cgso = 2.6482e-11
+ pa0 = 5.4920056e-14
+ cigc = 0.15259
+ ku0we = -0.0007
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 1.0391973e-9
+ pbs = 0.75
+ pk2 = 6.854543e-16
+ beta0 = 13.32
+ vfbsdoff = 0.01
+ pu0 = -1.2707891e-16
+ leta0 = -1.6826038999999998e-10
+ prt = 0
+ pua = -5.2218942e-24
+ pub = -3.6833051e-32
+ puc = -9.869134e-24
+ pud = 0
+ letab = 2.0996791e-8
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 8.9078668e-10
+ ub1 = -1.404024e-18
+ uc1 = 4.4088848e-11
+ ppclm = 7.4853015e-14
+ tpb = 0.0016
+ wa0 = -1.0981997e-6
+ ute = -1
+ wat = -0.026366825
+ web = 6628.3
+ wec = -16935.0
+ wk2 = -1.2621914e-8
+ wlc = 0
+ dlcig = 2.5e-9
+ permod = 1
+ wln = 1
+ wu0 = 1.2985144e-9
+ xgl = -8.2e-9
+ xgw = 0
+ bgidl = 1834800000.0
+ wua = -1.62426e-16
+ wub = 4.7085654e-25
+ wuc = 7.7079472e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ paramchk = 1
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ k2we = 5e-5
+ voffcv = -0.125
+ wpemod = 1
+ dsub = 0.5
+ dtox = 3.91e-10
+ ijthdfwd = 0.01
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ bigsd = 0.0003327
+ eta0 = 0.17434246
+ etab = -0.46008122
+ njtsswg = 6.489
+ wvoff = -4.5993296e-9
+ ijthdrev = 0.01
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ wvsat = -0.039767366
+ wvth0 = -1.4258701e-8
+ lpdiblc2 = 0
+ ckappad = 0.6
+ tpbswg = 0.001
+ ckappas = 0.6
+ waigc = -2.1370578e-11
+ pdiblc1 = 0
+ pdiblc2 = 0.00081573526
+ pdiblcb = 0
+ lketa = 9.0137227e-9
+ xpart = 1
+ ptvoff = 1.200911e-16
+ waigsd = 1.9051377e-12
+ bigbacc = 0.0054401
+ egidl = 0.001
+ lkvth0we = 3e-12
+ diomod = 1
+ kvth0we = -0.00022
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.7086399999999997e-10
+ pku0we = 0.0
+ cjswgs = 1.7086399999999997e-10
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ acnqsmod = 0
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ rbodymod = 0
+ mjswgd = 0.95
+ mjswgs = 0.95
+ pvfbsdoff = 0
+ tcjswg = 0.00128
+ keta = -0.21540901
+ pvoff = 1.7923089e-16
+ cdscb = 0
+ cdscd = 0
+ lags = -3.1969346e-8
+ pvsat = 2.3461931e-9
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ wk2we = 0.0
+ pvth0 = 1.4002649e-15
+ lcit = 1.7724378e-10
+ drout = 0.56
+ kt1l = 0
+ paigc = 2.5179991e-18
+ voffl = 0
+ wpdiblc2 = 1.6594883e-9
+ lint = 0
+ lkt1 = -7.598308999999999e-10
+ lkt2 = -4.7343777e-11
+ weta0 = 4.264371e-8
+ nfactor = 1
+ lmax = 9e-8
+ wetab = 1.3144359e-7
+ fprout = 200
+ lmin = 5.4e-8
+ lpclm = -1.0675035e-7
+ xrcrg1 = 12
+ xrcrg2 = 1
+ lpe0 = 6.44e-8
+ lpeb = 0
+ cgidl = 1
+ minv = -0.33
+ lua1 = -2.0580314e-17
+ lub1 = 3.261922e-26
+ luc1 = 9.999327e-18
+ wtvoff = -1.8141864e-9
+ ndep = 1e+18
+ lwlc = 0
+ moin = 5.5538
+ wkvth0we = 0.0
+ nigbacc = 10
+ pbswd = 0.9
+ nigc = 2.291
+ pbsws = 0.9
+ capmod = 2
+ trnqsmod = 0
+ wku0we = 1.5e-11
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ mobmod = 0
+ pdits = 0
+ nigbinv = 2.171
+ cigsd = 0.013281
+ pags = 2.8964227e-14
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ wtvfbsdoff = 0
+ ntox = 1.0
+ pcit = -6.8765404e-17
+ pclm = 2.5596902
+ rgatemod = 0
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ tnjtsswg = 1
+ ltvfbsdoff = 0
+ phin = 0.15
+ pkt1 = 1.17820041e-16
+ pkt2 = 1.7971063e-15
+ fnoimod = 1
+ tnoia = 0
+ eigbinv = 1.1
+ peta0 = -4.1797702e-15
+ petab = -6.6743123e-15
+ wketa = 8.0928346e-8
+ tpbsw = 0.0025
+ rbdb = 50
+ pua1 = 1.1954606e-22
+ prwb = 0
+ pub1 = -2.033661e-31
+ prwg = 0
+ puc1 = -2.1449333e-23
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ cjswd = 4.8144e-11
+ pvag = 2.1
+ cjsws = 4.8144e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ rdsw = 200
+ ptvfbsdoff = 0
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ cigbacc = 0.245
+ tnoimod = 0
+ rshg = 14.1
+ scref = 1e-6
+ pigcd = 2.572
+ cigbinv = 0.006
+ aigsd = 0.0063634291
+ lvoff = -2.6816163e-9
+ toxref = 3e-9
+ lvsat = -0.0059911154
+ lvth0 = -1.3102539000000001e-9
+ version = 4.5
+ ijthsfwd = 0.01
+ delta = 0.018814
+ tvfbsdoff = 0.1
+ tempmod = 0
+ laigc = -1.5433256e-11
+ tnom = 25
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ rnoia = 0
+ rnoib = 0
+ aigbacc = 0.012071
+ ltvoff = 1.2625293e-11
+ pketa = -4.6938441e-15
+ a0 = 3.5386076
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ ngate = 1.7e+20
+ at = 143383.81
+ cf = 8.17e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.0088402851
+ k3 = -2.5823
+ ijthsrev = 0.01
+ em = 20000000.0
+ ngcon = 1
+ ll = 0
+ lw = 0
+ u0 = 0.0050097056
+ wpclm = -1.0128863e-6
+ w0 = 0
+ ua = -1.1502605e-9
+ ub = 1.2511619e-18
+ uc = -9.619668e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ gbmin = 1e-12
+ wags = 9.0067526e-7
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ aigbinv = 0.009974
+ wcit = 7.2293275e-10
+ lku0we = 1.8e-11
+ wvfbsdoff = 0
+ epsrox = 3.9
+ lvfbsdoff = 0
+ voff = -0.11844975
+ acde = 0.5
+ vsat = 190294.39
+ ppdiblc2 = 0
+ rdsmod = 0
+ wint = 0
+ vth0 = -0.31147983999999995
+ igbmod = 1
+ wkt1 = -4.5227706e-9
+ wkt2 = -2.9740529e-8
+ wmax = 8.9974e-6
+ aigc = 0.0067091511
+ wmin = 8.974e-7
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ pbswgd = 0.8
+ ags = 3.2058772
+ pbswgs = 0.8
+ )

.model pch_sf_15 pmos (
+ level = 54
+ keta = 0.054978601
+ fnoimod = 1
+ pdits = 0
+ eigbinv = 1.1
+ cigsd = 0.013281
+ permod = 1
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 3.14566e-10
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ kt1l = 0
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ lint = 0
+ lkt1 = -1.3128112e-8
+ lkt2 = 1.0752811e-9
+ lmax = 5.4e-8
+ lmin = 4.5e-8
+ voffcv = -0.125
+ wpemod = 1
+ tnoia = 0
+ lpe0 = 6.44e-8
+ lpeb = 0
+ ijthsfwd = 0.01
+ cigbacc = 0.245
+ peta0 = 5.9656569000000005e-15
+ petab = -1.9628815e-15
+ minv = -0.33
+ lua1 = -1.9488641e-18
+ lub1 = 6.8003561e-26
+ wketa = -5.4843946e-8
+ luc1 = -2.115524e-18
+ tpbsw = 0.0025
+ ndep = 1e+18
+ tnoimod = 0
+ cjswd = 4.8144e-11
+ lwlc = 0
+ cjsws = 4.8144e-11
+ moin = 5.5538
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ nigc = 2.291
+ cigbinv = 0.006
+ ijthsrev = 0.01
+ tpbswg = 0.001
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ version = 4.5
+ tempmod = 0
+ ntox = 1.0
+ pcit = -6.9817065e-17
+ pclm = 1.3082183
+ scref = 1e-6
+ ptvoff = 9.8606268e-17
+ ppdiblc2 = 0
+ pigcd = 2.572
+ aigsd = 0.0063634291
+ waigsd = 1.9051377e-12
+ aigbacc = 0.012071
+ phin = 0.15
+ lvoff = -4.1725981e-9
+ diomod = 1
+ pkt1 = 1.3988109e-14
+ pkt2 = -4.0388508e-15
+ lvsat = -0.00020289408
+ lvth0 = -1.8026855e-9
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.7086399999999997e-10
+ pku0we = 0.0
+ cjswgs = 1.7086399999999997e-10
+ tvfbsdoff = 0.1
+ delta = 0.018814
+ aigbinv = 0.009974
+ laigc = -9.3796225e-12
+ rnoia = 0
+ rnoib = 0
+ rbdb = 50
+ pua1 = -1.9221227e-22
+ prwb = 0
+ pub1 = 2.2863324e-31
+ prwg = 0
+ puc1 = 2.3602641e-23
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ pkvth0we = 0.0
+ rbsb = 50
+ pvag = 2.1
+ mjswgd = 0.95
+ mjswgs = 0.95
+ rdsw = 200
+ pketa = 3.1809489e-15
+ ngate = 1.7e+20
+ ngcon = 1
+ tcjswg = 0.00128
+ wpclm = 1.8421624e-6
+ vfbsdoff = 0.01
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ poxedge = 1
+ paramchk = 1
+ rshg = 14.1
+ binunit = 2
+ ags = 2.6546816
+ cjd = 0.001270624
+ cit = -0.0031735079
+ cjs = 0.001270624
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 4.0349e-9
+ fprout = 200
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ ijthdfwd = 0.01
+ la0 = -1.5436392e-7
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0.0036843403
+ kt1 = -0.063173267
+ kt2 = -0.094912467
+ lk2 = 3.9587193e-9
+ llc = 0
+ tvoff = 0.0053332949
+ lln = 1
+ lu0 = -6.1056189e-11
+ wtvoff = -1.4437583e-9
+ tnom = 25
+ mjd = 0.335
+ mjs = 0.335
+ lua = -3.3837758e-17
+ lub = -3.4072549e-26
+ luc = -2.4014309e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = -3.174587e-14
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ xjbvd = 1
+ xjbvs = 1
+ nsd = 1e+20
+ pbd = 0.75
+ pat = -5.2399134e-10
+ lk2we = 0.0
+ pbs = 0.75
+ pk2 = 5.1035691e-16
+ pu0 = -9.701894e-17
+ prt = 0
+ pua = -1.0296702e-22
+ pub = 1.290002e-31
+ puc = 2.16225e-23
+ pud = 0
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ rsh = 15.2
+ wtvfbsdoff = 0
+ tcj = 0.000832
+ ua1 = 5.6955479e-10
+ ub1 = -2.0140988e-18
+ uc1 = 2.5296559e-10
+ ijthdrev = 0.01
+ capmod = 2
+ tpb = 0.0016
+ wa0 = 3.9604044e-7
+ ute = -1
+ wat = 0.00058470362
+ ku0we = -0.0007
+ web = 6628.3
+ wec = -16935.0
+ wk2 = -9.6029938e-9
+ wku0we = 1.5e-11
+ wlc = 0
+ beta0 = 13.32
+ wln = 1
+ wu0 = 7.8023907e-10
+ xgl = -8.2e-9
+ xgw = 0
+ lpdiblc2 = 0
+ wua = 1.5228349e-15
+ wub = -2.3883374e-24
+ leta0 = -1.8997369e-9
+ wuc = -4.6587973e-16
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ letab = 1.0403109e-8
+ ltvfbsdoff = 0
+ mobmod = 0
+ wags = 1.4000585e-6
+ ppclm = -9.0739811e-14
+ wcit = 7.4106483e-10
+ voff = -0.092743162
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ acde = 0.5
+ vsat = 90497.467
+ wint = 0
+ vth0 = -0.30298964
+ wkt1 = -2.4366569e-7
+ wkt2 = 7.087942e-8
+ wmax = 8.9974e-6
+ aigc = 0.0066047781
+ wmin = 8.974e-7
+ njtsswg = 6.489
+ dmcgt = 0
+ lkvth0we = 3e-12
+ tcjsw = 9.34e-5
+ ptvfbsdoff = 0
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ wua1 = 3.9047481e-15
+ wub1 = -4.8164385e-24
+ wuc1 = -5.0052376e-16
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.00081573526
+ pdiblcb = 0
+ bigc = 0.0012521
+ acnqsmod = 0
+ wwlc = 0
+ bigsd = 0.0003327
+ cdsc = 0
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ wvoff = 1.0199556e-9
+ rbodymod = 0
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigc = 0.15259
+ wvsat = -0.0078232946
+ bigbacc = 0.0054401
+ wvth0 = 5.0352399e-8
+ waigc = 1.173226e-10
+ kvth0we = -0.00022
+ lintnoi = -5e-9
+ lketa = -6.6687589e-9
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ xpart = 1
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ wpdiblc2 = 1.6594883e-9
+ toxref = 3e-9
+ egidl = 0.001
+ k2we = 5e-5
+ dsub = 0.5
+ dtox = 3.91e-10
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ eta0 = 0.2041955
+ etab = -0.27743155
+ ltvoff = -2.3219338e-10
+ wkvth0we = 0.0
+ pvfbsdoff = 0
+ trnqsmod = 0
+ nfactor = 1
+ pvoff = -1.4668765e-16
+ lku0we = 1.8e-11
+ cdscb = 0
+ cdscd = 0
+ epsrox = 3.9
+ pvsat = 4.9343693e-10
+ wk2we = 0.0
+ pvth0 = -2.3471789000000002e-15
+ drout = 0.56
+ paigc = -5.5262052e-18
+ rdsmod = 0
+ igbmod = 1
+ rgatemod = 0
+ voffl = 0
+ tnjtsswg = 1
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ nigbacc = 10
+ weta0 = -1.3227745e-7
+ wetab = 5.0212024e-8
+ pbswgd = 0.8
+ pbswgs = 0.8
+ lpclm = -3.4164983e-8
+ a0 = 2.1782471
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = -44109.368
+ cf = 8.17e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.015698968
+ k3 = -2.5823
+ em = 20000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.0096355868
+ w0 = 0
+ igcmod = 1
+ ua = 3.7489785e-10
+ ub = 2.0866896e-18
+ uc = 4.9437493e-10
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ cgidl = 1
+ nigbinv = 2.171
+ pbswd = 0.9
+ pbsws = 0.9
+ )

.model pch_sf_16 pmos (
+ level = 54
+ wpdiblc2 = 1.6594883e-9
+ voffcv = -0.125
+ wpemod = 1
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ bigbacc = 0.0054401
+ tnom = 25
+ kvth0we = -0.00022
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ bigsd = 0.0003327
+ lintnoi = -5e-9
+ wkvth0we = 0.0
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ wvoff = -9.7608128e-9
+ trnqsmod = 0
+ wvsat = -0.0020201595
+ tpbswg = 0.001
+ wvth0 = 9.7931233e-9
+ wags = 3.1454838e-6
+ waigc = -1.1150212e-11
+ wcit = -4.2593599e-9
+ voff = -0.099237323
+ acde = 0.5
+ lketa = 8.2510741e-9
+ ptvoff = -1.3565734e-16
+ xpart = 1
+ waigsd = 2.0479558e-12
+ vsat = 122744.64
+ wint = 0
+ rgatemod = 0
+ vth0 = -0.34523313
+ wkt1 = 3.1251908e-7
+ wkt2 = -1.0928272e-8
+ tnjtsswg = 1
+ wmax = 8.9974e-6
+ aigc = 0.0065575398
+ wmin = 8.974e-7
+ diomod = 1
+ egidl = 0.001
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.7086399999999997e-10
+ pku0we = 0.0
+ cjswgs = 1.7086399999999997e-10
+ nfactor = 1
+ wua1 = -3.8771176e-15
+ wub1 = 4.4904637e-24
+ wuc1 = 9.3089203e-17
+ bigc = 0.0012521
+ wwlc = 0
+ mjswgd = 0.95
+ mjswgs = 0.95
+ pvfbsdoff = 0
+ cdsc = 0
+ tcjswg = 0.00128
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigc = 0.15259
+ nigbacc = 10
+ pvoff = 3.8157e-16
+ cdscb = 0
+ cdscd = 0
+ pvsat = 2.0908331e-10
+ wk2we = 0.0
+ pvth0 = -3.597744e-16
+ drout = 0.56
+ paigc = 7.6896258e-19
+ nigbinv = 2.171
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ voffl = 0
+ dmdg = 0
+ fprout = 200
+ weta0 = 5.1544045e-9
+ xrcrg1 = 12
+ xrcrg2 = 1
+ wetab = 3.974597e-8
+ wtvfbsdoff = 0
+ lpclm = -2.1829165e-8
+ k2we = 5e-5
+ dsub = 0.5
+ dtox = 3.91e-10
+ ijthsfwd = 0.01
+ wtvoff = 3.3371317e-9
+ cgidl = 1
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ fnoimod = 1
+ ltvfbsdoff = 0
+ eigbinv = 1.1
+ eta0 = 0.11033512
+ etab = -0.14869011
+ capmod = 2
+ pbswd = 0.9
+ pbsws = 0.9
+ ijthsrev = 0.01
+ wku0we = 1.5e-11
+ mobmod = 0
+ pdits = 0
+ cigsd = 0.013281
+ ptvfbsdoff = 0
+ cigbacc = 0.245
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ ppdiblc2 = 0
+ tnoimod = 0
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ laigsd = 7.7486946e-16
+ cigbinv = 0.006
+ tnoia = 0
+ peta0 = -7.685038100000001e-16
+ petab = -1.4500449e-15
+ wketa = 4.9202854e-8
+ version = 4.5
+ tpbsw = 0.0025
+ tempmod = 0
+ cjswd = 4.8144e-11
+ pkvth0we = 0.0
+ cjsws = 4.8144e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ agidl = 3.2166e-9
+ aigbacc = 0.012071
+ vfbsdoff = 0.01
+ keta = -0.24950779
+ lags = 9.4399385e-8
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 1.8350138e-10
+ aigbinv = 0.009974
+ kt1l = 0
+ paramchk = 1
+ scref = 1e-6
+ pigcd = 2.572
+ aigsd = 0.0063634133
+ toxref = 3e-9
+ lint = 0
+ lvoff = -3.8543842e-9
+ lkt1 = 3.6838486e-10
+ lkt2 = 4.9336152e-10
+ lmax = 4.5e-8
+ lmin = 3.6e-8
+ lpe0 = 6.44e-8
+ lvsat = -0.0017830054
+ lpeb = 0
+ tvfbsdoff = 0.1
+ lvth0 = 2.67245694e-10
+ ijthdfwd = 0.01
+ delta = 0.018814
+ laigc = -7.0649434e-12
+ minv = -0.33
+ lua1 = -6.8231177e-17
+ lub1 = 7.1697841e-26
+ luc1 = 2.786749e-18
+ poxedge = 1
+ rnoia = 0
+ rnoib = 0
+ ndep = 1e+18
+ ltvoff = -9.8738127e-12
+ lwlc = 0
+ moin = 5.5538
+ binunit = 2
+ pketa = -1.9173443e-15
+ ngate = 1.7e+20
+ nigc = 2.291
+ ijthdrev = 0.01
+ ngcon = 1
+ wpclm = -3.2091624e-7
+ lpdiblc2 = 0
+ gbmin = 1e-12
+ lku0we = 1.8e-11
+ noff = 2.2684
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ epsrox = 3.9
+ ags = 0.72816353
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ cjd = 0.001270624
+ cit = -0.00049871975
+ cjs = 0.001270624
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ pags = -8.5525843e-14
+ dlc = 4.0349e-9
+ k3b = 2.1176
+ rdsmod = 0
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ ntox = 1.0
+ pcit = 1.7520375e-16
+ pclm = 1.0564669
+ igbmod = 1
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ la0 = -3.7737017e-8
+ jsd = 1.5e-7
+ phin = 0.15
+ jss = 1.5e-7
+ lat = -0.0025551022
+ jtsswgd = 1.75e-7
+ kt1 = -0.33861198
+ kt2 = -0.083036557
+ lk2 = 3.7383258000000006e-9
+ jtsswgs = 1.75e-7
+ llc = 0
+ lln = 1
+ pbswgd = 0.8
+ pbswgs = 0.8
+ lu0 = 1.5397989000000002e-10
+ mjd = 0.335
+ mjs = 0.335
+ lua = 2.9640356e-17
+ lub = 1.5163389e-26
+ luc = -2.5002144e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ lkvth0we = 3e-12
+ njd = 1.02
+ njs = 1.02
+ pa0 = -1.5136929e-14
+ pkt1 = -1.3264944e-14
+ pkt2 = -3.0273858e-17
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 2.5964497e-9
+ pbs = 0.75
+ pk2 = 4.883387e-16
+ igcmod = 1
+ pu0 = -4.5849539e-17
+ prt = 0
+ pua = 8.5912273e-23
+ pub = -1.727672e-31
+ puc = 8.2880171e-25
+ pud = 0
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 1.9222551e-9
+ ub1 = -2.0894923e-18
+ uc1 = 1.529192e-10
+ tvoff = 0.00079616085
+ tpb = 0.0016
+ wa0 = 5.7082474e-8
+ acnqsmod = 0
+ xjbvd = 1
+ ute = -1
+ wat = -0.063097766
+ xjbvs = 1
+ web = 6628.3
+ wec = -16935.0
+ rbdb = 50
+ wk2 = -9.1536426e-9
+ pua1 = 1.8909915e-22
+ prwb = 0
+ lk2we = 0.0
+ pub1 = -2.2740497e-31
+ prwg = 0
+ puc1 = -5.4843946e-24
+ wlc = 0
+ wln = 1
+ wu0 = -2.6403442e-10
+ xgl = -8.2e-9
+ rbpb = 50
+ rbpd = 50
+ xgw = 0
+ rbps = 50
+ rbsb = 50
+ wua = -2.3318447e-15
+ pvag = 2.1
+ wub = 3.770181e-24
+ wuc = -4.1518546e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ rdsw = 200
+ rbodymod = 0
+ paigsd = -6.9980875e-21
+ ku0we = -0.0007
+ beta0 = 13.32
+ njtsswg = 6.489
+ leta0 = 2.6994218e-9
+ letab = 4.094779e-9
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ ppclm = 1.5251044e-14
+ permod = 1
+ a0 = -0.20189383
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ ckappad = 0.6
+ at = 83226.192
+ cf = 8.17e-11
+ ckappas = 0.6
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.01120114
+ k3 = -2.5823
+ em = 20000000.0
+ dlcig = 2.5e-9
+ pdiblc1 = 0
+ pdiblc2 = 0.00081573526
+ ll = 0
+ lw = 0
+ bgidl = 1834800000.0
+ u0 = 0.0052470953999999995
+ w0 = 0
+ pdiblcb = 0
+ ua = -9.2057386e-10
+ ub = 1.0818745e-18
+ uc = 5.5311765e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ rshg = 14.1
+ )

.model pch_sf_17 pmos (
+ level = 54
+ tpbsw = 0.0025
+ aigbinv = 0.009974
+ eta0 = 0.191845
+ cjswd = 4.8144e-11
+ cjsws = 4.8144e-11
+ etab = -0.18516667
+ a0 = 2.6112
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ at = 72000
+ cf = 8.17e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.0045864754
+ k3 = -2.5823
+ em = 20000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.0096259667
+ w0 = 0
+ ua = 1.9119717e-10
+ ub = 1.0765761e-18
+ uc = -8.28048e-12
+ ud = 0
+ ijthdrev = 0.01
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ tpbswg = 0.001
+ lpdiblc2 = 0
+ ptvoff = 0
+ waigsd = 1.9350626e-12
+ scref = 1e-6
+ poxedge = 1
+ pigcd = 2.572
+ aigsd = 0.0063633642
+ diomod = 1
+ binunit = 2
+ lvoff = 0
+ pditsd = 0
+ lkvth0we = 3e-12
+ pditsl = 0
+ cjswgd = 1.7086399999999997e-10
+ pku0we = 0.0
+ cjswgs = 1.7086399999999997e-10
+ tvfbsdoff = 0.1
+ lvsat = -8.000000000000001e-6
+ lvth0 = 2.4e-10
+ delta = 0.018814
+ acnqsmod = 0
+ rnoia = 0
+ rnoib = 0
+ mjswgd = 0.95
+ mjswgs = 0.95
+ tcjswg = 0.00128
+ ngate = 1.7e+20
+ rbodymod = 0
+ ags = 0.98525249
+ ngcon = 1
+ wpclm = -5.08417e-8
+ cjd = 0.001270624
+ cit = 5e-6
+ cjs = 0.001270624
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ dlc = 1.0572421799999999e-8
+ k3b = 2.1176
+ dwb = 0
+ keta = -0.016063969
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ gbmin = 1e-12
+ wvfbsdoff = 0
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ lvfbsdoff = 0
+ wtvfbsdoff = 0
+ la0 = 0
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = -0.00064
+ lcit = -1.6e-11
+ kt1 = -0.18299632
+ lk2 = -3.2000000000000003e-10
+ kt2 = -0.042133438
+ llc = 0
+ lln = 1
+ lu0 = 8e-13
+ mjd = 0.335
+ kt1l = 0
+ mjs = 0.335
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 0
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ ltvfbsdoff = 0
+ pk2 = 0
+ wpdiblc2 = -1.7580235e-10
+ fprout = 200
+ pu0 = 0
+ prt = 0
+ pud = 0
+ lint = 6.5375218e-9
+ xrcrg1 = 12
+ xrcrg2 = 1
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 1.45515e-9
+ ub1 = -1.5029257e-18
+ uc1 = -4.3667733e-11
+ lkt1 = 4.8e-10
+ lmax = 2.001e-5
+ tpb = 0.0016
+ wa0 = 2.308488e-7
+ lmin = 8.9991e-6
+ ute = -0.96728333
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 1.3953799e-9
+ njtsswg = 6.489
+ lpe0 = 6.44e-8
+ wlc = 0
+ wln = 1
+ wu0 = 2.7482e-12
+ xgl = -8.2e-9
+ lpeb = 0
+ xgw = 0
+ wua = -1.5682603e-16
+ wub = 3.5681818e-26
+ wuc = 4.8873989e-18
+ wud = 0
+ wtvoff = -7.2458121e-11
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ tvoff = 0.0025973351
+ minv = -0.33
+ xjbvd = 1
+ xjbvs = 1
+ ckappad = 0.6
+ ckappas = 0.6
+ lk2we = 0.0
+ ndep = 1e+18
+ pdiblc1 = 0
+ pdiblc2 = 0.0032290423
+ pdiblcb = 0
+ lwlc = 0
+ ptvfbsdoff = 0
+ capmod = 2
+ wkvth0we = 0.0
+ moin = 5.5538
+ wku0we = 1.5e-11
+ nigc = 2.291
+ trnqsmod = 0
+ mobmod = 0
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = 4.8e-10
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ bigbacc = 0.0054401
+ ppclm = 0
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ kvth0we = -0.00022
+ ntox = 1.0
+ pcit = 8.000000000000001e-19
+ pclm = 1.2411167
+ rgatemod = 0
+ lintnoi = -5e-9
+ tnjtsswg = 1
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ phin = 0.15
+ vtsswgs = 1.1
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ pkt1 = 4e-17
+ bigsd = 0.0003327
+ rbdb = 50
+ prwb = 0
+ prwg = 0
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ rdsw = 200
+ wvoff = 3.276885e-9
+ wvsat = -0.017628054
+ wvth0 = 3.2194256000000006e-9
+ waigc = -7.2361068e-12
+ nfactor = 1
+ lketa = 0
+ rshg = 14.1
+ xpart = 1
+ toxref = 3e-9
+ egidl = 0.001
+ nigbacc = 10
+ ijthsfwd = 0.01
+ tnom = 25
+ ltvoff = 0
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ pvfbsdoff = 0
+ nigbinv = 2.171
+ ijthsrev = 0.01
+ lku0we = 1.8e-11
+ pvoff = -2e-17
+ epsrox = 3.9
+ wags = -3.1938756e-8
+ cdscb = 0
+ cdscd = 0
+ pvsat = 0
+ wk2we = 0.0
+ rdsmod = 0
+ pvth0 = 1.2e-16
+ fnoimod = 1
+ drout = 0.56
+ voff = -0.10917042
+ igbmod = 1
+ acde = 0.5
+ eigbinv = 1.1
+ ppdiblc2 = 0
+ vsat = 129757.01
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ wint = 0
+ voffl = 0
+ vth0 = -0.35924647
+ wkt1 = 1.4804073e-9
+ wkt2 = -8.3218931e-9
+ pbswgd = 0.8
+ pbswgs = 0.8
+ wmax = 8.974e-7
+ aigc = 0.0068422292
+ wmin = 5.374e-7
+ weta0 = -2.409757e-8
+ wetab = 1.3741e-8
+ igcmod = 1
+ lpclm = 0
+ wua1 = -5.289391e-16
+ wub1 = 6.5622425e-25
+ wuc1 = 2.3227786e-17
+ cgidl = 1
+ bigc = 0.0012521
+ wute = -1.003093e-7
+ cigbacc = 0.245
+ wwlc = 0
+ pkvth0we = 0.0
+ cdsc = 0
+ tnoimod = 0
+ pbswd = 0.9
+ pbsws = 0.9
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigc = 0.15259
+ vfbsdoff = 0.01
+ cigbinv = 0.006
+ permod = 1
+ pdits = 0
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ paramchk = 1
+ version = 4.5
+ tempmod = 0
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ voffcv = -0.125
+ wpemod = 1
+ aigbacc = 0.012071
+ k2we = 5e-5
+ tnoia = 0
+ dsub = 0.5
+ dtox = 3.91e-10
+ ijthdfwd = 0.01
+ peta0 = 1.6e-17
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ wketa = -3.7023239e-9
+ )

.model pch_sf_18 pmos (
+ level = 54
+ waigc = -9.2878513e-12
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ nigbacc = 10
+ ptvoff = 6.0745993e-16
+ pags = -1.6587566e-14
+ waigsd = 1.93751e-12
+ lketa = -8.0782883e-8
+ ntox = 1.0
+ pcit = 8.000000000000001e-19
+ pclm = 1.2411167
+ xpart = 1
+ ppdiblc2 = 2.0750737e-15
+ diomod = 1
+ nigbinv = 2.171
+ phin = 0.15
+ egidl = 0.001
+ pditsd = 0
+ pditsl = 0
+ a0 = 2.6572474
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ cjswgd = 1.7086399999999997e-10
+ pku0we = 0.0
+ cjswgs = 1.7086399999999997e-10
+ at = 72000
+ cf = 8.17e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.0050849127
+ k3 = -2.5823
+ em = 20000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.0095057581
+ pkt1 = 7.527886200000001e-15
+ pkt2 = 7.624365e-15
+ w0 = 0
+ ua = 1.8022848e-10
+ ub = 1.0497212e-18
+ uc = -5.9216956e-12
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ mjswgd = 0.95
+ mjswgs = 0.95
+ rbdb = 50
+ pua1 = 3.0135942e-22
+ prwb = 0
+ pub1 = -6.7644414e-31
+ prwg = 0
+ fnoimod = 1
+ puc1 = -4.7294542e-23
+ pvfbsdoff = 0
+ wtvfbsdoff = 0
+ tcjswg = 0.00128
+ pkvth0we = 0.0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ eigbinv = 1.1
+ pute = 3.5290383e-14
+ rdsw = 200
+ ltvfbsdoff = 0
+ vfbsdoff = 0.01
+ pvoff = 7.7887382e-16
+ cdscb = 0
+ cdscd = 0
+ pvsat = 0
+ wk2we = 0.0
+ pvth0 = -1.0464924e-15
+ drout = 0.56
+ paramchk = 1
+ paigc = 1.8445184e-17
+ rshg = 14.1
+ cigbacc = 0.245
+ fprout = 200
+ voffl = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ tnoimod = 0
+ ptvfbsdoff = 0
+ weta0 = -2.409757e-8
+ wetab = 1.3741e-8
+ lpclm = 0
+ wtvoff = -1.4002875e-10
+ cigbinv = 0.006
+ ijthdfwd = 0.01
+ cgidl = 1
+ tnom = 25
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ capmod = 2
+ version = 4.5
+ wku0we = 1.5e-11
+ tempmod = 0
+ pbswd = 0.9
+ pbsws = 0.9
+ ijthdrev = 0.01
+ mobmod = 0
+ lpdiblc2 = 3.0626629e-9
+ aigbacc = 0.012071
+ wags = -3.0093643e-8
+ pdits = 0
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ voff = -0.10728654
+ acde = 0.5
+ vsat = 129757.01
+ aigbinv = 0.009974
+ wint = 0
+ vth0 = -0.35817795999999996
+ laigsd = 5.7445099e-14
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ wkt1 = 6.4749443e-10
+ wkt2 = -9.1699871e-9
+ wmax = 8.974e-7
+ aigc = 0.0068507406
+ wmin = 5.374e-7
+ lkvth0we = 3e-12
+ tnoia = 0
+ peta0 = 1.6e-17
+ wua1 = -5.6246072e-16
+ wub1 = 7.3146831e-25
+ wuc1 = 2.8488581e-17
+ wketa = -8.2059163e-9
+ bigc = 0.0012521
+ wute = -1.0423482e-7
+ acnqsmod = 0
+ tpbsw = 0.0025
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ wwlc = 0
+ cjswd = 4.8144e-11
+ cjsws = 4.8144e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ poxedge = 1
+ cdsc = 0
+ rbodymod = 0
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigc = 0.15259
+ binunit = 2
+ toxref = 3e-9
+ scref = 1e-6
+ pigcd = 2.572
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ wpdiblc2 = -4.0662257e-10
+ aigsd = 0.0063633578
+ dmdg = 0
+ lvoff = -1.6936099e-8
+ tvfbsdoff = 0.1
+ k2we = 5e-5
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ lvsat = -8.000000000000001e-6
+ lvth0 = -9.3658678e-9
+ dsub = 0.5
+ dtox = 3.91e-10
+ delta = 0.018814
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ laigc = -7.651731e-11
+ ltvoff = -1.5996918e-9
+ ags = 0.95300429
+ rnoia = 0
+ rnoib = 0
+ cjd = 0.001270624
+ cit = 5e-6
+ cjs = 0.001270624
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 1.0572421799999999e-8
+ k3b = 2.1176
+ eta0 = 0.191845
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ etab = -0.18516667
+ dwj = 0
+ wkvth0we = 0.0
+ pketa = 4.0487295e-14
+ ngate = 1.7e+20
+ ngcon = 1
+ wpclm = -5.08417e-8
+ trnqsmod = 0
+ la0 = -4.1396638e-7
+ lku0we = 1.8e-11
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = -0.00064
+ kt1 = -0.17852273
+ kt2 = -0.039741464
+ lk2 = 4.1609517e-9
+ llc = 0
+ lln = 1
+ epsrox = 3.9
+ lu0 = 1.0814753e-9
+ mjd = 0.335
+ wvfbsdoff = 0
+ mjs = 0.335
+ lua = 9.8608496e-17
+ lub = 2.4142536e-25
+ luc = -2.1205472e-17
+ lud = 0
+ gbmin = 1e-12
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ lvfbsdoff = 0
+ njd = 1.02
+ njs = 1.02
+ pa0 = -1.9681175e-13
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ pk2 = -1.7465146e-15
+ njtsswg = 6.489
+ pu0 = -2.7146448e-18
+ rdsmod = 0
+ prt = 0
+ pua = -5.0852536e-23
+ pub = 3.3773548e-32
+ puc = 2.1258791e-23
+ pud = 0
+ igbmod = 1
+ xtsswgd = 0.32
+ rsh = 15.2
+ xtsswgs = 0.32
+ tcj = 0.000832
+ ua1 = 1.3709274e-9
+ ub1 = -1.4287011e-18
+ uc1 = -6.3574807e-11
+ tpb = 0.0016
+ wa0 = 2.527411e-7
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ ute = -0.97152091
+ ckappad = 0.6
+ ckappas = 0.6
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 1.5896529e-9
+ wlc = 0
+ rgatemod = 0
+ wln = 1
+ pdiblc1 = 0
+ pdiblc2 = 0.0028883679
+ wu0 = 3.0501627e-12
+ xgl = -8.2e-9
+ xgw = 0
+ pbswgd = 0.8
+ pdiblcb = 0
+ wua = -1.5116947e-16
+ pbswgs = 0.8
+ wub = 3.1925028e-26
+ wuc = 2.5226836e-18
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ tnjtsswg = 1
+ igcmod = 1
+ tvoff = 0.0027752763
+ bigbacc = 0.0054401
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ kvth0we = -0.00022
+ paigsd = -2.2002196e-20
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ ku0we = -0.0007
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ beta0 = 13.32
+ leta0 = 4.8e-10
+ keta = -0.0070781088
+ permod = 1
+ ppclm = 0
+ lags = 2.8991134e-7
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ dlcig = 2.5e-9
+ lcit = -1.6e-11
+ bgidl = 1834800000.0
+ kt1l = 0
+ voffcv = -0.125
+ wpemod = 1
+ lint = 6.5375218e-9
+ lkt1 = -3.9737527e-8
+ lkt2 = -2.1503841e-8
+ dmcgt = 0
+ lmax = 8.9991e-6
+ tcjsw = 9.34e-5
+ lmin = 8.9908e-7
+ lpe0 = 6.44e-8
+ lpeb = 0
+ ijthsfwd = 0.01
+ minv = -0.33
+ lua1 = 7.5716104e-16
+ lub1 = -6.6727951e-25
+ luc1 = 1.7896459e-16
+ nfactor = 1
+ bigsd = 0.0003327
+ ndep = 1e+18
+ lute = 3.8095772e-8
+ lwlc = 0
+ moin = 5.5538
+ wvoff = 3.1880225e-9
+ tpbswg = 0.001
+ ijthsrev = 0.01
+ nigc = 2.291
+ wvsat = -0.017628054
+ wvth0 = 3.3491800000000002e-9
+ noff = 2.2684
+ )

.model pch_sf_19 pmos (
+ level = 54
+ cjd = 0.001270624
+ cit = -8.7888889e-5
+ cjs = 0.001270624
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ lvsat = -8.000000000000001e-6
+ dlc = 1.0572421799999999e-8
+ k3b = 2.1176
+ lvth0 = 7.342612000000001e-11
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ ltvfbsdoff = 0
+ wua1 = -6.1430214e-16
+ wub1 = 1.1920544e-25
+ delta = 0.018814
+ wuc1 = -4.9561039e-17
+ laigc = -1.8208261e-11
+ mjswgd = 0.95
+ mjswgs = 0.95
+ njtsswg = 6.489
+ bigc = 0.0012521
+ wute = -1.2773023e-7
+ rnoia = 0
+ rnoib = 0
+ la0 = -9.6086602e-7
+ wwlc = 0
+ tcjswg = 0.00128
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = -0.00064
+ kt1 = -0.20738899
+ kt2 = -0.065812764
+ lk2 = -5.5080411e-10
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ llc = 0
+ lln = 1
+ lu0 = -1.5274407999999999e-9
+ mjd = 0.335
+ mjs = 0.335
+ lua = -3.205013e-16
+ lub = -3.7552526e-26
+ luc = 5.1848161e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 2.9499704e-13
+ pketa = -2.8529622e-14
+ ckappad = 0.6
+ cdsc = 0
+ ckappas = 0.6
+ ngate = 1.7e+20
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ pk2 = 8.8602334e-16
+ pdiblc1 = 0
+ pdiblc2 = -8.9657994e-6
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ ngcon = 1
+ xtis = 3
+ pdiblcb = 0
+ pu0 = 4.0536683e-16
+ wpclm = -5.08417e-8
+ prt = 0
+ pua = 3.1718399e-23
+ pub = 9.4535502e-32
+ puc = -3.7711192e-23
+ pud = 0
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigc = 0.15259
+ rsh = 15.2
+ wvfbsdoff = 0
+ tcj = 0.000832
+ ua1 = 2.985915e-9
+ ub1 = -2.7037422e-18
+ uc1 = 1.5248758e-10
+ lvfbsdoff = 0
+ gbmin = 1e-12
+ tpb = 0.0016
+ wa0 = -2.9985305e-7
+ jswgd = 3.69e-13
+ ptvfbsdoff = 0
+ jswgs = 3.69e-13
+ ute = -0.85901741
+ web = 6628.3
+ wec = -16935.0
+ wk2 = -1.3682549e-9
+ a0 = 3.2717414
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ wlc = 0
+ wln = 1
+ wu0 = -4.5546835e-10
+ at = 72000
+ cf = 8.17e-11
+ xgl = -8.2e-9
+ ef = 1.15
+ k1 = 0.30425
+ k2 = 0.00020919492
+ xgw = 0
+ k3 = -2.5823
+ em = 20000000.0
+ wua = -2.439458e-16
+ wub = -3.6346832e-26
+ wuc = 6.8781092e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ ll = 0
+ lw = 0
+ u0 = 0.012437123999999999
+ w0 = 0
+ ua = 6.5113837e-10
+ ub = 1.3631795e-18
+ uc = -8.8004429e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ bigbacc = 0.0054401
+ fprout = 200
+ xrcrg1 = 12
+ xrcrg2 = 1
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ kvth0we = -0.00022
+ lintnoi = -5e-9
+ wtvoff = 9.9743807e-10
+ bigbinv = 0.00149
+ k2we = 5e-5
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ dsub = 0.5
+ dtox = 3.91e-10
+ ijthsfwd = 0.01
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ tvoff = 0.00044287651
+ capmod = 2
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ wku0we = 1.5e-11
+ eta0 = 0.191845
+ etab = -0.18516667
+ mobmod = 0
+ ijthsrev = 0.01
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = 4.8e-10
+ ppclm = 0
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ nfactor = 1
+ laigsd = -3.6354984e-15
+ ppdiblc2 = -2.7249029e-15
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ nigbacc = 10
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ bigsd = 0.0003327
+ pkvth0we = 0.0
+ wvoff = 1.2743983e-8
+ nigbinv = 2.171
+ wvsat = -0.017628054
+ vfbsdoff = 0.01
+ wvth0 = 1.4292885800000004e-9
+ keta = -0.13767457
+ waigc = 2.7297355e-11
+ lags = 8.1183869e-8
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 6.6671111e-11
+ toxref = 3e-9
+ paramchk = 1
+ lketa = 3.5447968e-8
+ kt1l = 0
+ xpart = 1
+ fnoimod = 1
+ eigbinv = 1.1
+ lint = 6.5375218e-9
+ egidl = 0.001
+ lkt1 = -1.4046561e-8
+ lkt2 = 1.6996159e-9
+ lmax = 8.9908e-7
+ lmin = 4.4908e-7
+ lpe0 = 6.44e-8
+ lpeb = 0
+ ijthdfwd = 0.01
+ ltvoff = 4.7614406e-10
+ minv = -0.33
+ lua1 = -6.8017788e-16
+ lub1 = 4.6750711e-25
+ luc1 = -1.3330934e-17
+ pvfbsdoff = 0
+ ndep = 1e+18
+ lute = -6.2032341e-8
+ lwlc = 0
+ moin = 5.5538
+ cigbacc = 0.245
+ ijthdrev = 0.01
+ nigc = 2.291
+ lku0we = 1.8e-11
+ epsrox = 3.9
+ tnoimod = 0
+ lpdiblc2 = 5.64129e-9
+ pvoff = -7.7259313e-15
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ rdsmod = 0
+ cdscb = 0
+ cdscd = 0
+ cigbinv = 0.006
+ igbmod = 1
+ pvsat = 0
+ wk2we = 0.0
+ pvth0 = 6.6221102e-16
+ drout = 0.56
+ pags = 2.5130854e-13
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ paigc = -1.411565e-17
+ ntox = 1.0
+ pcit = 8.000000000000001e-19
+ pclm = 1.2411167
+ pbswgd = 0.8
+ pbswgs = 0.8
+ voffl = 0
+ version = 4.5
+ igcmod = 1
+ phin = 0.15
+ tempmod = 0
+ weta0 = -2.409757e-8
+ wetab = 1.3741e-8
+ lkvth0we = 3e-12
+ lpclm = 0
+ pkt1 = -4.6011548e-15
+ pkt2 = -3.0623252e-15
+ aigbacc = 0.012071
+ cgidl = 1
+ acnqsmod = 0
+ rbdb = 50
+ pua1 = 3.4749829e-22
+ prwb = 0
+ pub1 = -1.3153018e-31
+ prwg = 0
+ puc1 = 2.216962e-23
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ paigsd = 1.9849821e-21
+ rbsb = 50
+ pvag = 2.1
+ pute = 5.6201301e-14
+ rdsw = 200
+ rbodymod = 0
+ pbswd = 0.9
+ pbsws = 0.9
+ aigbinv = 0.009974
+ permod = 1
+ pdits = 0
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ rshg = 14.1
+ voffcv = -0.125
+ wpemod = 1
+ wpdiblc2 = 4.9866096e-9
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ poxedge = 1
+ tnoia = 0
+ binunit = 2
+ peta0 = 1.6e-17
+ wketa = 6.9341182e-8
+ tnom = 25
+ tpbsw = 0.0025
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ cjswd = 4.8144e-11
+ cjsws = 4.8144e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ wkvth0we = 0.0
+ agidl = 3.2166e-9
+ tpbswg = 0.001
+ trnqsmod = 0
+ wags = -3.311005e-7
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ ptvoff = -4.0488554e-16
+ waigsd = 1.9105581e-12
+ voff = -0.13228318
+ acde = 0.5
+ scref = 1e-6
+ diomod = 1
+ vsat = 129757.01
+ pigcd = 2.572
+ rgatemod = 0
+ wint = 0
+ aigsd = 0.0063634264
+ vth0 = -0.36878391
+ tnjtsswg = 1
+ wkt1 = 1.4275631e-8
+ wkt2 = 2.8375299e-9
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.7086399999999997e-10
+ pku0we = 0.0
+ wmax = 8.974e-7
+ wtvfbsdoff = 0
+ cjswgs = 1.7086399999999997e-10
+ aigc = 0.0067852248
+ lvoff = 5.3109112e-9
+ wmin = 5.374e-7
+ ags = 1.1875295
+ tvfbsdoff = 0.1
+ )

.model pch_sf_20 pmos (
+ level = 54
+ cjd = 0.001270624
+ cit = -0.00041212495
+ cjs = 0.001270624
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ lvsat = -8.000000000000001e-6
+ dlc = 1.38228675e-8
+ k3b = 2.1176
+ lvth0 = 6.7454743e-9
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ ltvfbsdoff = 0
+ wua1 = 2.4012676e-16
+ wub1 = -6.2487918e-26
+ delta = 0.018814
+ wuc1 = -3.9943707e-17
+ laigc = -2.2400472e-11
+ mjswgd = 0.95
+ mjswgs = 0.95
+ njtsswg = 6.489
+ bigc = 0.0012521
+ rnoia = 0
+ rnoib = 0
+ la0 = -7.2511148e-8
+ wwlc = 0
+ tcjswg = 0.00128
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = -0.00064
+ kt1 = -0.20886849
+ kt2 = -0.049681978
+ lk2 = 8.917426e-10
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ llc = -1.18e-13
+ lln = 0.7
+ lu0 = -4.801571499999999e-10
+ mjd = 0.335
+ mjs = 0.335
+ lua = -5.9775833e-17
+ lub = -8.2990392e-26
+ luc = -8.4878869e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = -2.0868237e-13
+ pketa = -1.8963071e-15
+ ckappad = 0.6
+ cdsc = 0
+ ckappas = 0.6
+ ngate = 1.7e+20
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ pk2 = -3.6576402e-16
+ pdiblc1 = 0
+ pdiblc2 = 0.01788848
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ ngcon = 1
+ xtis = 3
+ pdiblcb = 0
+ pu0 = -2.2283222e-17
+ wpclm = -5.08417e-8
+ prt = 0
+ pua = -3.7414239e-23
+ pub = 6.4271496e-32
+ puc = -3.5764571e-25
+ pud = 0
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigc = 0.15259
+ rsh = 15.2
+ wvfbsdoff = 0
+ tcj = 0.000832
+ ua1 = 1.3271195e-9
+ ub1 = -1.4620758e-18
+ uc1 = 1.6497662e-10
+ lvfbsdoff = 0
+ gbmin = 1e-12
+ tpb = 0.0016
+ wa0 = 8.4487289e-7
+ jswgd = 3.69e-13
+ ptvfbsdoff = 0
+ jswgs = 3.69e-13
+ ute = -1
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 1.4767164e-9
+ a0 = 1.2527531
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ wlc = 0
+ wln = 1
+ wu0 = 5.1646359e-10
+ at = 72000
+ cf = 8.17e-11
+ xgl = -8.2e-9
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.0030693202
+ xgw = 0
+ k3 = -2.5823
+ em = 20000000.0
+ wua = -8.6826164e-17
+ wub = 3.2435001e-26
+ wuc = -1.6113333e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ ll = -1.18e-13
+ lw = 0
+ u0 = 0.010056934
+ w0 = 0
+ ua = 5.8580479e-11
+ ub = 1.4664474e-18
+ uc = 4.9122952e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ bigbacc = 0.0054401
+ fprout = 200
+ xrcrg1 = 12
+ xrcrg2 = 1
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ kvth0we = -0.00022
+ lintnoi = -5e-9
+ wtvoff = -3.604609e-11
+ bigbinv = 0.00149
+ k2we = 5e-5
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ dsub = 0.5
+ dtox = 3.91e-10
+ ijthsfwd = 0.01
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ tvoff = 0.0020688013
+ capmod = 2
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ wku0we = 1.5e-11
+ eta0 = 0.191845
+ etab = -0.18516667
+ mobmod = 0
+ ijthsrev = 0.01
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = 4.8e-10
+ ppclm = 0
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ nfactor = 1
+ ppdiblc2 = 1.0915468e-15
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ nigbacc = 10
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ bigsd = 0.0003327
+ pkvth0we = 0.0
+ wvoff = -5.0330429e-9
+ nigbinv = 2.171
+ wvsat = -0.017628054
+ vfbsdoff = 0.01
+ wvth0 = 6.652660800000001e-9
+ keta = -0.023696099
+ waigc = -1.2459534e-12
+ lags = 6.5053339e-7
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 2.0933498e-10
+ toxref = 3e-9
+ paramchk = 1
+ lketa = -1.4702559e-8
+ kt1l = 0
+ xpart = 1
+ fnoimod = 1
+ eigbinv = 1.1
+ lint = 9.7879675e-9
+ egidl = 0.001
+ lkt1 = -1.3395579e-8
+ lkt2 = -5.3979298e-9
+ lmax = 4.4908e-7
+ lmin = 2.1577e-7
+ lpe0 = 6.44e-8
+ lpeb = 0
+ ijthdfwd = 0.01
+ ltvoff = -2.3926284e-10
+ minv = -0.33
+ lua1 = 4.9692128e-17
+ lub1 = -7.8826099e-26
+ luc1 = -1.8826114e-17
+ pvfbsdoff = 0
+ ndep = 1e+18
+ lwlc = 0
+ moin = 5.5538
+ cigbacc = 0.245
+ ijthdrev = 0.01
+ nigc = 2.291
+ lku0we = 1.8e-11
+ epsrox = 3.9
+ tnoimod = 0
+ lpdiblc2 = -2.233586e-9
+ pvoff = 9.596021e-17
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ rdsmod = 0
+ cdscb = 0
+ cdscd = 0
+ cigbinv = 0.006
+ igbmod = 1
+ pvsat = 0
+ wk2we = 0.0
+ pvth0 = -1.6360727e-15
+ drout = 0.56
+ pags = 1.3163813e-13
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ paigc = -1.5565945e-18
+ ntox = 1.0
+ pcit = -1.9700564e-17
+ pclm = 1.2411167
+ pbswgd = 0.8
+ pbswgs = 0.8
+ voffl = 0
+ version = 4.5
+ igcmod = 1
+ phin = 0.15
+ tempmod = 0
+ weta0 = -2.409757e-8
+ wetab = 1.3741e-8
+ lkvth0we = 3e-12
+ lpclm = 0
+ pkt1 = 1.1973276000000001e-15
+ pkt2 = 6.9635068e-17
+ aigbacc = 0.012071
+ cgidl = 1
+ acnqsmod = 0
+ rbdb = 50
+ pua1 = -2.8450432e-23
+ prwb = 0
+ pub1 = -5.1585101e-32
+ prwg = 0
+ puc1 = 1.7937993e-23
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ rdsw = 200
+ rbodymod = 0
+ pbswd = 0.9
+ pbsws = 0.9
+ aigbinv = 0.009974
+ permod = 1
+ pdits = 0
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ rshg = 14.1
+ voffcv = -0.125
+ wpemod = 1
+ wpdiblc2 = -3.6871397e-9
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ poxedge = 1
+ tnoia = 0
+ binunit = 2
+ peta0 = 1.6e-17
+ wketa = 8.8109206e-9
+ tnom = 25
+ tpbsw = 0.0025
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ cjswd = 4.8144e-11
+ cjsws = 4.8144e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ wkvth0we = 0.0
+ agidl = 3.2166e-9
+ tpbswg = 0.001
+ trnqsmod = 0
+ wags = -5.9122303e-8
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ ptvoff = 4.9847489e-17
+ wcit = 4.6592191e-11
+ waigsd = 1.9150694e-12
+ voff = -0.10909205
+ acde = 0.5
+ scref = 1e-6
+ diomod = 1
+ vsat = 129757.01
+ pigcd = 2.572
+ rgatemod = 0
+ wint = 0
+ aigsd = 0.0063634182
+ vth0 = -0.38394765999999997
+ tnjtsswg = 1
+ wkt1 = 1.0972613e-9
+ wkt2 = -4.2805615e-9
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.7086399999999997e-10
+ pku0we = 0.0
+ wmax = 8.974e-7
+ wtvfbsdoff = 0
+ cjswgs = 1.7086399999999997e-10
+ aigc = 0.0067947526
+ lvoff = -4.893186e-9
+ wmin = 5.374e-7
+ ags = -0.10644665
+ tvfbsdoff = 0.1
+ )

.model pch_sf_21 pmos (
+ level = 54
+ rbodymod = 0
+ version = 4.5
+ tempmod = 0
+ keta = -0.074839654
+ pvoff = 2.5972890000000003e-16
+ cdscb = 0
+ cdscd = 0
+ lags = 2.5597727e-7
+ pvsat = 0
+ aigbacc = 0.012071
+ wk2we = 0.0
+ pvth0 = 5.4710494e-16
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ drout = 0.56
+ fprout = 200
+ lcit = 1.3112816000000001e-10
+ kt1l = 0
+ paigc = 3.3660127e-18
+ xrcrg1 = 12
+ xrcrg2 = 1
+ voffl = 0
+ wpdiblc2 = 2.1803424e-9
+ lint = 9.7879675e-9
+ weta0 = -2.409757e-8
+ wtvoff = -4.3702924e-10
+ aigbinv = 0.009974
+ wetab = 1.3741e-8
+ lkt1 = -5.6843471e-9
+ lkt2 = -3.8990903e-9
+ lmax = 2.1577e-7
+ lpclm = 5.4900145e-8
+ lmin = 9e-8
+ lpe0 = 6.44e-8
+ lpeb = 0
+ cgidl = 1
+ minv = -0.33
+ capmod = 2
+ lua1 = -2.9544713e-16
+ lub1 = 3.7855773e-25
+ luc1 = 4.6029572e-17
+ wku0we = 1.5e-11
+ a0 = 0.98313605
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ ndep = 1e+18
+ at = 41320.114
+ cf = 8.17e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.016096302
+ k3 = -2.5823
+ em = 20000000.0
+ ll = -1.18e-13
+ lwlc = 0
+ lw = 0
+ u0 = 0.008606993
+ mobmod = 0
+ w0 = 0
+ wkvth0we = 0.0
+ ua = 2.7312462e-10
+ ub = 6.1180894e-19
+ uc = 6.0007215e-11
+ ud = 0
+ moin = 5.5538
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ pbswd = 0.9
+ pbsws = 0.9
+ nigc = 2.291
+ trnqsmod = 0
+ poxedge = 1
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ binunit = 2
+ pdits = 0
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ pags = -1.3976359e-13
+ ntox = 1.0
+ pcit = -3.558512e-17
+ pclm = 0.98092641
+ rgatemod = 0
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ tnjtsswg = 1
+ phin = 0.15
+ pkt1 = 1.582035e-15
+ pkt2 = 2.2793112e-15
+ tnoia = 0
+ peta0 = 1.6e-17
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ wketa = -2.2984762e-8
+ tpbsw = 0.0025
+ rbdb = 50
+ pua1 = 7.9342593e-23
+ prwb = 0
+ pub1 = -9.194958e-32
+ prwg = 0
+ puc1 = -2.9723056e-23
+ cjswd = 4.8144e-11
+ cjsws = 4.8144e-11
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ mjswd = 0.01
+ rbsb = 50
+ pvag = 2.1
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ rdsw = 200
+ toxref = 3e-9
+ njtsswg = 6.489
+ ags = 1.7634876
+ scref = 1e-6
+ rshg = 14.1
+ cjd = 0.001270624
+ cit = -4.1476524e-5
+ cjs = 0.001270624
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ xtsswgd = 0.32
+ pigcd = 2.572
+ xtsswgs = 0.32
+ dlc = 1.38228675e-8
+ aigsd = 0.0063634182
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ tvfbsdoff = 0.1
+ ckappad = 0.6
+ ckappas = 0.6
+ lvoff = -2.4249846e-9
+ pdiblc1 = 0
+ pdiblc2 = 0.011594472
+ pdiblcb = 0
+ la0 = -1.5621959e-8
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0.005833456
+ lvsat = -8.000000000000001e-6
+ kt1 = -0.24541461
+ kt2 = -0.056785482
+ lk2 = 3.6404228e-9
+ llc = -1.18e-13
+ lvth0 = 4.2239767e-9
+ lln = 0.7
+ ltvoff = -2.3342435e-10
+ lu0 = -1.7421950999999998e-10
+ mjd = 0.335
+ mjs = 0.335
+ lua = -1.0504465e-16
+ ijthsfwd = 0.01
+ lub = 9.7338322e-26
+ luc = -1.0784466e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ delta = 0.018814
+ pa0 = -2.5809676e-14
+ nsd = 1e+20
+ laigc = -2.5435198e-11
+ pbd = 0.75
+ pat = -8.1994638e-9
+ pbs = 0.75
+ pk2 = 1.2451684e-16
+ tnom = 25
+ pu0 = -7.9199366e-18
+ prt = 0
+ pua = 5.00917e-23
+ pub = -8.1076857e-32
+ puc = 8.6464743e-24
+ pud = 0
+ rnoia = 0
+ rnoib = 0
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 2.9628506e-9
+ ub1 = -3.6297717e-18
+ uc1 = -1.423963e-10
+ bigbacc = 0.0054401
+ tpb = 0.0016
+ wa0 = -2.1822352e-8
+ pketa = 4.8125819e-15
+ ute = -1
+ wat = 0.038860018
+ ngate = 1.7e+20
+ web = 6628.3
+ wec = -16935.0
+ lku0we = 1.8e-11
+ wk2 = -8.468563e-10
+ wlc = 0
+ wln = 1
+ ijthsrev = 0.01
+ wu0 = 4.4839114e-10
+ xgl = -8.2e-9
+ ngcon = 1
+ xgw = 0
+ epsrox = 3.9
+ wua = -5.0154626e-16
+ wub = 7.2128975e-25
+ wuc = -5.8786887e-17
+ wud = 0
+ wpclm = 1.8489068e-7
+ wwc = 0
+ kvth0we = -0.00022
+ wwl = 0
+ wwn = 1
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ gbmin = 1e-12
+ lintnoi = -5e-9
+ rdsmod = 0
+ jswgd = 3.69e-13
+ bigbinv = 0.00149
+ jswgs = 3.69e-13
+ wags = 1.2271418e-6
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ igbmod = 1
+ wcit = 1.2187445e-10
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ voff = -0.12078969
+ acde = 0.5
+ pbswgd = 0.8
+ pbswgs = 0.8
+ ppdiblc2 = -1.4649193e-16
+ vsat = 129757.01
+ wint = 0
+ vth0 = -0.37199742999999996
+ igcmod = 1
+ wkt1 = -7.259963e-10
+ wkt2 = -1.475296e-8
+ wmax = 8.974e-7
+ aigc = 0.0068091352
+ wmin = 5.374e-7
+ wua1 = -2.7074066e-16
+ wub1 = 1.2881293e-25
+ wuc1 = 1.8593804e-16
+ tvoff = 0.0020411307
+ bigc = 0.0012521
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ wwlc = 0
+ pkvth0we = 0.0
+ nfactor = 1
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ permod = 1
+ ku0we = -0.0007
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigc = 0.15259
+ beta0 = 13.32
+ vfbsdoff = 0.01
+ leta0 = 4.8e-10
+ ppclm = -4.9739531e-14
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ nigbacc = 10
+ paramchk = 1
+ voffcv = -0.125
+ wpemod = 1
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ nigbinv = 2.171
+ k2we = 5e-5
+ dsub = 0.5
+ ijthdfwd = 0.01
+ dtox = 3.91e-10
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ bigsd = 0.0003327
+ eta0 = 0.191845
+ tpbswg = 0.001
+ etab = -0.18516667
+ wvoff = -5.8091978e-9
+ fnoimod = 1
+ ijthdrev = 0.01
+ eigbinv = 1.1
+ wvsat = -0.017628054
+ wvth0 = -3.6941528999999994e-9
+ lpdiblc2 = -9.0555048e-10
+ wtvfbsdoff = 0
+ ptvoff = 1.3445493e-16
+ waigc = -2.4575845e-11
+ waigsd = 1.9150694e-12
+ ltvfbsdoff = 0
+ lketa = -3.9112692e-9
+ diomod = 1
+ xpart = 1
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.7086399999999997e-10
+ pku0we = 0.0
+ cjswgs = 1.7086399999999997e-10
+ cigbacc = 0.245
+ egidl = 0.001
+ lkvth0we = 3e-12
+ tnoimod = 0
+ mjswgd = 0.95
+ mjswgs = 0.95
+ cigbinv = 0.006
+ tcjswg = 0.00128
+ pvfbsdoff = 0
+ ptvfbsdoff = 0
+ acnqsmod = 0
+ )

.model pch_sf_22 pmos (
+ level = 54
+ xrcrg1 = 12
+ xrcrg2 = 1
+ paramchk = 1
+ rshg = 14.1
+ nfactor = 1
+ wtvoff = 2.0697628e-9
+ ijthdfwd = 0.01
+ capmod = 2
+ tvoff = -0.0031746364
+ tnom = 25
+ wku0we = 1.5e-11
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ mobmod = 0
+ nigbacc = 10
+ ijthdrev = 0.01
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = -9.571895e-9
+ lpdiblc2 = 0
+ letab = 1.4778454e-8
+ nigbinv = 2.171
+ wags = -2.597049e-7
+ ppclm = 2.5985382e-14
+ wcit = -2.4970451e-10
+ dlcig = 2.5e-9
+ laigsd = 2.2969081e-18
+ bgidl = 1834800000.0
+ voff = -0.11952627
+ acde = 0.5
+ vsat = 226790.48
+ wint = 0
+ vth0 = -0.33744588
+ a0 = 2.9368155
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ wkt1 = -1.289882e-8
+ wkt2 = 2.7006409e-8
+ at = 192293.99
+ cf = 8.17e-11
+ wmax = 8.974e-7
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.02088367
+ k3 = -2.5823
+ em = 20000000.0
+ fnoimod = 1
+ aigc = 0.0066428307
+ wmin = 5.374e-7
+ ll = 0
+ lw = 0
+ u0 = 0.0082035417
+ dmcgt = 0
+ w0 = 0
+ ua = -1.5734149e-9
+ ub = 3.4167628e-18
+ uc = -1.3540772e-10
+ ud = 0
+ tcjsw = 9.34e-5
+ wl = 0
+ lkvth0we = 3e-12
+ wr = 1
+ xj = 1.1e-7
+ eigbinv = 1.1
+ xl = 4e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ wua1 = 6.2697239e-16
+ wub1 = -9.8389336e-25
+ wuc1 = -5.3295995e-16
+ bigc = 0.0012521
+ acnqsmod = 0
+ bigsd = 0.0003327
+ wwlc = 0
+ wvoff = -3.6240027e-9
+ cdsc = 0
+ rbodymod = 0
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigbacc = 0.245
+ wvsat = -0.072832829
+ cigc = 0.15259
+ wvth0 = 9.2665364e-9
+ waigc = 3.8715701e-11
+ tnoimod = 0
+ toxref = 3e-9
+ lketa = 1.7736502e-8
+ cigbinv = 0.006
+ xpart = 1
+ wpdiblc2 = 6.2191766e-10
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ egidl = 0.001
+ version = 4.5
+ ltvoff = 2.5685776e-10
+ k2we = 5e-5
+ tempmod = 0
+ dsub = 0.5
+ dtox = 3.91e-10
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ pvfbsdoff = 0
+ aigbacc = 0.012071
+ eta0 = 0.29878005
+ etab = -0.34238426
+ wkvth0we = 0.0
+ lku0we = 1.8e-11
+ epsrox = 3.9
+ trnqsmod = 0
+ rdsmod = 0
+ aigbinv = 0.009974
+ pvoff = 5.4320557999999996e-17
+ igbmod = 1
+ cdscb = 0
+ cdscd = 0
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ pvsat = 5.1892488e-9
+ wk2we = 0.0
+ pvth0 = -6.711998500000001e-16
+ drout = 0.56
+ pbswgd = 0.8
+ pbswgs = 0.8
+ paigc = -2.5833927e-18
+ igcmod = 1
+ voffl = 0
+ rgatemod = 0
+ tnjtsswg = 1
+ weta0 = -7.0096749e-8
+ wetab = 2.4810139e-8
+ lpclm = -5.2812564e-8
+ poxedge = 1
+ cgidl = 1
+ binunit = 2
+ paigsd = -2.080997e-24
+ pbswd = 0.9
+ pbsws = 0.9
+ permod = 1
+ keta = -0.30513509
+ pdits = 0
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ jtsswgd = 1.75e-7
+ lcit = 1.0206861e-10
+ jtsswgs = 1.75e-7
+ voffcv = -0.125
+ wpemod = 1
+ kt1l = 0
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ lint = 0
+ lkt1 = -3.6389262e-9
+ lkt2 = 3.753071e-9
+ lmax = 9e-8
+ lmin = 5.4e-8
+ tnoia = 0
+ lpe0 = 6.44e-8
+ lpeb = 0
+ ijthsfwd = 0.01
+ peta0 = 4.3399229e-15
+ petab = -1.0404991e-15
+ wketa = 1.6222018e-7
+ minv = -0.33
+ wtvfbsdoff = 0
+ lua1 = 1.1693458e-16
+ lub1 = -2.0580342e-25
+ luc1 = -5.5456179e-17
+ tpbsw = 0.0025
+ tpbswg = 0.001
+ ndep = 1e+18
+ cjswd = 4.8144e-11
+ njtsswg = 6.489
+ cjsws = 4.8144e-11
+ mjswd = 0.01
+ lwlc = 0
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ moin = 5.5538
+ ltvfbsdoff = 0
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ ijthsrev = 0.01
+ nigc = 2.291
+ ckappad = 0.6
+ ckappas = 0.6
+ ags = 4.48665
+ pdiblc1 = 0
+ pdiblc2 = 0.0019609567
+ ptvoff = -1.0118352e-16
+ pdiblcb = 0
+ cjd = 0.001270624
+ cit = 0.00026766759
+ waigsd = 1.9150916e-12
+ cjs = 0.001270624
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ noff = 2.2684
+ bvs = 8.2
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ dlc = 4.0349e-9
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ diomod = 1
+ scref = 1e-6
+ ntox = 1.0
+ pcit = -6.566986999999999e-19
+ pclm = 2.1268063
+ la0 = -1.9926782e-7
+ pditsd = 0
+ pditsl = 0
+ ppdiblc2 = 0
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = -0.0083580887
+ cjswgd = 1.7086399999999997e-10
+ pku0we = 0.0
+ pigcd = 2.572
+ kt1 = -0.26717441
+ cjswgs = 1.7086399999999997e-10
+ kt2 = -0.13819145
+ lk2 = 4.0904354e-9
+ aigsd = 0.0063634181
+ bigbacc = 0.0054401
+ llc = 0
+ ptvfbsdoff = 0
+ lln = 1
+ lu0 = -1.3629508e-10
+ mjd = 0.335
+ mjs = 0.335
+ lua = 6.8530064e-17
+ lub = -1.6632734e-25
+ luc = 7.5845372e-18
+ lud = 0
+ tvfbsdoff = 0.1
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 2.4118768e-14
+ phin = 0.15
+ lvoff = -2.5437461e-9
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 2.0972465e-9
+ pbs = 0.75
+ pk2 = 2.0570947e-16
+ pu0 = 1.8416833e-16
+ kvth0we = -0.00022
+ prt = 0
+ pua = -1.7823119e-23
+ pub = 1.268951e-31
+ puc = -7.4643321e-24
+ pud = 0
+ pkt1 = 2.7262802999999997e-15
+ pkt2 = -1.6460695e-15
+ lvsat = -0.009129146
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = -1.4241889e-9
+ ub1 = 2.5868363e-18
+ mjswgd = 0.95
+ lvth0 = 9.761310900000001e-10
+ uc1 = 9.3723935e-10
+ mjswgs = 0.95
+ lintnoi = -5e-9
+ tpb = 0.0016
+ wa0 = -5.5297601e-7
+ delta = 0.018814
+ bigbinv = 0.00149
+ ute = -1
+ vtsswgd = 1.1
+ wat = -0.070679454
+ laigc = -9.8025804e-12
+ vtsswgs = 1.1
+ tcjswg = 0.00128
+ web = 6628.3
+ wec = -16935.0
+ wk2 = -1.7106076e-9
+ wlc = 0
+ wln = 1
+ wu0 = -1.5951011e-9
+ xgl = -8.2e-9
+ xgw = 0
+ wua = 2.2095182e-16
+ wub = -1.4911779e-24
+ wuc = 1.1260467e-16
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ rnoia = 0
+ rnoib = 0
+ rbdb = 50
+ pua1 = -5.0424332e-24
+ prwb = 0
+ pub1 = 1.2644812e-32
+ prwg = 0
+ puc1 = 3.7853356e-23
+ pkvth0we = 0.0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ pketa = -1.2596682e-14
+ ngate = 1.7e+20
+ rdsw = 200
+ ngcon = 1
+ wvfbsdoff = 0
+ wpclm = -6.2069351e-7
+ lvfbsdoff = 0
+ vfbsdoff = 0.01
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ fprout = 200
+ )

.model pch_sf_23 pmos (
+ level = 54
+ ijthsfwd = 0.01
+ dtox = 3.91e-10
+ cgidl = 1
+ wku0we = 1.5e-11
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ mobmod = 0
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ eta0 = 7.956713e-6
+ etab = -0.26192508
+ pbswd = 0.9
+ pbsws = 0.9
+ ijthsrev = 0.01
+ pdits = 0
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ ppdiblc2 = 0
+ njtsswg = 6.489
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ tnoia = 0
+ ckappad = 0.6
+ ckappas = 0.6
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ pdiblc1 = 0
+ pdiblc2 = 0.0019609567
+ pdiblcb = 0
+ peta0 = -2.7832439000000003e-15
+ petab = -1.6989745e-15
+ wketa = -4.2902456e-7
+ tpbsw = 0.0025
+ cjswd = 4.8144e-11
+ cjsws = 4.8144e-11
+ pkvth0we = 0.0
+ ags = 4.48665
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ cjd = 0.001270624
+ cit = -0.002877963
+ cjs = 0.001270624
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 4.0349e-9
+ bigbacc = 0.0054401
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ vfbsdoff = 0.01
+ a0 = 5.6551822
+ a1 = 0
+ a2 = 1
+ keta = 0.46798148
+ b0 = 0
+ b1 = 0
+ kvth0we = -0.00022
+ at = -40561.437
+ cf = 8.17e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.018874979
+ k3 = -2.5823
+ em = 20000000.0
+ la0 = -3.569331e-7
+ toxref = 3e-9
+ ll = 0
+ jsd = 1.5e-7
+ lw = 0
+ jss = 1.5e-7
+ lat = 0.0051475263
+ u0 = 0.0072084759
+ w0 = 0
+ kt1 = -0.46532049
+ kt2 = 0.0072316444
+ lk2 = 3.9739313e-9
+ ua = 5.3944309e-9
+ ub = -7.8004593e-18
+ uc = 1.0922891e-10
+ ud = 0
+ llc = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ lln = 1
+ xw = 8.600000000000001e-9
+ lu0 = -7.858127e-11
+ mjd = 0.335
+ lintnoi = -5e-9
+ mjs = 0.335
+ lua = -3.3560499e-16
+ lub = 4.8427154e-25
+ luc = -6.604387e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ bigbinv = 0.00149
+ njs = 1.02
+ pa0 = 1.517818e-13
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ nsd = 1e+20
+ lcit = 2.8451519e-10
+ pbd = 0.75
+ pat = -1.8496379e-9
+ pbs = 0.75
+ pk2 = 4.9657487e-16
+ paramchk = 1
+ pu0 = -8.1141216e-17
+ scref = 1e-6
+ kt1l = 0
+ prt = 0
+ pua = 1.7043409e-22
+ pub = -3.4061954e-31
+ puc = 5.8491101e-24
+ pud = 0
+ pigcd = 2.572
+ rsh = 15.2
+ aigsd = 0.0063634182
+ tcj = 0.000832
+ ua1 = 9.464156e-9
+ tvfbsdoff = 0.1
+ ub1 = -1.352433e-17
+ uc1 = -1.5339544e-9
+ tpb = 0.0016
+ wa0 = -2.7540628e-6
+ lint = 0
+ ute = -1
+ wat = -0.002629722
+ lvoff = -5.520199e-9
+ web = 6628.3
+ wec = -16935.0
+ wk2 = -6.7255282e-9
+ wlc = 0
+ wln = 1
+ lkt1 = 7.8535466e-9
+ lkt2 = -4.6814687e-9
+ wu0 = 2.9792015e-9
+ xgl = -8.2e-9
+ xgw = 0
+ ltvoff = -2.6406105e-10
+ wua = -3.0248621e-15
+ wub = 6.5694194e-24
+ wuc = -1.1693744e-16
+ wud = 0
+ lmax = 5.4e-8
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ lmin = 4.5e-8
+ lvsat = 0.005106104199999999
+ lpe0 = 6.44e-8
+ lvth0 = -6.5014368e-9
+ lpeb = 0
+ ijthdfwd = 0.01
+ delta = 0.018814
+ laigc = -1.6050622e-11
+ minv = -0.33
+ lua1 = -5.1458943e-16
+ lub1 = 7.2864421e-25
+ luc1 = 8.7873061e-17
+ rnoia = 0
+ rnoib = 0
+ ndep = 1e+18
+ lku0we = 1.8e-11
+ lwlc = 0
+ epsrox = 3.9
+ moin = 5.5538
+ pketa = 2.1695512e-14
+ ngate = 1.7e+20
+ wvfbsdoff = 0
+ ijthdrev = 0.01
+ lvfbsdoff = 0
+ ngcon = 1
+ nigc = 2.291
+ wpclm = -1.0386396e-6
+ nfactor = 1
+ rdsmod = 0
+ igbmod = 1
+ lpdiblc2 = 0
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ noff = 2.2684
+ pscbe1 = 926400000.0
+ noia = 2.86e+42
+ pscbe2 = 1e-20
+ noib = 2.5e+24
+ noic = 31000000000.0
+ pbswgd = 0.8
+ pbswgs = 0.8
+ igcmod = 1
+ ntox = 1.0
+ pcit = -4.2591024e-17
+ pclm = 4.4879115
+ nigbacc = 10
+ phin = 0.15
+ lkvth0we = 3e-12
+ pkt1 = -5.0212736e-15
+ pkt2 = 1.1767646e-15
+ nigbinv = 2.171
+ tvoff = 0.0058067224
+ acnqsmod = 0
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ rbdb = 50
+ pua1 = 2.7224008e-22
+ prwb = 0
+ pub1 = -3.6990718e-31
+ prwg = 0
+ puc1 = -5.7927018e-23
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ permod = 1
+ rbodymod = 0
+ rdsw = 200
+ ku0we = -0.0007
+ beta0 = 13.32
+ fnoimod = 1
+ leta0 = 7.7568866e-9
+ letab = 1.0111821e-8
+ eigbinv = 1.1
+ ppclm = 5.0226256e-14
+ voffcv = -0.125
+ wpemod = 1
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ rshg = 14.1
+ wtvfbsdoff = 0
+ wpdiblc2 = 6.2191766e-10
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ ltvfbsdoff = 0
+ cigbacc = 0.245
+ tnoimod = 0
+ tnom = 25
+ tpbswg = 0.001
+ bigsd = 0.0003327
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ cigbinv = 0.006
+ wkvth0we = 0.0
+ wvoff = -2.1208799e-8
+ trnqsmod = 0
+ wvsat = 0.09105966
+ ptvoff = 1.2747838e-16
+ ptvfbsdoff = 0
+ wvth0 = -3.5235008e-8
+ waigsd = 1.9150557e-12
+ version = 4.5
+ waigc = -1.4751759e-11
+ wags = -2.597049e-7
+ tempmod = 0
+ wcit = 4.7330111e-10
+ diomod = 1
+ voff = -0.068208113
+ lketa = -2.7104259e-8
+ acde = 0.5
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.7086399999999997e-10
+ pku0we = 0.0
+ cjswgs = 1.7086399999999997e-10
+ aigbacc = 0.012071
+ xpart = 1
+ rgatemod = 0
+ vsat = -18644.867
+ wint = 0
+ vth0 = -0.2085223
+ tnjtsswg = 1
+ wkt1 = 1.206797e-7
+ wkt2 = -2.1663145e-8
+ egidl = 0.001
+ wmax = 8.974e-7
+ aigc = 0.0067505556
+ wmin = 5.374e-7
+ mjswgd = 0.95
+ mjswgs = 0.95
+ aigbinv = 0.009974
+ tcjswg = 0.00128
+ pvfbsdoff = 0
+ wua1 = -4.1537606e-15
+ wub1 = 5.6118307e-24
+ wuc1 = 1.1184258e-15
+ bigc = 0.0012521
+ wwlc = 0
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigc = 0.15259
+ pvoff = 1.0742388e-15
+ poxedge = 1
+ cdscb = 0
+ cdscd = 0
+ fprout = 200
+ pvsat = -4.3165155e-9
+ wk2we = 0.0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ pvth0 = 1.9098897e-15
+ drout = 0.56
+ binunit = 2
+ paigc = 5.1772001e-19
+ voffl = 0
+ dmcg = 3.1e-8
+ wtvoff = -1.8726837e-9
+ dmci = 3.1e-8
+ dmdg = 0
+ weta0 = 5.2716471e-8
+ wetab = 3.6163164e-8
+ lpclm = -1.8975667e-7
+ k2we = 5e-5
+ capmod = 2
+ dsub = 0.5
+ )

.model pch_sf_24 pmos (
+ level = 54
+ beta0 = 13.32
+ leta0 = 9.3580824e-10
+ letab = 2.8639817e-9
+ cigbacc = 0.245
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ ppclm = -6.983762e-15
+ laigsd = -1.7489044e-14
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ tnoimod = 0
+ ntox = 1.0
+ pcit = -2.3859875e-16
+ pclm = 0.55996802
+ rgatemod = 0
+ cigbinv = 0.006
+ tnjtsswg = 1
+ phin = 0.15
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ pkt1 = 8.083990900000001e-15
+ pkt2 = -6.3201272e-16
+ version = 4.5
+ tempmod = 0
+ bigsd = 0.0003327
+ rbdb = 50
+ pua1 = -2.7866327e-22
+ prwb = 0
+ pub1 = 3.2786288e-31
+ prwg = 0
+ puc1 = 2.5974765e-23
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ aigbacc = 0.012071
+ wvoff = -2.6959456e-8
+ rdsw = 200
+ wvsat = 0.037826603
+ wvth0 = -2.9575681e-9
+ toxref = 3e-9
+ waigc = -9.7737582e-11
+ aigbinv = 0.009974
+ lketa = 1.4220453e-8
+ rshg = 14.1
+ xpart = 1
+ egidl = 0.001
+ ltvoff = -2.5344658e-10
+ pvfbsdoff = 0
+ ijthsfwd = 0.01
+ poxedge = 1
+ a0 = -2.5402778
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ tnom = 25
+ at = 213109.93
+ cf = 8.17e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.022656115
+ k3 = -2.5823
+ em = 20000000.0
+ lku0we = 1.8e-11
+ ll = 0
+ lw = 0
+ u0 = 0.0013178574
+ w0 = 0
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ ua = -6.0379704e-9
+ ub = 8.1069989e-18
+ uc = -2.2784413e-10
+ ud = 0
+ binunit = 2
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ epsrox = 3.9
+ xw = 8.600000000000001e-9
+ ijthsrev = 0.01
+ rdsmod = 0
+ igbmod = 1
+ pvoff = 1.3560210000000001e-15
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ wags = -2.597049e-7
+ cdscb = 0
+ cdscd = 0
+ pbswgd = 0.8
+ pbswgs = 0.8
+ pvsat = -1.7080957e-9
+ wcit = 4.4734589e-9
+ wk2we = 0.0
+ pvth0 = 3.2829517e-16
+ drout = 0.56
+ igcmod = 1
+ voff = -0.080254273
+ paigc = 4.5840253e-18
+ acde = 0.5
+ ppdiblc2 = 0
+ voffl = 0
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ vsat = 78763.66
+ wint = 0
+ vth0 = -0.33115952
+ wkt1 = -1.4677468e-7
+ wkt2 = 1.5250678e-8
+ wmax = 8.974e-7
+ weta0 = -2.1009528e-8
+ aigc = 0.0066531108
+ wetab = 8.325777e-9
+ wmin = 5.374e-7
+ lpclm = 2.7125638e-9
+ cgidl = 1
+ paigsd = 9.5490179e-21
+ wua1 = 7.089165e-15
+ wub1 = -8.6283747e-24
+ wuc1 = -5.9385548e-16
+ bigc = 0.0012521
+ wwlc = 0
+ pkvth0we = 0.0
+ permod = 1
+ cdsc = 0
+ pbswd = 0.9
+ pbsws = 0.9
+ njtsswg = 6.489
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ wtvfbsdoff = 0
+ cigc = 0.15259
+ vfbsdoff = 0.01
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ ckappad = 0.6
+ ckappas = 0.6
+ pdits = 0
+ voffcv = -0.125
+ wpemod = 1
+ pdiblc1 = 0
+ pdiblc2 = 0.0019609567
+ cigsd = 0.013281
+ ltvfbsdoff = 0
+ pdiblcb = 0
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ paramchk = 1
+ pk2we = 0.0
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ bigbacc = 0.0054401
+ tnoia = 0
+ k2we = 5e-5
+ ags = 4.48665
+ ijthdfwd = 0.01
+ dsub = 0.5
+ dtox = 3.91e-10
+ kvth0we = -0.00022
+ peta0 = 8.2933004e-16
+ ptvfbsdoff = 0
+ petab = -3.349425e-16
+ cjd = 0.001270624
+ cit = -0.010137593
+ cjs = 0.001270624
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dvt0 = 3.48
+ tpbswg = 0.001
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ wketa = 1.6324308e-7
+ dlc = 4.0349e-9
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ tpbsw = 0.0025
+ dwg = 0
+ lintnoi = -5e-9
+ dwj = 0
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ cjswd = 4.8144e-11
+ cjsws = 4.8144e-11
+ mjswd = 0.01
+ eta0 = 0.13921364
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ etab = -0.11400999
+ la0 = 4.4644444e-8
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = -0.0072823707
+ kt1 = 0.16833478
+ kt2 = -0.11193164
+ lk2 = 4.159207e-9
+ ijthdrev = 0.01
+ llc = 0
+ lln = 1
+ lu0 = 2.1005904e-10
+ mjd = 0.335
+ ptvoff = 8.5019581e-17
+ mjs = 0.335
+ lua = 2.2458267e-16
+ lub = -2.9519392e-25
+ luc = 9.9121919e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = -8.9774533e-14
+ waigsd = 1.7201778e-12
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 6.8793549e-9
+ pbs = 0.75
+ lpdiblc2 = 0
+ pk2 = 1.0702031e-16
+ pu0 = -9.6657248e-17
+ prt = 0
+ pua = -9.0705467e-23
+ pub = 1.0841652e-31
+ puc = -1.0416838e-23
+ pud = 0
+ diomod = 1
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = -1.018181e-8
+ ub1 = 1.2390462e-17
+ uc1 = 9.111363e-10
+ tpb = 0.0016
+ wa0 = 2.1756583e-6
+ ute = -1
+ wat = -0.18077244
+ pditsd = 0
+ web = 6628.3
+ wec = -16935.0
+ pditsl = 0
+ wk2 = 1.2245648e-9
+ cjswgd = 1.7086399999999997e-10
+ pku0we = 0.0
+ cjswgs = 1.7086399999999997e-10
+ wlc = 0
+ wln = 1
+ wu0 = 3.2958552e-9
+ xgl = -8.2e-9
+ xgw = 0
+ scref = 1e-6
+ wua = 2.3045166e-15
+ wub = -2.5945817e-24
+ wuc = 2.150207e-16
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ tvfbsdoff = 0.1
+ pigcd = 2.572
+ aigsd = 0.0063637751
+ lvoff = -4.9299372e-9
+ mjswgd = 0.95
+ mjswgs = 0.95
+ lkvth0we = 3e-12
+ nfactor = 1
+ lvsat = 0.00033308628000000004
+ tcjswg = 0.00128
+ lvth0 = -4.9221299e-10
+ delta = 0.018814
+ laigc = -1.1275829e-11
+ acnqsmod = 0
+ rnoia = 0
+ rnoib = 0
+ wvfbsdoff = 0
+ pketa = -7.3256019e-15
+ ngate = 1.7e+20
+ lvfbsdoff = 0
+ rbodymod = 0
+ nigbacc = 10
+ ngcon = 1
+ wpclm = 1.2891178e-7
+ gbmin = 1e-12
+ keta = -0.37538
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ fprout = 200
+ xrcrg1 = 12
+ xrcrg2 = 1
+ nigbinv = 2.171
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 6.4023704e-10
+ kt1l = 0
+ wtvoff = -1.0061777e-9
+ wpdiblc2 = 6.2191766e-10
+ lint = 0
+ lkt1 = -2.3195561e-8
+ lkt2 = 1.1575324e-9
+ lmax = 4.5e-8
+ lmin = 3.6e-8
+ capmod = 2
+ fnoimod = 1
+ lpe0 = 6.44e-8
+ lpeb = 0
+ wku0we = 1.5e-11
+ eigbinv = 1.1
+ tvoff = 0.0055901005
+ mobmod = 0
+ minv = -0.33
+ lua1 = 4.4806289e-16
+ lub1 = -5.4118058e-25
+ luc1 = -3.1936385e-17
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ ndep = 1e+18
+ wkvth0we = 0.0
+ lwlc = 0
+ moin = 5.5538
+ nigc = 2.291
+ trnqsmod = 0
+ ku0we = -0.0007
+ )

.model pch_sf_25 pmos (
+ level = 54
+ wint = 0
+ ags = 0.93810347
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ vth0 = -0.35398248
+ wkt1 = -1.5318394e-9
+ wkt2 = 2.21858e-9
+ cjd = 0.001270624
+ cit = 5e-6
+ cjs = 0.001270624
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ wmax = 5.374e-7
+ bvs = 8.2
+ aigc = 0.0068215676
+ wmin = 2.674e-7
+ dlc = 1.0572421799999999e-8
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ k3b = 2.1176
+ lkvth0we = 3e-12
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ tnoia = 0
+ peta0 = 1.6e-17
+ la0 = 0
+ wua1 = 1.6452204e-16
+ wub1 = -6.9710259e-26
+ wuc1 = 2.1709154e-17
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = -0.00064
+ wketa = 2.2687563e-8
+ kt1 = -0.17747938
+ lk2 = -3.2000000000000003e-10
+ kt2 = -0.061438333
+ llc = 0
+ lln = 1
+ lu0 = 8e-13
+ tpbsw = 0.0025
+ acnqsmod = 0
+ mjd = 0.335
+ bigc = 0.0012521
+ mjs = 0.335
+ wute = 3.2371733e-8
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ wwlc = 0
+ pa0 = 0
+ cjswd = 4.8144e-11
+ nsd = 1e+20
+ cjsws = 4.8144e-11
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ pk2 = 0
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ pu0 = 0
+ prt = 0
+ pud = 0
+ rbodymod = 0
+ cdsc = 0
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 1.8507467e-10
+ ub1 = -1.7337534e-19
+ uc1 = -4.0886356e-11
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ tpb = 0.0016
+ wa0 = -1.5013787e-7
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigc = 0.15259
+ ute = -1.2102889
+ toxref = 3e-9
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 4.440518e-10
+ wlc = 0
+ wln = 1
+ wu0 = 3.7953067e-11
+ xgl = -8.2e-9
+ xgw = 0
+ nfactor = 1
+ wua = -1.5196107e-16
+ wub = 9.0507286e-26
+ wuc = 5.3799588e-18
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ scref = 1e-6
+ tvfbsdoff = 0.1
+ pigcd = 2.572
+ aigsd = 0.0063632886
+ wpdiblc2 = -7.7579138e-11
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ ltvoff = 0
+ lvoff = 0
+ nigbacc = 10
+ lvsat = -8.000000000000001e-6
+ k2we = 5e-5
+ lvth0 = 2.4e-10
+ dsub = 0.5
+ dtox = 3.91e-10
+ delta = 0.018814
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ lku0we = 1.8e-11
+ rnoia = 0
+ rnoib = 0
+ epsrox = 3.9
+ nigbinv = 2.171
+ eta0 = 0.17962267
+ wvfbsdoff = 0
+ wkvth0we = 0.0
+ etab = -0.19577778
+ lvfbsdoff = 0
+ ngate = 1.7e+20
+ rdsmod = 0
+ ngcon = 1
+ igbmod = 1
+ wpclm = -1.1447315e-8
+ trnqsmod = 0
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ pbswgd = 0.8
+ pbswgs = 0.8
+ fnoimod = 1
+ eigbinv = 1.1
+ igcmod = 1
+ a0 = 3.3089778
+ a1 = 0
+ a2 = 1
+ rgatemod = 0
+ b0 = 0
+ b1 = 0
+ at = 72000
+ cf = 8.17e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.0028441163
+ k3 = -2.5823
+ em = 20000000.0
+ tnjtsswg = 1
+ ll = 0
+ lw = 0
+ u0 = 0.0095614889
+ w0 = 0
+ ua = 1.8228697e-10
+ ub = 9.7616315e-19
+ uc = -9.1826044e-12
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ wtvfbsdoff = 0
+ cigbacc = 0.245
+ tvoff = 0.0026578776
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ permod = 1
+ ltvfbsdoff = 0
+ tnoimod = 0
+ cigbinv = 0.006
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = 4.8e-10
+ keta = -0.064397096
+ voffcv = -0.125
+ wpemod = 1
+ ppclm = 0
+ version = 4.5
+ dlcig = 2.5e-9
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ bgidl = 1834800000.0
+ lcit = -1.6e-11
+ tempmod = 0
+ ptvfbsdoff = 0
+ kt1l = 0
+ aigbacc = 0.012071
+ lint = 6.5375218e-9
+ dmcgt = 0
+ lkt1 = 4.8e-10
+ tcjsw = 9.34e-5
+ lmax = 2.001e-5
+ lmin = 8.9991e-6
+ lpe0 = 6.44e-8
+ lpeb = 0
+ ijthsfwd = 0.01
+ tpbswg = 0.001
+ minv = -0.33
+ aigbinv = 0.009974
+ bigsd = 0.0003327
+ ndep = 1e+18
+ lwlc = 0
+ moin = 5.5538
+ wvoff = 2.5521431e-9
+ ptvoff = 0
+ ijthsrev = 0.01
+ nigc = 2.291
+ waigsd = 1.9763167e-12
+ wvsat = 0.0034765009
+ wvth0 = 3.452853000000003e-10
+ diomod = 1
+ waigc = 4.045116e-12
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.7086399999999997e-10
+ pku0we = 0.0
+ cjswgs = 1.7086399999999997e-10
+ poxedge = 1
+ lketa = 0
+ ntox = 1.0
+ xpart = 1
+ pcit = 8.000000000000001e-19
+ pclm = 1.1689658
+ ppdiblc2 = 0
+ binunit = 2
+ egidl = 0.001
+ mjswgd = 0.95
+ mjswgs = 0.95
+ phin = 0.15
+ tcjswg = 0.00128
+ pkt1 = 4e-17
+ pvfbsdoff = 0
+ rbdb = 50
+ prwb = 0
+ prwg = 0
+ pkvth0we = 0.0
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ jtsswgd = 1.75e-7
+ rdsw = 200
+ jtsswgs = 1.75e-7
+ vfbsdoff = 0.01
+ fprout = 200
+ pvoff = -2e-17
+ xrcrg1 = 12
+ xrcrg2 = 1
+ cdscb = 0
+ cdscd = 0
+ pvsat = 0
+ wk2we = 0.0
+ pvth0 = 1.2e-16
+ drout = 0.56
+ paramchk = 1
+ wtvoff = -1.0551434e-10
+ rshg = 14.1
+ voffl = 0
+ weta0 = -1.7424176e-8
+ wetab = 1.9534667e-8
+ njtsswg = 6.489
+ capmod = 2
+ lpclm = 0
+ wku0we = 1.5e-11
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ ijthdfwd = 0.01
+ cgidl = 1
+ mobmod = 0
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.0030491463
+ tnom = 25
+ pdiblcb = 0
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ pbswd = 0.9
+ pbsws = 0.9
+ ijthdrev = 0.01
+ lpdiblc2 = 0
+ bigbacc = 0.0054401
+ wags = -6.1953916e-9
+ pdits = 0
+ cigsd = 0.013281
+ kvth0we = -0.00022
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ voff = -0.10784306
+ acde = 0.5
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ vsat = 91103.982
+ pk2we = 0.0
+ )

.model pch_sf_26 pmos (
+ level = 54
+ bigsd = 0.0003327
+ poxedge = 1
+ pkvth0we = 0.0
+ wvoff = 2.9007224e-9
+ binunit = 2
+ toxref = 3e-9
+ wvsat = 0.0034765009
+ wvth0 = 2.837108000000003e-10
+ vfbsdoff = 0.01
+ keta = -0.06875265
+ waigc = 4.3476029e-12
+ lags = 1.0877241e-7
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = -1.6e-11
+ lketa = 3.9156432e-8
+ paramchk = 1
+ kt1l = 0
+ xpart = 1
+ ltvoff = -4.4286369e-10
+ egidl = 0.001
+ lint = 6.5375218e-9
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ lkt1 = -3.4373729e-8
+ lkt2 = -1.4641311e-8
+ lmax = 8.9991e-6
+ pvfbsdoff = 0
+ lmin = 8.9908e-7
+ lpe0 = 6.44e-8
+ ijthdfwd = 0.01
+ lpeb = 0
+ lku0we = 1.8e-11
+ minv = -0.33
+ epsrox = 3.9
+ lua1 = 1.4818924e-15
+ lub1 = -2.0711788e-24
+ luc1 = 2.2491171e-16
+ ndep = 1e+18
+ lute = 1.330224e-7
+ rdsmod = 0
+ lwlc = 0
+ moin = 5.5538
+ igbmod = 1
+ ijthdrev = 0.01
+ nigc = 2.291
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ lpdiblc2 = 8.2033961e-9
+ njtsswg = 6.489
+ pbswgd = 0.8
+ pvoff = -3.1537282e-15
+ pbswgs = 0.8
+ noff = 2.2684
+ cdscb = 0
+ cdscd = 0
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ igcmod = 1
+ pvsat = 0
+ wk2we = 0.0
+ pvth0 = 6.7355474e-16
+ drout = 0.56
+ ckappad = 0.6
+ ckappas = 0.6
+ pags = 8.2314292e-14
+ wtvfbsdoff = 0
+ pdiblc1 = 0
+ pdiblc2 = 0.002136644
+ paigc = -2.7193569e-18
+ pdiblcb = 0
+ ntox = 1.0
+ pcit = 8.000000000000001e-19
+ pclm = 1.1689658
+ voffl = 0
+ ltvfbsdoff = 0
+ weta0 = -1.7424176e-8
+ phin = 0.15
+ wetab = 1.9534667e-8
+ lkvth0we = 3e-12
+ lpclm = 0
+ paigsd = -4.5957918e-20
+ pkt1 = 4.5992525999999995e-15
+ pkt2 = 3.8774237e-15
+ bigbacc = 0.0054401
+ cgidl = 1
+ permod = 1
+ acnqsmod = 0
+ kvth0we = -0.00022
+ rbdb = 50
+ pua1 = -9.4343892e-23
+ prwb = 0
+ pub1 = 9.0084871e-32
+ prwg = 0
+ puc1 = -7.238167e-23
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ lintnoi = -5e-9
+ pute = -1.6539558e-14
+ bigbinv = 0.00149
+ rbodymod = 0
+ pbswd = 0.9
+ pbsws = 0.9
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ rdsw = 200
+ ptvfbsdoff = 0
+ a0 = 3.4253346
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 72000
+ cf = 8.17e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.0024652651
+ k3 = -2.5823
+ em = 20000000.0
+ ll = 0
+ voffcv = -0.125
+ lw = 0
+ wpemod = 1
+ u0 = 0.009445427499999999
+ w0 = 0
+ ua = 1.8429003e-10
+ ub = 9.3982253e-19
+ uc = -1.1498405e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ pdits = 0
+ cigsd = 0.013281
+ ags = 0.9260042
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ cjd = 0.001270624
+ cit = 5e-6
+ cjs = 0.001270624
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 1.0572421799999999e-8
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ rshg = 14.1
+ wpdiblc2 = 3.818702e-12
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ la0 = -1.0460478e-6
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = -0.00064
+ kt1 = -0.17360244
+ kt2 = -0.059809712
+ lk2 = -3.7258721e-9
+ llc = 0
+ lln = 1
+ lu0 = 1.0441917e-9
+ mjd = 0.335
+ mjs = 0.335
+ lua = -1.8007487e-17
+ lub = 3.2670219e-25
+ luc = 2.0819042e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ tnoia = 0
+ njd = 1.02
+ njs = 1.02
+ pa0 = 1.483047e-13
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ tpbswg = 0.001
+ pk2 = 2.5596912e-15
+ pu0 = 1.7642195e-17
+ nfactor = 1
+ peta0 = 1.6e-17
+ prt = 0
+ pua = 1.2819791e-23
+ pub = -1.2787603e-32
+ puc = -1.6865938e-24
+ pud = 0
+ wketa = 2.5468383e-8
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 2.0236805e-11
+ ub1 = 5.7011626e-20
+ uc1 = -6.5904343e-11
+ tnom = 25
+ tpbsw = 0.0025
+ tpb = 0.0016
+ wa0 = -1.666345e-7
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ ute = -1.2250856
+ cjswd = 4.8144e-11
+ cjsws = 4.8144e-11
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 1.5932531e-10
+ mjswd = 0.01
+ wlc = 0
+ mjsws = 0.01
+ wln = 1
+ agidl = 3.2166e-9
+ wu0 = 3.5990642e-11
+ wkvth0we = 0.0
+ xgl = -8.2e-9
+ xgw = 0
+ wua = -1.5338707e-16
+ wub = 9.1929712e-26
+ wuc = 5.5675666e-18
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ ptvoff = -2.4168192e-17
+ waigsd = 1.9814288e-12
+ trnqsmod = 0
+ nigbacc = 10
+ diomod = 1
+ wags = -1.5351598e-8
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.7086399999999997e-10
+ pku0we = 0.0
+ cjswgs = 1.7086399999999997e-10
+ tvfbsdoff = 0.1
+ voff = -0.10676035
+ scref = 1e-6
+ acde = 0.5
+ nigbinv = 2.171
+ pigcd = 2.572
+ rgatemod = 0
+ aigsd = 0.0063632773
+ vsat = 91103.982
+ wint = 0
+ vth0 = -0.35256355
+ tnjtsswg = 1
+ mjswgd = 0.95
+ mjswgs = 0.95
+ wkt1 = -2.0389865e-9
+ wkt2 = 1.7872759e-9
+ lvoff = -9.7335308e-9
+ wmax = 5.374e-7
+ aigc = 0.0068257672
+ wmin = 2.674e-7
+ tcjswg = 0.00128
+ lvsat = -8.000000000000001e-6
+ lvth0 = -1.2516136999999998e-8
+ delta = 0.018814
+ laigc = -3.7754415e-11
+ wua1 = 1.7501635e-16
+ wub1 = -7.9730823e-26
+ wuc1 = 2.9760508e-17
+ fnoimod = 1
+ rnoia = 0
+ rnoib = 0
+ bigc = 0.0012521
+ eigbinv = 1.1
+ wute = 3.4211506e-8
+ wwlc = 0
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ pketa = -2.4999571e-14
+ ngate = 1.7e+20
+ cdsc = 0
+ ngcon = 1
+ cgbo = 0
+ wpclm = -1.1447315e-8
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ fprout = 200
+ cigc = 0.15259
+ gbmin = 1e-12
+ xrcrg1 = 12
+ xrcrg2 = 1
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ cigbacc = 0.245
+ wtvoff = -1.02826e-10
+ tnoimod = 0
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ capmod = 2
+ cigbinv = 0.006
+ wku0we = 1.5e-11
+ k2we = 5e-5
+ mobmod = 0
+ ijthsfwd = 0.01
+ dsub = 0.5
+ dtox = 3.91e-10
+ tvoff = 0.0027071394
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ xjbvd = 1
+ xjbvs = 1
+ version = 4.5
+ lk2we = 0.0
+ tempmod = 0
+ eta0 = 0.17962267
+ etab = -0.19577778
+ ijthsrev = 0.01
+ ku0we = -0.0007
+ aigbacc = 0.012071
+ beta0 = 13.32
+ leta0 = 4.8e-10
+ laigsd = 1.0132005e-13
+ ppclm = 0
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ aigbinv = 0.009974
+ ppdiblc2 = -7.3176658e-16
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ )

.model pch_sf_27 pmos (
+ level = 54
+ tvfbsdoff = 0.1
+ fnoimod = 1
+ scref = 1e-6
+ eigbinv = 1.1
+ rshg = 14.1
+ ltvoff = -3.7535707e-10
+ pigcd = 2.572
+ aigsd = 0.0063633912
+ lvoff = -1.1639377e-8
+ lvsat = -8.000000000000001e-6
+ lvth0 = 1.2906701e-9
+ ijthsfwd = 0.01
+ lku0we = 1.8e-11
+ delta = 0.018814
+ laigc = -5.5983746e-11
+ epsrox = 3.9
+ tnom = 25
+ rnoia = 0
+ rnoib = 0
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ cigbacc = 0.245
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ rdsmod = 0
+ igbmod = 1
+ pketa = 5.6398736e-15
+ ngate = 1.7e+20
+ wtvfbsdoff = 0
+ ijthsrev = 0.01
+ ngcon = 1
+ tnoimod = 0
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ wpclm = -1.1447315e-8
+ pbswgd = 0.8
+ pbswgs = 0.8
+ gbmin = 1e-12
+ cigbinv = 0.006
+ jswgd = 3.69e-13
+ ltvfbsdoff = 0
+ jswgs = 3.69e-13
+ igcmod = 1
+ wags = 3.4820603e-7
+ voff = -0.10461895
+ acde = 0.5
+ version = 4.5
+ ppdiblc2 = 9.4893758e-16
+ vsat = 91103.982
+ tempmod = 0
+ wint = 0
+ vth0 = -0.36807681999999997
+ wkt1 = 1.4552168e-8
+ wkt2 = 6.9668931e-9
+ wmax = 5.374e-7
+ aigc = 0.0068462496
+ wmin = 2.674e-7
+ aigbacc = 0.012071
+ ptvfbsdoff = 0
+ tvoff = 0.0026312893
+ wua1 = 1.777316e-16
+ wub1 = 1.5048515e-26
+ wuc1 = -3.1929257e-17
+ permod = 1
+ xjbvd = 1
+ xjbvs = 1
+ bigc = 0.0012521
+ wute = 6.965504e-8
+ lk2we = 0.0
+ wwlc = 0
+ pkvth0we = 0.0
+ aigbinv = 0.009974
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ ku0we = -0.0007
+ beta0 = 13.32
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ voffcv = -0.125
+ wpemod = 1
+ cigc = 0.15259
+ vfbsdoff = 0.01
+ leta0 = 4.8e-10
+ ppclm = 0
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ paramchk = 1
+ poxedge = 1
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ binunit = 2
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ tpbswg = 0.001
+ k2we = 5e-5
+ ijthdfwd = 0.01
+ dsub = 0.5
+ dtox = 3.91e-10
+ a0 = 2.4559917
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 72000
+ cf = 8.17e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.0065510297
+ k3 = -2.5823
+ em = 20000000.0
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ ll = 0
+ lw = 0
+ u0 = 0.010979968
+ w0 = 0
+ ua = 2.2475737e-10
+ ub = 1.3971204e-18
+ uc = 8.9671176e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ bigsd = 0.0003327
+ ptvoff = 6.0034078e-17
+ eta0 = 0.17962267
+ etab = -0.19577778
+ waigsd = 1.9297907e-12
+ wvoff = -2.3606869e-9
+ ijthdrev = 0.01
+ wvsat = 0.0034765009
+ diomod = 1
+ wvth0 = 1.0432152000000004e-9
+ lpdiblc2 = -1.0873556e-9
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ waigc = -6.0221967e-12
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.7086399999999997e-10
+ pku0we = 0.0
+ cjswgs = 1.7086399999999997e-10
+ lketa = -2.7133526e-8
+ xpart = 1
+ mjswgd = 0.95
+ mjswgs = 0.95
+ egidl = 0.001
+ tcjswg = 0.00128
+ pvfbsdoff = 0
+ lkvth0we = 3e-12
+ njtsswg = 6.489
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ acnqsmod = 0
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.012575691
+ pdiblcb = 0
+ rbodymod = 0
+ fprout = 200
+ xrcrg1 = 12
+ xrcrg2 = 1
+ pvoff = 1.5289261e-15
+ keta = 0.0057304489
+ cdscb = 0
+ cdscd = 0
+ pvsat = 0
+ bigbacc = 0.0054401
+ lags = 9.833094e-7
+ wk2we = 0.0
+ pvth0 = -2.4041799999999865e-18
+ wtvoff = -1.9743529e-10
+ drout = 0.56
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 6.6671111e-11
+ paigc = 6.5097646e-18
+ kt1l = 0
+ kvth0we = -0.00022
+ voffl = 0
+ wpdiblc2 = -1.8846129e-9
+ lintnoi = -5e-9
+ capmod = 2
+ lint = 6.5375218e-9
+ bigbinv = 0.00149
+ weta0 = -1.7424176e-8
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ wetab = 1.9534667e-8
+ wku0we = 1.5e-11
+ lkt1 = -3.8529349e-9
+ lkt2 = -2.567581e-9
+ lpclm = 0
+ lmax = 8.9908e-7
+ lmin = 4.4908e-7
+ mobmod = 0
+ lpe0 = 6.44e-8
+ lpeb = 0
+ cgidl = 1
+ minv = -0.33
+ lua1 = 1.3348283e-16
+ lub1 = 2.1611253e-25
+ luc1 = 5.928335e-17
+ ndep = 1e+18
+ lute = 1.2896693e-7
+ wkvth0we = 0.0
+ lwlc = 0
+ moin = 5.5538
+ pbswd = 0.9
+ pbsws = 0.9
+ ags = -0.056621626
+ nigc = 2.291
+ trnqsmod = 0
+ cjd = 0.001270624
+ cit = -8.7888889e-5
+ cjs = 0.001270624
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 1.0572421799999999e-8
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ pdits = 0
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ cigsd = 0.013281
+ nfactor = 1
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ la0 = -1.8333262e-7
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = -0.00064
+ pags = -2.41252e-13
+ kt1 = -0.20789546
+ kt2 = -0.0733757
+ lk2 = -8.954158000000004e-11
+ llc = 0
+ lln = 1
+ lu0 = -3.2154965000000003e-10
+ mjd = 0.335
+ mjs = 0.335
+ lua = -5.402342e-17
+ lub = -8.029291e-26
+ luc = -6.9221885e-17
+ lud = 0
+ ntox = 1.0
+ lwc = 0
+ lwl = 0
+ pcit = 8.000000000000001e-19
+ lwn = 1
+ pclm = 1.1689658
+ njd = 1.02
+ njs = 1.02
+ pa0 = -1.295362e-13
+ rgatemod = 0
+ nsd = 1e+20
+ pbd = 0.75
+ pk2we = 0.0
+ pat = 0
+ pbs = 0.75
+ pk2 = 6.34174e-16
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ tnjtsswg = 1
+ pu0 = -2.5304972e-16
+ prt = 0
+ pua = -1.1377853e-22
+ pub = 1.1787175e-31
+ puc = 2.8393052e-23
+ pud = 0
+ phin = 0.15
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 1.5353037e-9
+ ub1 = -2.5129786e-18
+ uc1 = 1.2019494e-10
+ tpb = 0.0016
+ tnoia = 0
+ wa0 = 1.4554629e-7
+ pkt1 = -1.0166873999999999e-14
+ pkt2 = -7.3243565e-16
+ ute = -1.2205289
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 2.3228278e-9
+ nigbacc = 10
+ wlc = 0
+ wln = 1
+ wu0 = 3.4013886e-10
+ xgl = -8.2e-9
+ xgw = 0
+ peta0 = 1.6e-17
+ wua = -1.1141771e-17
+ wub = -5.4878553e-26
+ wuc = -2.8229789e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ wketa = -8.9579586e-9
+ tpbsw = 0.0025
+ cjswd = 4.8144e-11
+ cjsws = 4.8144e-11
+ rbdb = 50
+ pua1 = -9.6760461e-23
+ prwb = 0
+ pub1 = 5.7312604e-33
+ prwg = 0
+ puc1 = -1.747778e-23
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ nigbinv = 2.171
+ pute = -4.8084303e-14
+ rdsw = 200
+ toxref = 3e-9
+ )

.model pch_sf_28 pmos (
+ level = 54
+ wtvfbsdoff = 0
+ lku0we = 1.8e-11
+ k2we = 5e-5
+ epsrox = 3.9
+ dsub = 0.5
+ dtox = 3.91e-10
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ ltvfbsdoff = 0
+ bigbacc = 0.0054401
+ rdsmod = 0
+ igbmod = 1
+ wkvth0we = 0.0
+ eta0 = 0.17962267
+ etab = -0.19577778
+ kvth0we = -0.00022
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ trnqsmod = 0
+ pbswgd = 0.8
+ lintnoi = -5e-9
+ pbswgs = 0.8
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ pvoff = -2.4654209e-16
+ igcmod = 1
+ cdscb = 0
+ cdscd = 0
+ pvsat = 0
+ wk2we = 0.0
+ pvth0 = -5.767691400000001e-16
+ ptvfbsdoff = 0
+ drout = 0.56
+ paigc = -3.9499473e-18
+ voffl = 0
+ rgatemod = 0
+ tnjtsswg = 1
+ weta0 = -1.7424176e-8
+ wetab = 1.9534667e-8
+ lpclm = 0
+ cgidl = 1
+ permod = 1
+ ags = -1.2539967
+ nfactor = 1
+ cjd = 0.001270624
+ cit = -0.00036538451
+ cjs = 0.001270624
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 1.38228675e-8
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ pbswd = 0.9
+ pbsws = 0.9
+ voffcv = -0.125
+ wpemod = 1
+ la0 = -4.7253353e-7
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = -0.00064
+ kt1 = -0.16257215
+ kt2 = -0.066291072
+ lk2 = 6.0447077e-10
+ llc = -1.18e-13
+ lln = 0.7
+ lu0 = -5.4210454e-10
+ keta = -0.0061234738
+ mjd = 0.335
+ mjs = 0.335
+ lua = -1.0290148e-16
+ lub = -5.3060964e-27
+ luc = -4.0794824e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pdits = 0
+ pa0 = 9.7298482e-15
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ cigsd = 0.013281
+ pk2 = -2.0891363e-16
+ nigbacc = 10
+ lags = 1.5101544e-6
+ pu0 = 1.1540053e-17
+ dvt0w = 0
+ dvt1w = 0
+ prt = 0
+ dvt2w = 0
+ pua = -1.3867635e-23
+ pub = 2.1855871e-32
+ puc = -2.7646346e-24
+ pud = 0
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 1.8876918e-10
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 1.7313241e-9
+ ub1 = -1.3316629e-18
+ uc1 = 2.2670111e-10
+ kt1l = 0
+ tpb = 0.0016
+ wa0 = -1.7096745e-7
+ ute = -0.86054925
+ web = 6628.3
+ wec = -16935.0
+ pk2we = 0.0
+ wk2 = 4.238936e-9
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ wlc = 0
+ wln = 1
+ wu0 = -2.6120153e-10
+ xgl = -8.2e-9
+ xgw = 0
+ wua = -2.3821198e-16
+ wub = 1.6333936e-25
+ wuc = 4.2583136e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ nigbinv = 2.171
+ lint = 9.7879675e-9
+ tpbswg = 0.001
+ lkt1 = -2.3795191999999997e-8
+ lkt2 = -5.6848171e-9
+ lmax = 4.4908e-7
+ tnoia = 0
+ lmin = 2.1577e-7
+ lpe0 = 6.44e-8
+ ijthsfwd = 0.01
+ lpeb = 0
+ peta0 = 1.6e-17
+ wketa = -7.8373297e-10
+ minv = -0.33
+ tpbsw = 0.0025
+ lua1 = 4.723388e-17
+ lub1 = -3.0366637e-25
+ luc1 = 1.2420632e-17
+ ptvoff = 5.0195791e-17
+ cjswd = 4.8144e-11
+ cjsws = 4.8144e-11
+ ndep = 1e+18
+ fnoimod = 1
+ mjswd = 0.01
+ lute = -2.9424109e-8
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ waigsd = 1.9297907e-12
+ lwlc = 0
+ eigbinv = 1.1
+ moin = 5.5538
+ ijthsrev = 0.01
+ nigc = 2.291
+ diomod = 1
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.7086399999999997e-10
+ pku0we = 0.0
+ cjswgs = 1.7086399999999997e-10
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ tvfbsdoff = 0.1
+ pags = -3.3771496e-13
+ scref = 1e-6
+ a0 = 3.1132665
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 72000
+ cf = 8.17e-11
+ ntox = 1.0
+ mjswgd = 0.95
+ ef = 1.15
+ mjswgs = 0.95
+ k1 = 0.30425
+ k2 = -0.0081283305
+ k3 = -2.5823
+ pcit = -8.471640299999999e-18
+ em = 20000000.0
+ ppdiblc2 = -3.8737293e-16
+ pclm = 1.1689658
+ pigcd = 2.572
+ cigbacc = 0.245
+ ll = -1.18e-13
+ aigsd = 0.0063633912
+ lw = 0
+ u0 = 0.01148123
+ w0 = 0
+ ua = 3.3584387e-10
+ ub = 1.2266958e-18
+ uc = -5.8379738e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ tcjswg = 0.00128
+ lvoff = -4.2658924e-9
+ phin = 0.15
+ tnoimod = 0
+ lvsat = -8.000000000000001e-6
+ pkt1 = 6.8755166e-15
+ pkt2 = 2.2627554e-16
+ lvth0 = 4.8053579e-9
+ cigbinv = 0.006
+ delta = 0.018814
+ laigc = -1.8017042e-11
+ wvfbsdoff = 0
+ rnoia = 0
+ rnoib = 0
+ lvfbsdoff = 0
+ rbdb = 50
+ pua1 = -2.7108228e-23
+ pkvth0we = 0.0
+ prwb = 0
+ pub1 = 7.1177686e-32
+ prwg = 0
+ puc1 = 8.7727027e-25
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ pketa = 2.0432143e-15
+ version = 4.5
+ ngate = 1.7e+20
+ pute = 1.6065563e-14
+ fprout = 200
+ rdsw = 200
+ ngcon = 1
+ tempmod = 0
+ wpclm = -1.1447315e-8
+ xrcrg1 = 12
+ xrcrg2 = 1
+ vfbsdoff = 0.01
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ aigbacc = 0.012071
+ wtvoff = -1.7507555e-10
+ paramchk = 1
+ rshg = 14.1
+ capmod = 2
+ aigbinv = 0.009974
+ wku0we = 1.5e-11
+ mobmod = 0
+ ijthdfwd = 0.01
+ tvoff = 0.002323434
+ tnom = 25
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ poxedge = 1
+ ijthdrev = 0.01
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = 4.8e-10
+ lpdiblc2 = 4.7505822e-10
+ binunit = 2
+ ppclm = 0
+ wags = 5.6744004e-7
+ wcit = 2.107191e-11
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ voff = -0.12137687
+ acde = 0.5
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ vsat = 91103.982
+ wint = 0
+ vth0 = -0.37606475
+ wkt1 = -2.4180539e-8
+ wkt2 = 4.7880041e-9
+ wmax = 5.374e-7
+ dmcgt = 0
+ aigc = 0.0067599617
+ wmin = 2.674e-7
+ tcjsw = 9.34e-5
+ lkvth0we = 3e-12
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ wua1 = 1.9431072e-17
+ wub1 = -1.3369336e-25
+ wuc1 = -7.3645279e-17
+ acnqsmod = 0
+ bigc = 0.0012521
+ bigsd = 0.0003327
+ wute = -7.6140111e-8
+ wwlc = 0
+ wvoff = 1.674468e-9
+ toxref = 3e-9
+ rbodymod = 0
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ wvsat = 0.0034765009
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ wvth0 = 2.3485901000000005e-9
+ cigc = 0.15259
+ waigc = 1.7749876e-11
+ njtsswg = 6.489
+ lketa = -2.19178e-8
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ ltvoff = -2.3990075e-10
+ xpart = 1
+ ckappad = 0.6
+ wpdiblc2 = 1.1524564e-9
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.0090247504
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ pdiblcb = 0
+ egidl = 0.001
+ pvfbsdoff = 0
+ )

.model pch_sf_29 pmos (
+ level = 54
+ ijthdrev = 0.01
+ ngcon = 1
+ pbswgd = 0.8
+ pbswgs = 0.8
+ wpclm = -1.2079184e-7
+ aigbinv = 0.009974
+ nigc = 2.291
+ igcmod = 1
+ lpdiblc2 = -1.1954251e-9
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ ntox = 1.0
+ pcit = -7.329839099999999e-18
+ pclm = 1.5407845
+ poxedge = 1
+ phin = 0.15
+ lkvth0we = 3e-12
+ pkt1 = -1.17482e-15
+ pkt2 = -1.4992738e-15
+ binunit = 2
+ permod = 1
+ tvoff = 0.00085372815
+ acnqsmod = 0
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ rbdb = 50
+ pua1 = 1.9617826e-23
+ prwb = 0
+ pub1 = -3.1346313e-32
+ prwg = 0
+ puc1 = 1.1713402e-23
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ rbodymod = 0
+ voffcv = -0.125
+ wpemod = 1
+ rdsw = 200
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = 4.8e-10
+ ppclm = 2.3071337e-14
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ rshg = 14.1
+ wpdiblc2 = -7.3926191e-10
+ tpbswg = 0.001
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ njtsswg = 6.489
+ ptvoff = -3.132788e-17
+ tnom = 25
+ bigsd = 0.0003327
+ waigsd = 1.9297907e-12
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ wkvth0we = 0.0
+ wvoff = 3.1859801e-10
+ diomod = 1
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.016941733
+ trnqsmod = 0
+ pdiblcb = 0
+ wvsat = 0.0032472346
+ pditsd = 0
+ wvth0 = -2.8069424999999994e-9
+ pditsl = 0
+ cjswgd = 1.7086399999999997e-10
+ pku0we = 0.0
+ cjswgs = 1.7086399999999997e-10
+ waigc = -1.7260908e-11
+ wags = -1.0331048e-6
+ wcit = 1.566053e-11
+ lketa = 7.1935383e-9
+ voff = -0.13201276
+ mjswgd = 0.95
+ mjswgs = 0.95
+ bigbacc = 0.0054401
+ acde = 0.5
+ xpart = 1
+ rgatemod = 0
+ tcjswg = 0.00128
+ vsat = 91523.884
+ wint = 0
+ tnjtsswg = 1
+ vth0 = -0.37362236
+ pvfbsdoff = 0
+ kvth0we = -0.00022
+ egidl = 0.001
+ wkt1 = 1.3972715e-8
+ wkt2 = 1.2965963e-8
+ wmax = 5.374e-7
+ aigc = 0.0067957378
+ wmin = 2.674e-7
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ wua1 = -2.0201942e-16
+ wub1 = 3.5220237e-25
+ wuc1 = -1.2500135e-16
+ bigc = 0.0012521
+ wwlc = 0
+ fprout = 200
+ cdsc = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ a0 = 1.1444157
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ at = 108550.2
+ xtid = 3
+ cf = 8.17e-11
+ xtis = 3
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.025395241
+ k3 = -2.5823
+ em = 20000000.0
+ ll = -1.18e-13
+ lw = 0
+ u0 = 0.0098417592
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ w0 = 0
+ ua = -3.1599722e-11
+ ub = 1.4008434e-18
+ uc = -1.6299488e-10
+ ud = 0
+ cigc = 0.15259
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ pvoff = 3.9546471e-17
+ wtvoff = 2.1129256e-10
+ cdscb = 0
+ cdscd = 0
+ pvsat = 4.83709e-11
+ wk2we = 0.0
+ pvth0 = 5.1104824e-16
+ drout = 0.56
+ paigc = 3.4373281e-18
+ nfactor = 1
+ capmod = 2
+ voffl = 0
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ wku0we = 1.5e-11
+ dmdg = 0
+ weta0 = -1.7424176e-8
+ wetab = 1.9534667e-8
+ mobmod = 0
+ ags = 5.9031333
+ lpclm = -7.8453093e-8
+ cjd = 0.001270624
+ cit = 0.00015305446
+ cjs = 0.001270624
+ clc = 1e-7
+ cle = 0.6
+ k2we = 5e-5
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 1.38228675e-8
+ ijthsfwd = 0.01
+ k3b = 2.1176
+ dsub = 0.5
+ cgidl = 1
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ dtox = 3.91e-10
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ nigbacc = 10
+ la0 = -5.7105222e-8
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = -0.0083520921
+ kt1 = -0.27233533
+ kt2 = -0.10755274
+ lk2 = 4.2477889e-9
+ eta0 = 0.17962267
+ llc = -1.18e-13
+ lln = 0.7
+ lu0 = -1.961763e-10
+ etab = -0.19577778
+ mjd = 0.335
+ mjs = 0.335
+ lua = -2.5370884e-17
+ lub = -4.2051244e-26
+ luc = 1.7994313e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ pbswd = 0.9
+ pbsws = 0.9
+ njd = 1.02
+ njs = 1.02
+ pa0 = -3.159814e-15
+ ijthsrev = 0.01
+ nsd = 1e+20
+ pbd = 0.75
+ pat = -4.5415452e-10
+ pbs = 0.75
+ pk2 = -2.0710507e-16
+ pu0 = 4.0684676e-18
+ prt = 0
+ pua = 6.5898257e-24
+ pub = -4.9701536e-33
+ puc = -7.066739e-24
+ pud = 0
+ nigbinv = 2.171
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 2.8369875e-9
+ ub1 = -4.0389099e-18
+ uc1 = 4.2708978e-10
+ tpb = 0.0016
+ wa0 = -1.0988104e-7
+ pdits = 0
+ ute = -1
+ wat = 0.0021523911
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 4.2303646e-9
+ cigsd = 0.013281
+ wlc = 0
+ wln = 1
+ wu0 = -2.2579117e-10
+ xgl = -8.2e-9
+ xgw = 0
+ wua = -3.3516677e-16
+ dvt0w = 0
+ wub = 2.9047692e-25
+ wuc = 6.2972257e-17
+ wud = 0
+ dvt1w = 0
+ dvt2w = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ ppdiblc2 = 1.1779633e-17
+ pk2we = 0.0
+ fnoimod = 1
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ eigbinv = 1.1
+ tnoia = 0
+ peta0 = 1.6e-17
+ wketa = 1.4826965e-8
+ tpbsw = 0.0025
+ cjswd = 4.8144e-11
+ cjsws = 4.8144e-11
+ pkvth0we = 0.0
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ toxref = 3e-9
+ cigbacc = 0.245
+ vfbsdoff = 0.01
+ tnoimod = 0
+ keta = -0.1440919
+ tvfbsdoff = 0.1
+ wtvfbsdoff = 0
+ cigbinv = 0.006
+ ltvoff = 7.0207177e-11
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 7.937856e-11
+ paramchk = 1
+ scref = 1e-6
+ kt1l = 0
+ pigcd = 2.572
+ aigsd = 0.0063633912
+ ltvfbsdoff = 0
+ version = 4.5
+ lvoff = -2.0217201e-9
+ lint = 9.7879675e-9
+ tempmod = 0
+ lkt1 = -6.351622e-10
+ lkt2 = 3.021395e-9
+ lku0we = 1.8e-11
+ lmax = 2.1577e-7
+ lvsat = -9.65914e-5
+ lmin = 9e-8
+ epsrox = 3.9
+ lvth0 = 4.2900147e-9
+ lpe0 = 6.44e-8
+ ijthdfwd = 0.01
+ lpeb = 0
+ delta = 0.018814
+ laigc = -2.5565813e-11
+ aigbacc = 0.012071
+ wvfbsdoff = 0
+ rdsmod = 0
+ lvfbsdoff = 0
+ minv = -0.33
+ rnoia = 0
+ rnoib = 0
+ lua1 = -1.8606111e-16
+ lub1 = 2.6756274e-25
+ luc1 = -2.9861377e-17
+ igbmod = 1
+ ndep = 1e+18
+ ptvfbsdoff = 0
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ lwlc = 0
+ pketa = -1.250643e-15
+ ngate = 1.7e+20
+ moin = 5.5538
+ )

.model pch_sf_30 pmos (
+ level = 54
+ ijthdrev = 0.01
+ ngcon = 1
+ pbswgd = 0.8
+ pbswgs = 0.8
+ wpclm = 4.9341412e-7
+ aigbinv = 0.009974
+ nigc = 2.291
+ igcmod = 1
+ lpdiblc2 = 0
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ ntox = 1.0
+ pcit = -5.378864999999999e-18
+ pclm = 0.08631615
+ paigsd = 8.4526218e-25
+ poxedge = 1
+ phin = 0.15
+ lkvth0we = 3e-12
+ pkt1 = -1.6724191e-15
+ pkt2 = 2.1480498e-17
+ binunit = 2
+ permod = 1
+ tvoff = 0.0012365685
+ acnqsmod = 0
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ rbdb = 50
+ pua1 = 4.1792962e-25
+ prwb = 0
+ pub1 = 6.1746384e-33
+ prwg = 0
+ puc1 = 2.9246063e-24
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ rbodymod = 0
+ voffcv = -0.125
+ wpemod = 1
+ rdsw = 200
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = -8.0858832e-9
+ letab = 1.7579973e-8
+ ppclm = -3.4664022e-14
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ rshg = 14.1
+ wpdiblc2 = -6.1394667e-10
+ tpbswg = 0.001
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ njtsswg = 6.489
+ ptvoff = 2.0376593e-17
+ tnom = 25
+ bigsd = 0.0003327
+ waigsd = 1.9297817e-12
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ wkvth0we = 0.0
+ wvoff = -2.8254962e-9
+ diomod = 1
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.0042244444
+ trnqsmod = 0
+ pdiblcb = 0
+ wvsat = 0.017016245
+ pditsd = 0
+ wvth0 = -1.6431860999999996e-9
+ pditsl = 0
+ cjswgd = 1.7086399999999997e-10
+ pku0we = 0.0
+ cjswgs = 1.7086399999999997e-10
+ waigc = 7.1461687e-12
+ wags = -1.0331048e-6
+ wcit = -5.09452e-12
+ lketa = -1.1878561e-8
+ voff = -0.12098873
+ mjswgd = 0.95
+ mjswgs = 0.95
+ bigbacc = 0.0054401
+ acde = 0.5
+ xpart = 1
+ rgatemod = 0
+ tcjswg = 0.00128
+ vsat = 62231.739
+ wint = 0
+ tnjtsswg = 1
+ vth0 = -0.31746471
+ pvfbsdoff = 0
+ kvth0we = -0.00022
+ egidl = 0.001
+ wkt1 = 1.9266322e-8
+ wkt2 = -3.2122744e-9
+ wmax = 5.374e-7
+ aigc = 0.0067006504
+ wmin = 2.674e-7
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ wua1 = 2.2347963e-18
+ wub1 = -4.6956688e-26
+ wuc1 = -3.1503526e-17
+ bigc = 0.0012521
+ wwlc = 0
+ fprout = 200
+ cdsc = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ a0 = 3.9744452
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ at = 69068.642
+ xtid = 3
+ cf = 8.17e-11
+ xtis = 3
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.022825095
+ k3 = -2.5823
+ em = 20000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.0040056963
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ w0 = 0
+ ua = -9.2439852e-11
+ ub = -1.6232125e-18
+ uc = 5.3507127e-11
+ ud = 0
+ cigc = 0.15259
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ pvoff = 3.3509132e-16
+ wtvoff = -3.3875503e-10
+ cdscb = 0
+ cdscd = 0
+ pvsat = -1.2459161e-9
+ wk2we = 0.0
+ pvth0 = 4.0165514e-16
+ drout = 0.56
+ paigc = 1.1430629e-18
+ nfactor = 1
+ capmod = 2
+ voffl = 0
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ wku0we = 1.5e-11
+ dmdg = 0
+ weta0 = -5.4791839e-8
+ wetab = 4.6876459e-8
+ mobmod = 0
+ ags = 5.9031333
+ lpclm = 5.8266931e-8
+ cjd = 0.001270624
+ cit = -0.00018033605
+ cjs = 0.001270624
+ clc = 1e-7
+ cle = 0.6
+ k2we = 5e-5
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 4.0349e-9
+ ijthsfwd = 0.01
+ k3b = 2.1176
+ dsub = 0.5
+ cgidl = 1
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ dtox = 3.91e-10
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ nigbacc = 10
+ la0 = -3.23128e-7
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = -0.0046408257
+ kt1 = -0.32608492
+ kt2 = -0.08284588
+ lk2 = 4.006195200000001e-9
+ eta0 = 0.27074908
+ llc = 0
+ lln = 1
+ lu0 = 3.5241361999999997e-10
+ etab = -0.38279877
+ mjd = 0.335
+ mjs = 0.335
+ lua = -1.9651912e-17
+ lub = 2.4221001e-25
+ luc = -2.356876e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ pbswd = 0.9
+ pbsws = 0.9
+ njd = 1.02
+ njs = 1.02
+ pa0 = 9.1746422e-14
+ laigsd = -3.0625433e-18
+ ijthsrev = 0.01
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 6.7620954e-11
+ pbs = 0.75
+ pk2 = 2.5170462e-16
+ pu0 = -8.2666616e-17
+ prt = 0
+ pua = 3.032424e-23
+ pub = -9.6166295e-32
+ puc = -2.0363205e-24
+ pud = 0
+ nigbinv = 2.171
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = -2.7998083e-10
+ ub1 = 8.7083504e-19
+ uc1 = 1.8820988e-11
+ tpb = 0.0016
+ wa0 = -1.1195219e-6
+ pdits = 0
+ ute = -1
+ wat = -0.0033984119
+ web = 6628.3
+ wec = -16935.0
+ wk2 = -6.5058945e-10
+ cigsd = 0.013281
+ wlc = 0
+ wln = 1
+ wu0 = 6.9692249e-10
+ xgl = -8.2e-9
+ xgw = 0
+ wua = -5.8766054e-16
+ dvt0w = 0
+ wub = 1.2606486e-24
+ wuc = 9.4571662e-18
+ wud = 0
+ dvt1w = 0
+ dvt2w = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ ppdiblc2 = 0
+ pk2we = 0.0
+ fnoimod = 1
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ eigbinv = 1.1
+ tnoia = 0
+ peta0 = 3.5285603e-15
+ petab = -2.5701285e-15
+ wketa = -3.6489897e-8
+ tpbsw = 0.0025
+ cjswd = 4.8144e-11
+ cjsws = 4.8144e-11
+ pkvth0we = 0.0
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ toxref = 3e-9
+ cigbacc = 0.245
+ vfbsdoff = 0.01
+ tnoimod = 0
+ keta = 0.058802768
+ tvfbsdoff = 0.1
+ wtvfbsdoff = 0
+ cigbinv = 0.006
+ ltvoff = 3.4220189e-11
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 1.1071727e-10
+ paramchk = 1
+ scref = 1e-6
+ kt1l = 0
+ pigcd = 2.572
+ aigsd = 0.0063633912
+ ltvfbsdoff = 0
+ version = 4.5
+ lvoff = -3.0579783e-9
+ lint = 0
+ tempmod = 0
+ lkt1 = 4.4172999e-9
+ lkt2 = 6.989501e-10
+ lku0we = 1.8e-11
+ lmax = 9e-8
+ lvsat = 0.0026568702999999996
+ lmin = 5.4e-8
+ epsrox = 3.9
+ lvth0 = -9.888048e-10
+ lpe0 = 6.44e-8
+ ijthdfwd = 0.01
+ lpeb = 0
+ delta = 0.018814
+ laigc = -1.6627591e-11
+ aigbacc = 0.012071
+ wvfbsdoff = 0
+ rdsmod = 0
+ lvfbsdoff = 0
+ minv = -0.33
+ rnoia = 0
+ rnoib = 0
+ lua1 = 1.0693391e-16
+ lub1 = -1.9395329e-25
+ luc1 = 8.5158894e-18
+ igbmod = 1
+ ndep = 1e+18
+ ptvfbsdoff = 0
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ lwlc = 0
+ pketa = 3.573142e-15
+ ngate = 1.7e+20
+ moin = 5.5538
+ )

.model pch_sf_31 pmos (
+ level = 54
+ paigc = -3.8652128e-18
+ voff = -0.11425646
+ nigbacc = 10
+ ags = 5.9031333
+ acde = 0.5
+ ppdiblc2 = 0
+ voffl = 0
+ cjd = 0.001270624
+ cit = -0.0023632098
+ cjs = 0.001270624
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ vsat = 205509.49
+ dlc = 4.0349e-9
+ wint = 0
+ k3b = 2.1176
+ vth0 = -0.29741972
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ weta0 = 4.5793198e-8
+ wkt1 = -9.053012e-8
+ wkt2 = -4.5663135e-8
+ wetab = 2.1214781e-8
+ wmax = 5.374e-7
+ aigc = 0.0065523001
+ wmin = 2.674e-7
+ lpclm = -1.6067206e-7
+ permod = 1
+ nigbinv = 2.171
+ la0 = 2.2449695e-9
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = -0.00158527867
+ kt1 = -0.078489325
+ kt2 = 0.051187672
+ lk2 = 5.103110100000001e-9
+ llc = 0
+ lln = 1
+ cgidl = 1
+ lu0 = -6.406920299999999e-10
+ mjd = 0.335
+ mjs = 0.335
+ lua = -5.2618623e-17
+ lub = -3.080728e-25
+ luc = -2.0280652e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ wua1 = 2.8402308e-15
+ njs = 1.02
+ wub1 = -3.9062366e-24
+ wuc1 = 2.0276364e-16
+ pa0 = -4.432942e-14
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 1.8264736e-9
+ pbs = 0.75
+ pk2 = -1.1995676e-16
+ pu0 = 2.2577126e-16
+ bigc = 0.0012521
+ prt = 0
+ pua = 1.5923531e-23
+ pub = 9.2000466e-32
+ puc = 3.3504384e-24
+ pud = 0
+ wwlc = 0
+ pkvth0we = 0.0
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = -3.345352e-9
+ ub1 = 3.9080279e-18
+ uc1 = 1.4308247e-10
+ tpb = 0.0016
+ voffcv = -0.125
+ wpemod = 1
+ pbswd = 0.9
+ pbsws = 0.9
+ wa0 = 1.2266134e-6
+ cdsc = 0
+ ute = -1
+ wat = -0.033723458
+ web = 6628.3
+ wec = -16935.0
+ fnoimod = 1
+ wk2 = 5.7573654e-9
+ wlc = 0
+ cgbo = 0
+ wln = 1
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ wu0 = -4.6209719e-9
+ xtid = 3
+ xgl = -8.2e-9
+ xtis = 3
+ xgw = 0
+ wua = -3.3937245e-16
+ wub = -1.9836059e-24
+ wuc = -8.3417988e-17
+ wud = 0
+ eigbinv = 1.1
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ vfbsdoff = 0.01
+ cigc = 0.15259
+ pdits = 0
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ paramchk = 1
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ tpbswg = 0.001
+ cigbacc = 0.245
+ tnoia = 0
+ k2we = 5e-5
+ tnoimod = 0
+ ijthdfwd = 0.01
+ peta0 = -2.3053718000000003e-15
+ dsub = 0.5
+ petab = -1.0817512e-15
+ dtox = 3.91e-10
+ wketa = 7.0696889e-8
+ ptvoff = -1.3332507e-17
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ tpbsw = 0.0025
+ waigsd = 1.9297962e-12
+ cigbinv = 0.006
+ cjswd = 4.8144e-11
+ cjsws = 4.8144e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ eta0 = 0.012687945
+ etab = -0.23454709
+ diomod = 1
+ ijthdrev = 0.01
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.7086399999999997e-10
+ pku0we = 0.0
+ version = 4.5
+ cjswgs = 1.7086399999999997e-10
+ lpdiblc2 = 0
+ tempmod = 0
+ tvfbsdoff = 0.1
+ aigbacc = 0.012071
+ mjswgd = 0.95
+ mjswgs = 0.95
+ scref = 1e-6
+ tcjswg = 0.00128
+ pigcd = 2.572
+ aigsd = 0.0063633912
+ lvoff = -3.4484499e-9
+ lkvth0we = 3e-12
+ aigbinv = 0.009974
+ lvsat = -0.0056532393000000005
+ lvth0 = -2.1514143e-9
+ delta = 0.018814
+ wvfbsdoff = 0
+ laigc = -8.0232722e-12
+ lvfbsdoff = 0
+ rnoia = 0
+ rnoib = 0
+ acnqsmod = 0
+ fprout = 200
+ pketa = -2.6436916e-15
+ ngate = 1.7e+20
+ xrcrg1 = 12
+ xrcrg2 = 1
+ rbodymod = 0
+ ngcon = 1
+ wpclm = -6.9641486e-7
+ poxedge = 1
+ gbmin = 1e-12
+ wtvoff = 2.4243635e-10
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ keta = -0.44725926
+ binunit = 2
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 2.3732395e-10
+ capmod = 2
+ kt1l = 0
+ wku0we = 1.5e-11
+ wpdiblc2 = -6.1394667e-10
+ mobmod = 0
+ lint = 0
+ lkt1 = -9.943245e-9
+ lkt2 = -7.0749959e-9
+ lmax = 5.4e-8
+ lmin = 4.5e-8
+ a0 = -1.6354335
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 16386.797
+ cf = 8.17e-11
+ lpe0 = 6.44e-8
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.041737421
+ k3 = -2.5823
+ em = 20000000.0
+ lpeb = 0
+ ll = 0
+ lw = 0
+ u0 = 0.021128207
+ w0 = 0
+ tvoff = 0.0019328761
+ ua = 4.7595173e-10
+ ub = 7.8644222e-18
+ uc = 4.7837975e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ minv = -0.33
+ xjbvd = 1
+ xjbvs = 1
+ lua1 = 2.8472544e-16
+ lub1 = -3.7011047e-25
+ lk2we = 0.0
+ luc1 = 1.3087235e-18
+ ndep = 1e+18
+ wkvth0we = 0.0
+ lwlc = 0
+ moin = 5.5538
+ ku0we = -0.0007
+ trnqsmod = 0
+ nigc = 2.291
+ beta0 = 13.32
+ leta0 = 6.8816629e-9
+ letab = 8.9813755e-9
+ ppclm = 3.4346058e-14
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ njtsswg = 6.489
+ ntox = 1.0
+ pcit = -1.682461e-17
+ pclm = 3.8611263
+ rgatemod = 0
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ tnjtsswg = 1
+ dmcgt = 0
+ ckappad = 0.6
+ phin = 0.15
+ ckappas = 0.6
+ tcjsw = 9.34e-5
+ pdiblc1 = 0
+ pdiblc2 = 0.0042244444
+ pdiblcb = 0
+ pkt1 = 4.6957745e-15
+ pkt2 = 2.4836304e-15
+ bigsd = 0.0003327
+ toxref = 3e-9
+ rbdb = 50
+ pua1 = -1.6418584e-22
+ prwb = 0
+ pub1 = 2.3001287e-31
+ prwg = 0
+ puc1 = -1.0662889e-23
+ wtvfbsdoff = 0
+ bigbacc = 0.0054401
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ wvoff = 3.9335999e-9
+ rdsw = 200
+ wvsat = -0.031328619
+ kvth0we = -0.00022
+ ltvfbsdoff = 0
+ wvth0 = 1.3302981e-8
+ waigc = 9.3495749e-11
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ ltvoff = -6.1656569e-12
+ lketa = 1.7473037e-8
+ xpart = 1
+ rshg = 14.1
+ pvfbsdoff = 0
+ egidl = 0.001
+ ptvfbsdoff = 0
+ lku0we = 1.8e-11
+ epsrox = 3.9
+ ijthsfwd = 0.01
+ rdsmod = 0
+ igbmod = 1
+ tnom = 25
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ nfactor = 1
+ pbswgd = 0.8
+ pbswgs = 0.8
+ ijthsrev = 0.01
+ igcmod = 1
+ pvoff = -5.6936248e-17
+ cdscb = 0
+ cdscd = 0
+ wags = -1.0331048e-6
+ pvsat = 1.5580861e-9
+ wk2we = 0.0
+ pvth0 = -4.6522254e-16
+ wcit = 1.9224593e-10
+ drout = 0.56
+ )

.model pch_sf_32 pmos (
+ level = 54
+ tvoff = 0.0050068134
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ voffcv = -0.125
+ wpemod = 1
+ njtsswg = 6.489
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = 3.1914638e-9
+ ckappad = 0.6
+ letab = 1.8240871e-9
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.0042244444
+ pdiblcb = 0
+ keta = -0.10111506
+ ppclm = 1.7398739e-15
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = -2.0839499999999998e-11
+ kt1l = 0
+ tpbswg = 0.001
+ bigbacc = 0.0054401
+ lint = 0
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ lkt1 = -1.2929032e-8
+ lkt2 = 2.2261728e-10
+ lmax = 4.5e-8
+ kvth0we = -0.00022
+ lmin = 3.6e-8
+ lpe0 = 6.44e-8
+ ijthsfwd = 0.01
+ lpeb = 0
+ ptvoff = 3.2244316e-17
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ waigsd = 1.9257033e-12
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ minv = -0.33
+ bigsd = 0.0003327
+ lua1 = -1.7116539e-16
+ lub1 = 1.8549471e-25
+ luc1 = 2.2025561e-17
+ ndep = 1e+18
+ diomod = 1
+ lwlc = 0
+ wvoff = 1.094003e-8
+ moin = 5.5538
+ ijthsrev = 0.01
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.7086399999999997e-10
+ pku0we = 0.0
+ cjswgs = 1.7086399999999997e-10
+ nigc = 2.291
+ wvsat = -0.018712604
+ wvth0 = 1.7742333e-8
+ waigc = 1.753535e-10
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ mjswgd = 0.95
+ mjswgs = 0.95
+ lketa = 5.1197136e-10
+ tcjswg = 0.00128
+ xpart = 1
+ ntox = 1.0
+ ppdiblc2 = 0
+ pcit = 1.2234904e-16
+ pclm = 0.85281474
+ pvfbsdoff = 0
+ nfactor = 1
+ egidl = 0.001
+ phin = 0.15
+ pkt1 = 2.4784659999999998e-15
+ pkt2 = -1.2154904e-16
+ fprout = 200
+ pkvth0we = 0.0
+ rbdb = 50
+ pua1 = 5.9435365e-23
+ prwb = 0
+ pub1 = -6.8901825e-32
+ prwg = 0
+ puc1 = -3.4884574e-24
+ xrcrg1 = 12
+ xrcrg2 = 1
+ nigbacc = 10
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ rdsw = 200
+ wtvoff = -6.8770288e-10
+ vfbsdoff = 0.01
+ pvoff = -4.0025133e-16
+ ags = 5.9031333
+ nigbinv = 2.171
+ cdscb = 0
+ cdscd = 0
+ cjd = 0.001270624
+ cit = 0.0029054321
+ cjs = 0.001270624
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ pvsat = 9.3990127e-10
+ dlc = 4.0349e-9
+ wk2we = 0.0
+ pvth0 = -6.827508000000001e-16
+ k3b = 2.1176
+ dwb = 0
+ drout = 0.56
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ capmod = 2
+ paramchk = 1
+ paigc = -7.8762427e-18
+ wku0we = 1.5e-11
+ rshg = 14.1
+ voffl = 0
+ la0 = -2.1218621e-7
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0.009868083
+ mobmod = 0
+ kt1 = -0.017554887
+ kt2 = -0.09774321
+ lk2 = 3.737225800000001e-9
+ llc = 0
+ lln = 1
+ lu0 = -2.427917e-10
+ mjd = 0.335
+ mjs = 0.335
+ lua = 4.1444844e-17
+ lub = -1.5666965e-25
+ luc = -1.4956542e-17
+ lud = 0
+ lwc = 0
+ weta0 = 6.9541382e-9
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ wetab = -5.613608e-9
+ njs = 1.02
+ pa0 = 5.0455005e-14
+ fnoimod = 1
+ nsd = 1e+20
+ pbd = 0.75
+ pat = -2.4847929e-9
+ pbs = 0.75
+ pk2 = 3.3742201e-16
+ lpclm = -1.3264792e-8
+ pu0 = 1.5059926e-16
+ eigbinv = 1.1
+ prt = 0
+ pua = 9.2877876e-24
+ pub = 3.2782262e-32
+ puc = 3.1614905e-24
+ pud = 0
+ ijthdfwd = 0.01
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 5.9585425e-9
+ ub1 = -7.4308533e-18
+ uc1 = -2.7971012e-10
+ cgidl = 1
+ tpb = 0.0016
+ wa0 = -7.0776268e-7
+ ute = -1
+ wat = 0.054261574
+ web = 6628.3
+ wec = -16935.0
+ wk2 = -3.5768953e-9
+ wlc = 0
+ wln = 1
+ wu0 = -3.0868494e-9
+ tnom = 25
+ xgl = -8.2e-9
+ xgw = 0
+ wua = -2.0394912e-16
+ wub = -7.7507108e-25
+ wuc = -7.9561907e-17
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ laigsd = -3.6731852e-16
+ pbswd = 0.9
+ pbsws = 0.9
+ ijthdrev = 0.01
+ cigbacc = 0.245
+ lpdiblc2 = 0
+ pdits = 0
+ wags = -1.0331048e-6
+ cigsd = 0.013281
+ tnoimod = 0
+ dvt0w = 0
+ dvt1w = 0
+ wcit = -2.6480326e-9
+ dvt2w = 0
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ a0 = 2.7407131
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = -217355.29
+ cf = 8.17e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.013862232
+ k3 = -2.5823
+ em = 20000000.0
+ voff = -0.14966725
+ ll = 0
+ lw = 0
+ u0 = 0.013007793
+ w0 = 0
+ cigbinv = 0.006
+ acde = 0.5
+ ua = -1.4437109e-9
+ ub = 4.7745619e-18
+ uc = 3.1168444e-10
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ vsat = 182315.32
+ wint = 0
+ vth0 = -0.36907143
+ wkt1 = -4.5278925e-8
+ wkt2 = 7.5037926e-9
+ wtvfbsdoff = 0
+ wmax = 5.374e-7
+ aigc = 0.006152944
+ wmin = 2.674e-7
+ lkvth0we = 3e-12
+ tnoia = 0
+ version = 4.5
+ tempmod = 0
+ peta0 = -4.0225789e-16
+ ltvfbsdoff = 0
+ petab = 2.3283989e-16
+ wketa = 1.3494424e-8
+ wua1 = -1.7234672e-15
+ wub1 = 2.1940634e-24
+ wuc1 = 5.6346661e-17
+ tpbsw = 0.0025
+ acnqsmod = 0
+ toxref = 3e-9
+ bigc = 0.0012521
+ aigbacc = 0.012071
+ cjswd = 4.8144e-11
+ cjsws = 4.8144e-11
+ wwlc = 0
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ rbodymod = 0
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigc = 0.15259
+ aigbinv = 0.009974
+ tvfbsdoff = 0.1
+ ptvfbsdoff = 0
+ ltvoff = -1.5678858e-10
+ scref = 1e-6
+ pigcd = 2.572
+ aigsd = 0.0063633987
+ wpdiblc2 = -6.1394667e-10
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ lku0we = 1.8e-11
+ lvoff = -1.7133213e-9
+ epsrox = 3.9
+ lvsat = -0.0045167251000000005
+ poxedge = 1
+ lvth0 = 1.3595196e-9
+ k2we = 5e-5
+ wvfbsdoff = 0
+ rdsmod = 0
+ lvfbsdoff = 0
+ delta = 0.018814
+ dsub = 0.5
+ dtox = 3.91e-10
+ laigc = 1.1545174e-11
+ igbmod = 1
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ binunit = 2
+ rnoia = 0
+ rnoib = 0
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ pbswgd = 0.8
+ wkvth0we = 0.0
+ pbswgs = 0.8
+ eta0 = 0.08799813
+ pketa = 1.5922924e-16
+ etab = -0.088479977
+ ngate = 1.7e+20
+ ngcon = 1
+ igcmod = 1
+ wpclm = -3.0982532e-8
+ trnqsmod = 0
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ paigsd = 2.0055591e-22
+ rgatemod = 0
+ tnjtsswg = 1
+ permod = 1
+ )

.model pch_sf_33 pmos (
+ level = 54
+ version = 4.5
+ pdits = 0
+ cigsd = 0.013281
+ tempmod = 0
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ tpbswg = 0.001
+ rshg = 14.1
+ aigbacc = 0.012071
+ wpdiblc2 = 3.3638075e-10
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ tnoia = 0
+ ptvoff = 0
+ aigbinv = 0.009974
+ peta0 = 1.6e-17
+ waigsd = 1.9846811e-12
+ wketa = -1.9384664e-9
+ tpbsw = 0.0025
+ tnom = 25
+ diomod = 1
+ cjswd = 4.8144e-11
+ cjsws = 4.8144e-11
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ wkvth0we = 0.0
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.7086399999999997e-10
+ pku0we = 0.0
+ cjswgs = 1.7086399999999997e-10
+ trnqsmod = 0
+ tvfbsdoff = 0.1
+ poxedge = 1
+ mjswgd = 0.95
+ wags = 5.1942014e-9
+ mjswgs = 0.95
+ tcjswg = 0.00128
+ binunit = 2
+ scref = 1e-6
+ voff = -0.10372023
+ acde = 0.5
+ pigcd = 2.572
+ aigsd = 0.0063632583
+ rgatemod = 0
+ vsat = 108525.44
+ tnjtsswg = 1
+ wint = 0
+ vth0 = -0.34887115999999996
+ lvoff = 0
+ wkt1 = -3.0503659e-9
+ wkt2 = -7.2833333e-10
+ wmax = 2.674e-7
+ aigc = 0.0068302204
+ wmin = 1.08e-7
+ lvsat = -8.000000000000001e-6
+ lvth0 = 2.4e-10
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ delta = 0.018814
+ wua1 = -5.5326541e-17
+ wub1 = -1.0689498e-25
+ wuc1 = -1.2119467e-17
+ fprout = 200
+ rnoia = 0
+ rnoib = 0
+ bigc = 0.0012521
+ wute = -7.6523556e-8
+ xrcrg1 = 12
+ xrcrg2 = 1
+ wwlc = 0
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ ngate = 1.7e+20
+ ngcon = 1
+ cdsc = 0
+ wpclm = 7.1298978e-9
+ cgbo = 0
+ cgdl = 3.0105e-11
+ wtvoff = -7.3630015e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigc = 0.15259
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ capmod = 2
+ wku0we = 1.5e-11
+ mobmod = 0
+ njtsswg = 6.489
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ k2we = 5e-5
+ ckappad = 0.6
+ ckappas = 0.6
+ ijthsfwd = 0.01
+ pdiblc1 = 0
+ pdiblc2 = 0.0015492917
+ dsub = 0.5
+ pdiblcb = 0
+ dtox = 3.91e-10
+ tvoff = 0.0025423547
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ eta0 = 0.10792519
+ etab = -0.13555556
+ ijthsrev = 0.01
+ ku0we = -0.0007
+ bigbacc = 0.0054401
+ beta0 = 13.32
+ leta0 = 4.8e-10
+ wtvfbsdoff = 0
+ kvth0we = -0.00022
+ ppclm = 0
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ dlcig = 2.5e-9
+ lintnoi = -5e-9
+ bgidl = 1834800000.0
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ ltvfbsdoff = 0
+ ppdiblc2 = 0
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ toxref = 3e-9
+ bigsd = 0.0003327
+ ptvfbsdoff = 0
+ pkvth0we = 0.0
+ wvoff = 1.4142431e-9
+ a0 = 2.5876667
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ at = 72000
+ cf = 8.17e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.015389268
+ k3 = -2.5823
+ em = 20000000.0
+ ll = 0
+ lw = 0
+ u0 = 0.0094871852
+ w0 = 0
+ ua = -1.9215717e-10
+ ub = 1.2747184e-18
+ uc = -1.7585185e-12
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ wvsat = -0.0013318206
+ nfactor = 1
+ wvth0 = -1.0654371999999995e-9
+ vfbsdoff = 0.01
+ waigc = 1.6569661e-12
+ keta = 0.02482765
+ ltvoff = 0
+ jswd = 3.69e-13
+ lketa = 0
+ jsws = 3.69e-13
+ paramchk = 1
+ lcit = -1.6e-11
+ xpart = 1
+ pvfbsdoff = 0
+ kt1l = 0
+ lku0we = 1.8e-11
+ nigbacc = 10
+ egidl = 0.001
+ epsrox = 3.9
+ lint = 6.5375218e-9
+ lkt1 = 4.8e-10
+ lmax = 2.001e-5
+ lmin = 8.9991e-6
+ rdsmod = 0
+ ijthdfwd = 0.01
+ lpe0 = 6.44e-8
+ igbmod = 1
+ lpeb = 0
+ nigbinv = 2.171
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ minv = -0.33
+ pbswgd = 0.8
+ pbswgs = 0.8
+ ndep = 1e+18
+ ags = 0.89683683
+ lwlc = 0
+ igcmod = 1
+ moin = 5.5538
+ ijthdrev = 0.01
+ cjd = 0.001270624
+ cit = 5e-6
+ cjs = 0.001270624
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 1.0572421799999999e-8
+ nigc = 2.291
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ lpdiblc2 = 0
+ fnoimod = 1
+ pvoff = -2e-17
+ eigbinv = 1.1
+ cdscb = 0
+ cdscd = 0
+ la0 = 0
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ jsd = 1.5e-7
+ pvsat = 0
+ jss = 1.5e-7
+ lat = -0.00064
+ kt1 = -0.17197747
+ lk2 = -3.2000000000000003e-10
+ kt2 = -0.050761111
+ wk2we = 0.0
+ pvth0 = 1.2e-16
+ llc = 0
+ lln = 1
+ lu0 = 8e-13
+ drout = 0.56
+ mjd = 0.335
+ mjs = 0.335
+ lub = 0
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 0
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ pk2 = 0
+ pu0 = 0
+ ntox = 1.0
+ voffl = 0
+ prt = 0
+ pub = 0
+ pcit = 8.000000000000001e-19
+ pud = 0
+ pclm = 1.101657
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 9.8162749e-10
+ ub1 = -3.8648101e-20
+ uc1 = 8.1681111e-11
+ tpb = 0.0016
+ weta0 = 2.3643289e-9
+ permod = 1
+ wa0 = 4.8944e-8
+ wetab = 2.9133333e-9
+ ute = -0.81574074
+ phin = 0.15
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 3.9065138e-9
+ lkvth0we = 3e-12
+ lpclm = 0
+ wlc = 0
+ wln = 1
+ wu0 = 5.8460889e-11
+ xgl = -8.2e-9
+ xgw = 0
+ wua = -4.8614483e-17
+ wub = 8.106039e-27
+ wuc = 3.3309111e-18
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ cigbacc = 0.245
+ pkt1 = 4e-17
+ cgidl = 1
+ tnoimod = 0
+ acnqsmod = 0
+ voffcv = -0.125
+ wpemod = 1
+ rbdb = 50
+ prwb = 0
+ prwg = 0
+ rbpb = 50
+ rbpd = 50
+ cigbinv = 0.006
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ pbswd = 0.9
+ rbodymod = 0
+ pbsws = 0.9
+ rdsw = 200
+ )

.model pch_sf_34 pmos (
+ level = 54
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ nfactor = 1
+ ptvoff = -5.393716e-17
+ k2we = 5e-5
+ waigsd = 1.9861139e-12
+ ijthdfwd = 0.01
+ dsub = 0.5
+ dtox = 3.91e-10
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ diomod = 1
+ bigsd = 0.0003327
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.7086399999999997e-10
+ pku0we = 0.0
+ cjswgs = 1.7086399999999997e-10
+ eta0 = 0.10792519
+ wvoff = 1.3100722e-9
+ etab = -0.13555556
+ ijthdrev = 0.01
+ nigbacc = 10
+ wvsat = -0.0013318206
+ wvth0 = -1.1611130999999997e-9
+ lpdiblc2 = 6.2970633e-9
+ waigc = 1.4905459e-12
+ mjswgd = 0.95
+ mjswgs = 0.95
+ tcjswg = 0.00128
+ nigbinv = 2.171
+ lketa = -5.5366519e-8
+ pvfbsdoff = 0
+ xpart = 1
+ egidl = 0.001
+ lkvth0we = 3e-12
+ fnoimod = 1
+ ags = 0.84380759
+ eigbinv = 1.1
+ fprout = 200
+ cjd = 0.001270624
+ cit = 5e-6
+ cjs = 0.001270624
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ acnqsmod = 0
+ dlc = 1.0572421799999999e-8
+ xrcrg1 = 12
+ xrcrg2 = 1
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ rbodymod = 0
+ la0 = -3.9401851e-7
+ wtvoff = -6.7630331e-11
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = -0.00064
+ kt1 = -0.17107141
+ kt2 = -0.050597496
+ lk2 = 5.211940300000001e-9
+ llc = 0
+ lln = 1
+ lu0 = 9.9758999e-10
+ mjd = 0.335
+ mjs = 0.335
+ lua = -7.2048384e-17
+ lub = 4.3514377e-25
+ luc = 1.4270275e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = -3.1655381e-14
+ pvoff = 9.1649624e-16
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ pk2 = 9.285497e-17
+ keta = 0.030986328
+ pu0 = 3.0504276e-17
+ prt = 0
+ cdscb = 0
+ cdscd = 0
+ pua = 2.7735079e-23
+ pub = -4.2717478e-32
+ puc = 1.20866e-25
+ pud = 0
+ cigbacc = 0.245
+ capmod = 2
+ pvsat = 0
+ rsh = 15.2
+ wk2we = 0.0
+ tcj = 0.000832
+ ua1 = 8.0734953e-10
+ pvth0 = 9.8012639e-16
+ ub1 = 2.6826436e-19
+ uc1 = 8.9789043e-11
+ drout = 0.56
+ lags = 4.7673289e-7
+ wku0we = 1.5e-11
+ tpb = 0.0016
+ wa0 = 5.2465177e-8
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ ute = -0.817454
+ paigc = 1.4961177e-18
+ lcit = -1.6e-11
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 3.8961851e-9
+ tnoimod = 0
+ mobmod = 0
+ wlc = 0
+ wln = 1
+ wu0 = 5.5067755e-11
+ xgl = -8.2e-9
+ xgw = 0
+ kt1l = 0
+ wua = -5.1699586e-17
+ wub = 1.2857705e-26
+ wuc = 3.3174666e-18
+ wud = 0
+ voffl = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ wpdiblc2 = 3.5925269e-10
+ cigbinv = 0.006
+ weta0 = 2.3643289e-9
+ wetab = 2.9133333e-9
+ lint = 6.5375218e-9
+ lpclm = 0
+ lkt1 = -7.6654893e-9
+ lkt2 = -1.4709041e-9
+ lmax = 8.9991e-6
+ lmin = 8.9908e-7
+ lpe0 = 6.44e-8
+ cgidl = 1
+ lpeb = 0
+ version = 4.5
+ tempmod = 0
+ minv = -0.33
+ wtvfbsdoff = 0
+ laigsd = -1.8524358e-14
+ lua1 = 1.5667589e-15
+ lub1 = -2.759143e-24
+ luc1 = -7.2890309e-17
+ ndep = 1e+18
+ wkvth0we = 0.0
+ lute = 1.5402209e-8
+ lwlc = 0
+ pbswd = 0.9
+ pbsws = 0.9
+ moin = 5.5538
+ aigbacc = 0.012071
+ ltvfbsdoff = 0
+ trnqsmod = 0
+ nigc = 2.291
+ pdits = 0
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ noff = 2.2684
+ cigsd = 0.013281
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ aigbinv = 0.009974
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ pags = -1.92428e-14
+ ntox = 1.0
+ pcit = 8.000000000000001e-19
+ rgatemod = 0
+ pclm = 1.101657
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ ptvfbsdoff = 0
+ tnjtsswg = 1
+ phin = 0.15
+ tnoia = 0
+ pkt1 = -2.7722214e-15
+ pkt2 = 2.4239149e-16
+ peta0 = 1.6e-17
+ toxref = 3e-9
+ wketa = -2.0595747e-9
+ poxedge = 1
+ tpbsw = 0.0025
+ cjswd = 4.8144e-11
+ cjsws = 4.8144e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ rbdb = 50
+ pua1 = -1.1776704e-22
+ binunit = 2
+ prwb = 0
+ pub1 = 2.7996299e-31
+ prwg = 0
+ puc1 = 9.811687e-24
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ pute = 1.5923616e-14
+ rdsw = 200
+ tvfbsdoff = 0.1
+ ltvoff = -3.3500511e-10
+ scref = 1e-6
+ pigcd = 2.572
+ rshg = 14.1
+ aigsd = 0.0063632604
+ lku0we = 1.8e-11
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ epsrox = 3.9
+ lvoff = -2.4480721e-8
+ a0 = 2.6314952
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ rdsmod = 0
+ wvfbsdoff = 0
+ at = 72000
+ cf = 8.17e-11
+ lvsat = -8.000000000000001e-6
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.016004612
+ k3 = -2.5823
+ em = 20000000.0
+ lvfbsdoff = 0
+ lvth0 = -1.3626904e-8
+ igbmod = 1
+ ll = 0
+ lw = 0
+ u0 = 0.0093763075
+ w0 = 0
+ ua = -1.8414289e-10
+ ub = 1.2263153e-18
+ uc = -3.3458683e-12
+ ud = 0
+ ijthsfwd = 0.01
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ delta = 0.018814
+ laigc = -5.3027874e-11
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ rnoia = 0
+ rnoib = 0
+ pbswgd = 0.8
+ pbswgs = 0.8
+ tnom = 25
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ igcmod = 1
+ pketa = 1.0887638e-15
+ ngate = 1.7e+20
+ ngcon = 1
+ ijthsrev = 0.01
+ wpclm = 7.1298978e-9
+ njtsswg = 6.489
+ gbmin = 1e-12
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ wags = 7.3346686e-9
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.00084883969
+ pdiblcb = 0
+ paigsd = -1.2880862e-20
+ voff = -0.10099712
+ acde = 0.5
+ ppdiblc2 = -2.0561872e-16
+ vsat = 108525.44
+ wint = 0
+ permod = 1
+ vth0 = -0.34732868
+ wkt1 = -2.7375492e-9
+ wkt2 = -7.5529568e-10
+ wmax = 2.674e-7
+ aigc = 0.0068361189
+ wmin = 1.08e-7
+ bigbacc = 0.0054401
+ tvoff = 0.0025796189
+ kvth0we = -0.00022
+ wua1 = -4.222676e-17
+ wub1 = -1.3803658e-25
+ wuc1 = -1.3210867e-17
+ xjbvd = 1
+ xjbvs = 1
+ voffcv = -0.125
+ wpemod = 1
+ lk2we = 0.0
+ lintnoi = -5e-9
+ bigc = 0.0012521
+ wute = -7.8294814e-8
+ bigbinv = 0.00149
+ pkvth0we = 0.0
+ wwlc = 0
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ cdsc = 0
+ ku0we = -0.0007
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ beta0 = 13.32
+ leta0 = 4.8e-10
+ vfbsdoff = 0.01
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigc = 0.15259
+ ppclm = 0
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ paramchk = 1
+ tpbswg = 0.001
+ )

.model pch_sf_35 pmos (
+ level = 54
+ cjsws = 4.8144e-11
+ cjswgd = 1.7086399999999997e-10
+ pku0we = 0.0
+ cjswgs = 1.7086399999999997e-10
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ ndep = 1e+18
+ lute = -1.0958354e-8
+ lwlc = 0
+ moin = 5.5538
+ ijthsrev = 0.01
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ tvfbsdoff = 0.1
+ nigc = 2.291
+ mjswgd = 0.95
+ mjswgs = 0.95
+ tcjswg = 0.00128
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ scref = 1e-6
+ pags = 1.1742809e-13
+ ppdiblc2 = -6.1367245e-16
+ pigcd = 2.572
+ ntox = 1.0
+ aigsd = 0.0063632396
+ pcit = 8.000000000000001e-19
+ pclm = 1.101657
+ lvoff = -2.4340257e-9
+ phin = 0.15
+ wvfbsdoff = 0
+ njtsswg = 6.489
+ lvfbsdoff = 0
+ lvsat = -8.000000000000001e-6
+ lvth0 = 2.1200595e-10
+ pkt1 = 5.7873331999999995e-15
+ pkt2 = -5.7270183e-16
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ delta = 0.018814
+ fprout = 200
+ laigc = -3.3884553e-11
+ xrcrg1 = 12
+ xrcrg2 = 1
+ ckappad = 0.6
+ ckappas = 0.6
+ rnoia = 0
+ rnoib = 0
+ pdiblc1 = 0
+ pdiblc2 = 0.0027845581
+ pdiblcb = 0
+ pkvth0we = 0.0
+ rbdb = 50
+ pua1 = -9.8048843e-24
+ prwb = 0
+ pub1 = -2.3189739e-32
+ prwg = 0
+ puc1 = -4.5795492e-24
+ pketa = -3.0075994e-15
+ rbpb = 50
+ rbpd = 50
+ ngate = 1.7e+20
+ rbps = 50
+ rbsb = 50
+ wtvoff = -2.2790108e-10
+ pvag = 2.1
+ pute = -9.4649237e-15
+ ngcon = 1
+ wpclm = 7.1298978e-9
+ rdsw = 200
+ vfbsdoff = 0.01
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ bigbacc = 0.0054401
+ capmod = 2
+ wku0we = 1.5e-11
+ kvth0we = -0.00022
+ mobmod = 0
+ paramchk = 1
+ lintnoi = -5e-9
+ rshg = 14.1
+ bigbinv = 0.00149
+ wtvfbsdoff = 0
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ ltvfbsdoff = 0
+ ijthdfwd = 0.01
+ tvoff = 0.0027416725
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ tnom = 25
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ ijthdrev = 0.01
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = 4.8e-10
+ lpdiblc2 = 4.574275e-9
+ ptvfbsdoff = 0
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ nfactor = 1
+ ppclm = 0
+ wags = -1.4622812e-7
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ voff = -0.12576869
+ acde = 0.5
+ vsat = 108525.44
+ wint = 0
+ vth0 = -0.36287801999999997
+ wkt1 = -1.2355026e-8
+ wkt2 = 1.605395e-10
+ dmcgt = 0
+ wmax = 2.674e-7
+ tcjsw = 9.34e-5
+ lkvth0we = 3e-12
+ aigc = 0.0068146096
+ wmin = 1.08e-7
+ nigbacc = 10
+ toxref = 3e-9
+ wua1 = -1.6353255e-16
+ wub1 = 2.0258446e-25
+ wuc1 = 2.9590615e-18
+ acnqsmod = 0
+ bigsd = 0.0003327
+ bigc = 0.0012521
+ wute = -4.9768365e-8
+ nigbinv = 2.171
+ wwlc = 0
+ wvoff = 3.4766421e-9
+ rbodymod = 0
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ wvsat = -0.0013318206
+ xtid = 3
+ xtis = 3
+ wvth0 = -3.9165319999999977e-10
+ ltvoff = -4.7923289e-10
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigc = 0.15259
+ waigc = 2.7104678e-12
+ fnoimod = 1
+ eigbinv = 1.1
+ pvfbsdoff = 0
+ lketa = 4.197898e-9
+ xpart = 1
+ lku0we = 1.8e-11
+ epsrox = 3.9
+ wpdiblc2 = 8.1773971e-10
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ ags = 1.7348065
+ dmdg = 0
+ egidl = 0.001
+ cjd = 0.001270624
+ rdsmod = 0
+ cit = -8.7888889e-5
+ cjs = 0.001270624
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 1.0572421799999999e-8
+ igbmod = 1
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ k2we = 5e-5
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ dsub = 0.5
+ dtox = 3.91e-10
+ pbswgd = 0.8
+ la0 = -1.044589e-6
+ cigbacc = 0.245
+ pbswgs = 0.8
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = -0.00064
+ kt1 = -0.11040563
+ kt2 = -0.048714998
+ lk2 = 2.7690726e-9
+ llc = 0
+ lln = 1
+ lu0 = -1.8164817999999999e-9
+ mjd = 0.335
+ mjs = 0.335
+ lua = -6.2776752e-16
+ lub = 4.4518935e-25
+ luc = 5.1177769e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ igcmod = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 1.0817056e-13
+ wkvth0we = 0.0
+ nsd = 1e+20
+ pbd = 0.75
+ tnoimod = 0
+ pat = 0
+ pbs = 0.75
+ pk2 = -1.5480351e-16
+ eta0 = 0.10792519
+ etab = -0.13555556
+ pu0 = 1.5955157e-16
+ prt = 0
+ pua = 4.4574845e-23
+ pub = -2.7161351e-32
+ puc = -4.8372521e-24
+ pud = 0
+ rsh = 15.2
+ trnqsmod = 0
+ tcj = 0.000832
+ ua1 = 2.771768e-9
+ ub1 = -3.1924567e-18
+ uc1 = -6.2120134e-12
+ cigbinv = 0.006
+ tpb = 0.0016
+ wa0 = -1.0464262e-7
+ ute = -0.78783539
+ pvoff = -1.01175093e-15
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 4.174453e-9
+ wlc = 0
+ wln = 1
+ wu0 = -8.9929205e-11
+ xgl = -8.2e-9
+ xgw = 0
+ wua = -7.0620672e-17
+ wub = -4.621089e-27
+ wuc = 8.8883858e-18
+ wud = 0
+ cdscb = 0
+ cdscd = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ pvsat = 0
+ a0 = 3.3624733
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ wk2we = 0.0
+ pvth0 = 2.9530712e-16
+ at = 72000
+ cf = 8.17e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.013259817
+ k3 = -2.5823
+ em = 20000000.0
+ drout = 0.56
+ version = 4.5
+ ll = 0
+ lw = 0
+ u0 = 0.012538186
+ w0 = 0
+ ua = 4.4026063e-10
+ ub = 1.2150282e-18
+ uc = -4.4814963e-11
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ paigc = 4.1038726e-19
+ xw = 8.600000000000001e-9
+ tempmod = 0
+ voffl = 0
+ rgatemod = 0
+ permod = 1
+ tnjtsswg = 1
+ weta0 = 2.3643289e-9
+ wetab = 2.9133333e-9
+ aigbacc = 0.012071
+ lpclm = 0
+ cgidl = 1
+ voffcv = -0.125
+ wpemod = 1
+ aigbinv = 0.009974
+ pbswd = 0.9
+ pbsws = 0.9
+ keta = -0.035939983
+ pdits = 0
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ lags = -3.1625612e-7
+ tpbswg = 0.001
+ poxedge = 1
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 6.6671111e-11
+ kt1l = 0
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ binunit = 2
+ lint = 6.5375218e-9
+ ptvoff = 8.8703803e-17
+ lkt1 = -6.1658035e-8
+ lkt2 = -3.1463267e-9
+ tnoia = 0
+ lmax = 8.9908e-7
+ waigsd = 1.9716411e-12
+ lmin = 4.4908e-7
+ ijthsfwd = 0.01
+ peta0 = 1.6e-17
+ lpe0 = 6.44e-8
+ lpeb = 0
+ wketa = 2.5430806e-9
+ diomod = 1
+ tpbsw = 0.0025
+ minv = -0.33
+ lua1 = -1.8157361e-16
+ lub1 = 3.2089876e-25
+ luc1 = 1.2550631e-17
+ pditsd = 0
+ cjswd = 4.8144e-11
+ pditsl = 0
+ )

.model pch_sf_36 pmos (
+ level = 54
+ ags = 0.79842724
+ pvfbsdoff = 0
+ wcit = 5.8162887e-11
+ lketa = -1.0850486e-8
+ cigbacc = 0.245
+ cjd = 0.001270624
+ cit = -0.00049977211
+ cjs = 0.001270624
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ voff = -0.11894985
+ xpart = 1
+ dlc = 1.38228675e-8
+ k3b = 2.1176
+ acde = 0.5
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ rgatemod = 0
+ tnjtsswg = 1
+ vsat = 108525.44
+ tnoimod = 0
+ wint = 0
+ vth0 = -0.36950626
+ egidl = 0.001
+ wkt1 = 8.365112e-10
+ wkt2 = -1.4765978e-9
+ la0 = -3.2362015e-7
+ wmax = 2.674e-7
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = -0.00064
+ aigc = 0.0068096243
+ wmin = 1.08e-7
+ kt1 = -0.25321364
+ kt2 = -0.04359324
+ lk2 = -6.627309e-10
+ llc = -1.18e-13
+ lln = 0.7
+ cigbinv = 0.006
+ lu0 = -4.4979608e-10
+ mjd = 0.335
+ mjs = 0.335
+ lua = -1.7021816e-16
+ lub = 1.0550853e-25
+ luc = -1.2975077e-17
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ fprout = 200
+ njs = 1.02
+ pa0 = -3.1370244e-14
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 0
+ pbs = 0.75
+ pk2 = 1.4083403e-16
+ xrcrg1 = 12
+ xrcrg2 = 1
+ pu0 = -1.3937081e-17
+ prt = 0
+ pua = 4.7117679e-24
+ pub = -8.7289665e-33
+ puc = -3.0945045e-25
+ pud = 0
+ wua1 = -2.3000717e-16
+ wub1 = 1.2114667e-25
+ wuc1 = -1.9684753e-17
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 2.6350858e-9
+ ub1 = -2.2549964e-18
+ uc1 = 3.1191962e-11
+ bigc = 0.0012521
+ wute = -1.1762912e-7
+ version = 4.5
+ tpb = 0.0016
+ wa0 = 2.1249557e-7
+ wwlc = 0
+ ute = -0.71022675
+ wtvoff = -1.1036076e-10
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 3.5025496e-9
+ tempmod = 0
+ wlc = 0
+ wln = 1
+ wu0 = 3.0436319e-10
+ xgl = -8.2e-9
+ xgw = 0
+ wua = 1.9977231e-17
+ wub = -4.6512873e-26
+ wuc = -1.4020724e-18
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ wtvfbsdoff = 0
+ aigbacc = 0.012071
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigc = 0.15259
+ pvoff = 7.5942711e-17
+ capmod = 2
+ cdscb = 0
+ cdscd = 0
+ wku0we = 1.5e-11
+ pvsat = 0
+ wk2we = 0.0
+ pvth0 = -1.1393785e-16
+ ltvfbsdoff = 0
+ drout = 0.56
+ mobmod = 0
+ paigc = -1.759214e-19
+ aigbinv = 0.009974
+ voffl = 0
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ weta0 = 2.3643289e-9
+ wetab = 2.9133333e-9
+ lpclm = 0
+ k2we = 5e-5
+ ijthsfwd = 0.01
+ cgidl = 1
+ dsub = 0.5
+ ptvfbsdoff = 0
+ dtox = 3.91e-10
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ poxedge = 1
+ eta0 = 0.10792519
+ pbswd = 0.9
+ etab = -0.13555556
+ pbsws = 0.9
+ ijthsrev = 0.01
+ binunit = 2
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ pdits = 0
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ ppdiblc2 = 9.2177422e-17
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ tnoia = 0
+ toxref = 3e-9
+ peta0 = 1.6e-17
+ wketa = -1.9938172e-9
+ tpbsw = 0.0025
+ cjswd = 4.8144e-11
+ cjsws = 4.8144e-11
+ pkvth0we = 0.0
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ tvfbsdoff = 0.1
+ ltvoff = -1.9203223e-10
+ vfbsdoff = 0.01
+ njtsswg = 6.489
+ keta = -0.0017391106
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ lags = 9.5750741e-8
+ lku0we = 1.8e-11
+ paramchk = 1
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ scref = 1e-6
+ ckappad = 0.6
+ ckappas = 0.6
+ lcit = 2.4789973e-10
+ pdiblc1 = 0
+ pdiblc2 = 0.016049816
+ epsrox = 3.9
+ pdiblcb = 0
+ pigcd = 2.572
+ kt1l = 0
+ aigsd = 0.0063632396
+ rdsmod = 0
+ lvoff = -5.4343156e-9
+ wvfbsdoff = 0
+ lint = 9.7879675e-9
+ igbmod = 1
+ lvfbsdoff = 0
+ lkt1 = 1.177866e-9
+ lkt2 = -5.3999005e-9
+ lvsat = -8.000000000000001e-6
+ lmax = 4.4908e-7
+ lvth0 = 3.1284329e-9
+ lmin = 2.1577e-7
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ ijthdfwd = 0.01
+ lpe0 = 6.44e-8
+ delta = 0.018814
+ bigbacc = 0.0054401
+ lpeb = 0
+ pbswgd = 0.8
+ laigc = -3.1691048e-11
+ pbswgs = 0.8
+ rnoia = 0
+ rnoib = 0
+ minv = -0.33
+ igcmod = 1
+ lua1 = -1.2143343e-16
+ lub1 = -9.158653e-26
+ luc1 = -3.907118e-18
+ kvth0we = -0.00022
+ ndep = 1e+18
+ lute = -4.5106156e-8
+ pketa = -1.0113644e-15
+ ngate = 1.7e+20
+ lwlc = 0
+ lintnoi = -5e-9
+ moin = 5.5538
+ ijthdrev = 0.01
+ ngcon = 1
+ bigbinv = 0.00149
+ wpclm = 7.1298978e-9
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ nigc = 2.291
+ lpdiblc2 = -1.262443e-9
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ pags = 5.2660461e-14
+ permod = 1
+ ntox = 1.0
+ pcit = -2.4791670000000003e-17
+ pclm = 1.101657
+ phin = 0.15
+ lkvth0we = 3e-12
+ pkt1 = -1.70475e-17
+ pkt2 = 1.4763857e-16
+ voffcv = -0.125
+ wpemod = 1
+ tvoff = 0.0020889601
+ nfactor = 1
+ xjbvd = 1
+ acnqsmod = 0
+ xjbvs = 1
+ lk2we = 0.0
+ a0 = 1.7239078
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ rbdb = 50
+ pua1 = 1.9443948e-23
+ prwb = 0
+ pub1 = 1.2643651e-32
+ prwg = 0
+ at = 72000
+ puc1 = 5.3837292e-24
+ cf = 8.17e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.0054602636
+ k3 = -2.5823
+ em = 20000000.0
+ rbpb = 50
+ rbpd = 50
+ ll = -1.18e-13
+ lw = 0
+ rbps = 50
+ u0 = 0.009432082
+ rbsb = 50
+ pvag = 2.1
+ w0 = 0
+ rbodymod = 0
+ ua = -5.9962427e-10
+ ub = 1.98703e-18
+ uc = 1.0098696e-10
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ pute = 2.0393808e-14
+ xw = 8.600000000000001e-9
+ rdsw = 200
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = 4.8e-10
+ nigbacc = 10
+ ppclm = 0
+ tpbswg = 0.001
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ rshg = 14.1
+ nigbinv = 2.171
+ wpdiblc2 = -7.8646151e-10
+ ptvoff = 3.6984079e-17
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ waigsd = 1.9716411e-12
+ diomod = 1
+ fnoimod = 1
+ pditsd = 0
+ pditsl = 0
+ bigsd = 0.0003327
+ cjswgd = 1.7086399999999997e-10
+ pku0we = 0.0
+ tnom = 25
+ cjswgs = 1.7086399999999997e-10
+ eigbinv = 1.1
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ wkvth0we = 0.0
+ wvoff = 1.0046111e-9
+ trnqsmod = 0
+ wvsat = -0.0013318206
+ mjswgd = 0.95
+ wvth0 = 5.384490000000004e-10
+ mjswgs = 0.95
+ tcjswg = 0.00128
+ waigc = 4.0429874e-12
+ wags = 9.7102189e-10
+ )

.model pch_sf_37 pmos (
+ level = 54
+ fprout = 200
+ lvth0 = 5.7674905e-9
+ xrcrg1 = 12
+ xrcrg2 = 1
+ delta = 0.018814
+ wtvfbsdoff = 0
+ laigc = -4.357169e-12
+ rnoia = 0
+ rnoib = 0
+ acnqsmod = 0
+ wtvoff = 1.2048366e-10
+ ltvfbsdoff = 0
+ pketa = 4.1278959e-16
+ ngate = 1.7e+20
+ rbodymod = 0
+ ngcon = 1
+ wpclm = 6.8691006e-8
+ capmod = 2
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ wku0we = 1.5e-11
+ keta = -0.058692164
+ mobmod = 0
+ nfactor = 1
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 9.291477e-12
+ ptvfbsdoff = 0
+ kt1l = 0
+ wpdiblc2 = -7.28246e-10
+ lint = 9.7879675e-9
+ lkt1 = -4.1970694e-9
+ lkt2 = -3.7791597e-9
+ lmax = 2.1577e-7
+ lmin = 9e-8
+ lpe0 = 6.44e-8
+ nigbacc = 10
+ lpeb = 0
+ tvoff = 0.0011827459
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ minv = -0.33
+ lua1 = -2.1218464e-16
+ lub1 = 2.7818737e-25
+ luc1 = 2.2554944e-17
+ ndep = 1e+18
+ wkvth0we = 0.0
+ lute = 1.5508066e-9
+ lwlc = 0
+ moin = 5.5538
+ nigbinv = 2.171
+ ku0we = -0.0007
+ trnqsmod = 0
+ beta0 = 13.32
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ nigc = 2.291
+ leta0 = 4.8e-10
+ ppclm = -1.2989269e-14
+ noff = 2.2684
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ fnoimod = 1
+ eigbinv = 1.1
+ ntox = 1.0
+ rgatemod = 0
+ pcit = 1.2014196000000001e-17
+ pclm = 0.85425247
+ tnjtsswg = 1
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ phin = 0.15
+ toxref = 3e-9
+ pkt1 = -1.917336e-16
+ pkt2 = 3.7767926e-16
+ bigsd = 0.0003327
+ cigbacc = 0.245
+ rbdb = 50
+ pua1 = 2.6827919e-23
+ prwb = 0
+ pub1 = -3.4278711e-32
+ prwg = 0
+ puc1 = -2.7535024e-24
+ wvoff = 8.5374562e-10
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ pute = -4.2802262e-16
+ ltvoff = -8.1627e-13
+ rdsw = 200
+ tnoimod = 0
+ wvsat = -0.00089129698
+ ags = 1.2522222
+ wvth0 = -4.909479999999996e-10
+ cjd = 0.001270624
+ cit = 0.00063107268
+ cjs = 0.001270624
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 1.38228675e-8
+ waigc = 1.4660694e-11
+ k3b = 2.1176
+ cigbinv = 0.006
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ pvfbsdoff = 0
+ lku0we = 1.8e-11
+ lketa = 1.1666086e-9
+ epsrox = 3.9
+ la0 = 6.219346e-9
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = -0.0081843287
+ xpart = 1
+ kt1 = -0.22773883
+ kt2 = -0.051274476
+ lk2 = 3.3511471e-9
+ llc = -1.18e-13
+ lln = 0.7
+ lu0 = -1.6234862e-10
+ mjd = 0.335
+ version = 4.5
+ mjs = 0.335
+ lua = 1.3101868e-17
+ lub = -8.7271368e-26
+ luc = -1.2812174e-17
+ lud = 0
+ rshg = 14.1
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = -2.0637395e-14
+ rdsmod = 0
+ nsd = 1e+20
+ pbd = 0.75
+ tempmod = 0
+ pat = -5.0045721e-10
+ pbs = 0.75
+ pk2 = 4.0368065e-17
+ egidl = 0.001
+ igbmod = 1
+ pu0 = -5.2679707e-18
+ prt = 0
+ pua = -4.0286539e-24
+ pub = 7.5106005e-33
+ puc = 1.4358513e-24
+ pud = 0
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 3.0651863e-9
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ ub1 = -4.0074881e-18
+ uc1 = -9.4220652e-11
+ tpb = 0.0016
+ aigbacc = 0.012071
+ wa0 = 1.6162969e-7
+ pbswgd = 0.8
+ pbswgs = 0.8
+ ute = -0.93134979
+ ijthsfwd = 0.01
+ wat = 0.0023718351
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 3.9786916e-9
+ wlc = 0
+ wln = 1
+ wu0 = 2.6327735e-10
+ xgl = -8.2e-9
+ xgw = 0
+ wua = 6.1401032e-17
+ wub = -1.2347765e-25
+ wuc = -9.6736445e-18
+ wud = 0
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ igcmod = 1
+ tnom = 25
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ aigbinv = 0.009974
+ ijthsrev = 0.01
+ pvoff = 1.0777532e-16
+ cdscb = 0
+ cdscd = 0
+ pvsat = -9.2948987e-11
+ wags = 2.5054667e-7
+ wk2we = 0.0
+ pvth0 = 1.03264908e-16
+ drout = 0.56
+ wcit = -1.162725e-10
+ paigc = -2.4162575e-18
+ permod = 1
+ voff = -0.1339517
+ acde = 0.5
+ ppdiblc2 = 7.9894307e-17
+ voffl = 0
+ poxedge = 1
+ vsat = 106518.57
+ wint = 0
+ vth0 = -0.38201365
+ weta0 = 2.3643289e-9
+ wetab = 2.9133333e-9
+ wkt1 = 1.664079e-9
+ wkt2 = -2.566838e-9
+ wmax = 2.674e-7
+ lpclm = 5.2201277e-8
+ binunit = 2
+ aigc = 0.0066800799
+ wmin = 1.08e-7
+ voffcv = -0.125
+ wpemod = 1
+ cgidl = 1
+ wua1 = -2.6500229e-16
+ wub1 = 3.4352994e-25
+ wuc1 = 1.8880326e-17
+ bigc = 0.0012521
+ wute = -1.8947457e-8
+ pkvth0we = 0.0
+ wwlc = 0
+ pbswd = 0.9
+ pbsws = 0.9
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ vfbsdoff = 0.01
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigc = 0.15259
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ pdits = 0
+ tpbswg = 0.001
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ paramchk = 1
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ ptvoff = -1.1725409e-17
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ a0 = 0.16068118
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ waigsd = 1.9716411e-12
+ at = 107755.11
+ cf = 8.17e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.024483382
+ k3 = -2.5823
+ em = 20000000.0
+ ll = -1.18e-13
+ lw = 0
+ u0 = 0.0080697718
+ tnoia = 0
+ w0 = 0
+ ua = -1.4684396e-9
+ ub = 2.9006788e-18
+ uc = 1.0021491e-10
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ diomod = 1
+ k2we = 5e-5
+ ijthdfwd = 0.01
+ peta0 = 1.6e-17
+ njtsswg = 6.489
+ dsub = 0.5
+ dtox = 3.91e-10
+ wketa = -8.743362e-9
+ pditsd = 0
+ pditsl = 0
+ cjswgd = 1.7086399999999997e-10
+ pku0we = 0.0
+ cjswgs = 1.7086399999999997e-10
+ tpbsw = 0.0025
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ cjswd = 4.8144e-11
+ cjsws = 4.8144e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ ckappad = 0.6
+ ckappas = 0.6
+ pdiblc1 = 0
+ pdiblc2 = 0.01690182
+ eta0 = 0.10792519
+ pdiblcb = 0
+ etab = -0.13555556
+ tvfbsdoff = 0.1
+ ijthdrev = 0.01
+ mjswgd = 0.95
+ mjswgs = 0.95
+ lpdiblc2 = -1.4422174e-9
+ tcjswg = 0.00128
+ bigbacc = 0.0054401
+ scref = 1e-6
+ pigcd = 2.572
+ aigsd = 0.0063632396
+ kvth0we = -0.00022
+ wvfbsdoff = 0
+ lvoff = -2.268926e-9
+ lintnoi = -5e-9
+ lvfbsdoff = 0
+ bigbinv = 0.00149
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ lkvth0we = 3e-12
+ lvsat = 0.00041543719
+ )

.model pch_sf_38 pmos (
+ level = 54
+ poxedge = 1
+ ptvfbsdoff = 0
+ rdsw = 200
+ capmod = 2
+ vfbsdoff = 0.01
+ wku0we = 1.5e-11
+ pvoff = -1.6373467e-16
+ binunit = 2
+ cdscb = 0
+ cdscd = 0
+ mobmod = 0
+ pvsat = 1.729604e-10
+ wk2we = 0.0
+ pvth0 = 1.76763134e-16
+ drout = 0.56
+ paramchk = 1
+ paigc = -1.1563004e-18
+ voffl = 0
+ rshg = 14.1
+ weta0 = 1.3181501e-8
+ wetab = 4.1458967e-9
+ lpclm = -1.0127779e-7
+ ijthdfwd = 0.01
+ jtsswgd = 1.75e-7
+ cgidl = 1
+ jtsswgs = 1.75e-7
+ tnom = 25
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ pbswd = 0.9
+ pbsws = 0.9
+ ijthdrev = 0.01
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ lpdiblc2 = -1.4113545e-11
+ pdits = 0
+ cigsd = 0.013281
+ wags = 2.5054667e-7
+ dvt0w = 0
+ dvt1w = 0
+ njtsswg = 6.489
+ dvt2w = 0
+ wcit = 7.0487744e-11
+ xtsswgd = 0.32
+ voff = -0.14478455
+ xtsswgs = 0.32
+ acde = 0.5
+ pk2we = 0.0
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ ckappad = 0.6
+ ckappas = 0.6
+ vsat = 137363.5
+ wint = 0
+ pdiblc1 = 0
+ pdiblc2 = 0.0017092259
+ vth0 = -0.31880653
+ pdiblcb = 0
+ wkt1 = -1.350742e-8
+ wkt2 = 1.8825744e-9
+ toxref = 3e-9
+ wmax = 2.674e-7
+ lkvth0we = 3e-12
+ aigc = 0.0067219883
+ wmin = 1.08e-7
+ tnoia = 0
+ peta0 = -1.0008142e-15
+ petab = -1.1586096e-16
+ wketa = -6.6698086e-9
+ wua1 = 1.6631395e-16
+ wub1 = -2.121384e-25
+ wuc1 = 2.5860689e-17
+ tpbsw = 0.0025
+ acnqsmod = 0
+ bigbacc = 0.0054401
+ cjswd = 4.8144e-11
+ bigc = 0.0012521
+ cjsws = 4.8144e-11
+ wute = -6.1363432e-8
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ wwlc = 0
+ tvfbsdoff = 0.1
+ ltvoff = 3.7319947e-11
+ rbodymod = 0
+ kvth0we = -0.00022
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ xtid = 3
+ xtis = 3
+ lintnoi = -5e-9
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ bigbinv = 0.00149
+ cigc = 0.15259
+ vtsswgd = 1.1
+ vtsswgs = 1.1
+ lku0we = 1.8e-11
+ epsrox = 3.9
+ scref = 1e-6
+ pigcd = 2.572
+ aigsd = 0.0063632396
+ rdsmod = 0
+ wpdiblc2 = 8.0253658e-11
+ igbmod = 1
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ lvoff = -1.2506377e-9
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ lvsat = -0.0024839865000000003
+ pbswgd = 0.8
+ pbswgs = 0.8
+ lvth0 = -1.739787e-10
+ k2we = 5e-5
+ delta = 0.018814
+ laigc = -8.2965642e-12
+ dsub = 0.5
+ igcmod = 1
+ dtox = 3.91e-10
+ rnoia = 0
+ rnoib = 0
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ nfactor = 1
+ wkvth0we = 0.0
+ pketa = 2.1787556e-16
+ ngate = 1.7e+20
+ eta0 = 0.024468866
+ etab = -0.22797789
+ ngcon = 1
+ wpclm = -1.6917696e-7
+ trnqsmod = 0
+ gbmin = 1e-12
+ jswgd = 3.69e-13
+ jswgs = 3.69e-13
+ nigbacc = 10
+ permod = 1
+ rgatemod = 0
+ tnjtsswg = 1
+ nigbinv = 2.171
+ voffcv = -0.125
+ wpemod = 1
+ tvoff = 0.00077704148
+ xjbvd = 1
+ xjbvs = 1
+ lk2we = 0.0
+ fnoimod = 1
+ eigbinv = 1.1
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = 8.324894e-9
+ letab = 8.6876992e-9
+ tpbswg = 0.001
+ ppclm = 9.3703198e-15
+ keta = -0.049241031
+ dlcig = 2.5e-9
+ bgidl = 1834800000.0
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 1.1130569000000001e-10
+ kt1l = 0
+ ptvoff = 1.952106e-17
+ cigbacc = 0.245
+ waigsd = 1.9716411e-12
+ dmcgt = 0
+ lint = 0
+ tcjsw = 9.34e-5
+ tnoimod = 0
+ lkt1 = -6.1146074e-9
+ lkt2 = 9.2375447e-10
+ diomod = 1
+ lmax = 9e-8
+ lmin = 5.4e-8
+ ijthsfwd = 0.01
+ lpe0 = 6.44e-8
+ pditsd = 0
+ pditsl = 0
+ lpeb = 0
+ cigbinv = 0.006
+ cjswgd = 1.7086399999999997e-10
+ pku0we = 0.0
+ cjswgs = 1.7086399999999997e-10
+ bigsd = 0.0003327
+ minv = -0.33
+ ags = 1.2522222
+ lua1 = 1.5814311e-16
+ lub1 = -2.3663254e-25
+ luc1 = 3.1466117e-17
+ cjd = 0.001270624
+ cit = -0.00045418481
+ cjs = 0.001270624
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ ndep = 1e+18
+ bvs = 8.2
+ lute = -1.2895214e-8
+ dlc = 4.0349e-9
+ wvoff = 3.7421498e-9
+ k3b = 2.1176
+ lwlc = 0
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ version = 4.5
+ moin = 5.5538
+ mjswgd = 0.95
+ mjswgs = 0.95
+ ijthsrev = 0.01
+ tempmod = 0
+ wvsat = -0.0037201203
+ nigc = 2.291
+ tcjswg = 0.00128
+ wvth0 = -1.2728439999999995e-9
+ la0 = 3.4503642e-8
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = -0.0086928059
+ kt1 = -0.20733948
+ kt2 = -0.10130548
+ lk2 = 5.227863e-9
+ waigc = 1.256895e-12
+ llc = 0
+ lln = 1
+ a0 = -0.1402156
+ a1 = 0
+ a2 = 1
+ b0 = 0
+ b1 = 0
+ lu0 = 4.660914e-11
+ mjd = 0.335
+ mjs = 0.335
+ lua = 1.1003971e-16
+ lub = -1.3258131e-25
+ luc = -1.072064e-17
+ at = 113164.44
+ lud = 0
+ cf = 8.17e-11
+ lwc = 0
+ pvfbsdoff = 0
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.044448444
+ k3 = -2.5823
+ lwl = 0
+ lwn = 1
+ em = 20000000.0
+ aigbacc = 0.012071
+ njd = 1.02
+ njs = 1.02
+ ll = 0
+ noff = 2.2684
+ pa0 = -6.959911e-15
+ lw = 0
+ u0 = 0.0058468169
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ w0 = 0
+ nsd = 1e+20
+ pbd = 0.75
+ pat = 1.1859675e-9
+ ua = -2.4996932e-9
+ ub = 3.3826995e-18
+ uc = 7.7964547e-11
+ ud = 0
+ pbs = 0.75
+ pk2 = -8.547569e-17
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ pu0 = 1.7354187e-18
+ prt = 0
+ lketa = 2.7820203e-10
+ pua = -5.4706466e-24
+ pub = 7.2761107e-33
+ puc = 2.7207836e-25
+ pud = 0
+ wtvfbsdoff = 0
+ xpart = 1
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = -8.7447052e-10
+ ub1 = 1.4693195e-18
+ uc1 = -1.8902037e-10
+ ppdiblc2 = 3.8953385e-18
+ ntox = 1.0
+ tpb = 0.0016
+ pcit = -5.5412666999999994e-18
+ pclm = 2.4870084
+ wa0 = 1.612455e-8
+ ute = -0.77766872
+ wat = -0.015568853
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 5.3174549e-9
+ aigbinv = 0.009974
+ wlc = 0
+ egidl = 0.001
+ wln = 1
+ wu0 = 1.8877321e-10
+ xgl = -8.2e-9
+ xgw = 0
+ wua = 7.6741379e-17
+ wub = -1.2098307e-25
+ wuc = 2.7069183e-18
+ wud = 0
+ wwc = 0
+ ltvfbsdoff = 0
+ wwl = 0
+ wwn = 1
+ phin = 0.15
+ fprout = 200
+ xrcrg1 = 12
+ xrcrg2 = 1
+ pkt1 = 1.2343873e-15
+ pkt2 = -4.056551e-17
+ wtvoff = -2.1192558e-10
+ pkvth0we = 0.0
+ rbdb = 50
+ pua1 = -1.3715808e-23
+ prwb = 0
+ pub1 = 1.7954113e-32
+ prwg = 0
+ puc1 = -3.4096566e-24
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbsb = 50
+ pvag = 2.1
+ pute = 3.5590791e-15
+ )

.model pch_sf_39 pmos (
+ level = 54
+ fnoimod = 1
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ eigbinv = 1.1
+ k2we = 5e-5
+ ijthsfwd = 0.01
+ tvoff = 0.00092289205
+ dsub = 0.5
+ dtox = 3.91e-10
+ xjbvd = 1
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ xjbvs = 1
+ lk2we = 0.0
+ eta0 = 0.19463541
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ etab = -0.16706384
+ ijthsrev = 0.01
+ cigbacc = 0.245
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = -1.5447657000000001e-9
+ letab = 5.1546845e-9
+ tnoimod = 0
+ ppclm = 7.8094068e-15
+ dlcig = 2.5e-9
+ cigbinv = 0.006
+ bgidl = 1834800000.0
+ ppdiblc2 = 0
+ toxref = 3e-9
+ version = 4.5
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ tempmod = 0
+ ags = 1.2522222
+ cjd = 0.001270624
+ cit = -0.0026753087
+ cjs = 0.001270624
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 4.0349e-9
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ aigbacc = 0.012071
+ bigsd = 0.0003327
+ pkvth0we = 0.0
+ la0 = -1.4904033e-7
+ ltvoff = 2.8860613e-11
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0.008732509
+ kt1 = -0.53950997
+ kt2 = -0.12590838
+ lk2 = 3.8965993000000006e-9
+ wvoff = 1.4341134e-10
+ llc = 0
+ lln = 1
+ lu0 = 4.1731088999999996e-10
+ mjd = 0.335
+ mjs = 0.335
+ lua = 7.9060667e-17
+ lub = -2.7964918e-26
+ luc = 5.5424848e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = -2.574678e-15
+ nsd = 1e+20
+ pbd = 0.75
+ pat = -1.0212358e-9
+ wvsat = -0.0027183681
+ pbs = 0.75
+ pk2 = 2.1304022e-16
+ aigbinv = 0.009974
+ wvth0 = -2.2127999999999575e-11
+ pu0 = -6.6237547e-17
+ vfbsdoff = 0.01
+ prt = 0
+ pua = -2.0419953e-23
+ pub = 1.469069e-32
+ puc = 1.2609666e-24
+ pud = 0
+ waigc = 6.0357037e-12
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 8.3453493e-9
+ ub1 = -1.1410668e-17
+ pvfbsdoff = 0
+ uc1 = 1.6197295e-9
+ keta = -0.31465021
+ lku0we = 1.8e-11
+ tpb = 0.0016
+ wa0 = -5.9482929e-8
+ epsrox = 3.9
+ ute = -1
+ wat = 0.022486376
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 1.7062889e-10
+ wlc = 0
+ wln = 1
+ wu0 = 1.3607209e-9
+ xgl = -8.2e-9
+ xgw = 0
+ wua = 3.3448805e-16
+ wub = -2.4882066e-25
+ wuc = -1.434288e-17
+ wud = 0
+ lketa = 1.5671934e-8
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ paramchk = 1
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 2.4013086e-10
+ xpart = 1
+ rdsmod = 0
+ kt1l = 0
+ igbmod = 1
+ egidl = 0.001
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ lint = 0
+ poxedge = 1
+ pbswgd = 0.8
+ pbswgs = 0.8
+ lkt1 = 1.3151281e-8
+ lkt2 = 2.350723e-9
+ lmax = 5.4e-8
+ lmin = 4.5e-8
+ ijthdfwd = 0.01
+ igcmod = 1
+ binunit = 2
+ lpe0 = 6.44e-8
+ lpeb = 0
+ minv = -0.33
+ lua1 = -3.7660644e-16
+ lub1 = 5.1040674e-25
+ luc1 = -7.3441373e-17
+ ndep = 1e+18
+ lwlc = 0
+ ijthdrev = 0.01
+ moin = 5.5538
+ nigc = 2.291
+ lpdiblc2 = 0
+ pvoff = 4.4992157999999996e-17
+ cdscb = 0
+ cdscd = 0
+ pvsat = 1.1485877e-10
+ noff = 2.2684
+ wk2we = 0.0
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ pvth0 = 1.04221603e-16
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ permod = 1
+ drout = 0.56
+ paigc = -1.4334713e-18
+ voffl = 0
+ ntox = 1.0
+ pcit = -1.7599318000000002e-17
+ pclm = 1.8533357
+ weta0 = -4.4243037e-9
+ wetab = 2.5894049e-9
+ lpclm = -6.4524768e-8
+ lkvth0we = 3e-12
+ phin = 0.15
+ voffcv = -0.125
+ wpemod = 1
+ pkt1 = -1.6783146e-15
+ pkt2 = -1.1786798e-16
+ cgidl = 1
+ acnqsmod = 0
+ njtsswg = 6.489
+ rbdb = 50
+ pua1 = 1.8341764e-23
+ prwb = 0
+ pub1 = -1.3009877e-32
+ prwg = 0
+ puc1 = 9.9681375e-24
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ pbswd = 0.9
+ rbpb = 50
+ rbpd = 50
+ pbsws = 0.9
+ rbps = 50
+ rbodymod = 0
+ rbsb = 50
+ pvag = 2.1
+ ckappad = 0.6
+ ckappas = 0.6
+ rdsw = 200
+ pdiblc1 = 0
+ pdiblc2 = 0.0014658889
+ pdiblcb = 0
+ tpbswg = 0.001
+ pdits = 0
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ bigbacc = 0.0054401
+ ptvoff = -2.2999757e-17
+ pk2we = 0.0
+ wpdiblc2 = 1.4741467e-10
+ rshg = 14.1
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ waigsd = 1.9716411e-12
+ kvth0we = -0.00022
+ diomod = 1
+ tnoia = 0
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ pditsd = 0
+ pditsl = 0
+ vtsswgd = 1.1
+ peta0 = 2.03224906e-17
+ vtsswgs = 1.1
+ cjswgd = 1.7086399999999997e-10
+ pku0we = 0.0
+ cjswgs = 1.7086399999999997e-10
+ petab = -2.558443e-17
+ wketa = 3.409679e-8
+ tpbsw = 0.0025
+ tnom = 25
+ cjswd = 4.8144e-11
+ cjsws = 4.8144e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ tvfbsdoff = 0.1
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ wkvth0we = 0.0
+ mjswgd = 0.95
+ mjswgs = 0.95
+ wtvfbsdoff = 0
+ tcjswg = 0.00128
+ trnqsmod = 0
+ ltvfbsdoff = 0
+ wags = 2.5054667e-7
+ wcit = 2.7838518e-10
+ scref = 1e-6
+ voff = -0.1005239
+ pigcd = 2.572
+ acde = 0.5
+ aigsd = 0.0063632396
+ nfactor = 1
+ rgatemod = 0
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ tnjtsswg = 1
+ vsat = 101849.16
+ wint = 0
+ lvoff = -3.8177557e-9
+ vth0 = -0.24914034
+ fprout = 200
+ wkt1 = 3.6711578e-8
+ wkt2 = 3.2153756e-9
+ wmax = 2.674e-7
+ xrcrg1 = 12
+ xrcrg2 = 1
+ aigc = 0.0068691843
+ wmin = 1.08e-7
+ lvsat = -0.00042415496
+ lvth0 = -4.2146177e-9
+ ptvfbsdoff = 0
+ delta = 0.018814
+ laigc = -1.683393e-11
+ wtvoff = 5.2119196e-10
+ wua1 = -3.864028e-16
+ wub1 = 3.2172349e-25
+ wuc1 = -2.0479093e-16
+ rnoia = 0
+ rnoib = 0
+ a0 = 3.0243356
+ a1 = 0
+ a2 = 1
+ nigbacc = 10
+ b0 = 0
+ b1 = 0
+ at = -187272.02
+ cf = 8.17e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.021495622
+ k3 = -2.5823
+ em = 20000000.0
+ bigc = 0.0012521
+ ll = 0
+ lw = 0
+ u0 = -0.00054459259
+ w0 = 0
+ wwlc = 0
+ ua = -1.9655718e-9
+ ub = 1.5789686e-18
+ uc = -2.0243416e-10
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ pketa = -2.1465872e-15
+ ngate = 1.7e+20
+ ngcon = 1
+ capmod = 2
+ wpclm = -1.4226467e-7
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ wku0we = 1.5e-11
+ xtid = 3
+ xtis = 3
+ gbmin = 1e-12
+ nigbinv = 2.171
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigc = 0.15259
+ jswgd = 3.69e-13
+ mobmod = 0
+ jswgs = 3.69e-13
+ )

.model pch_sf_40 pmos (
+ level = 54
+ fnoimod = 1
+ dmcg = 3.1e-8
+ dmci = 3.1e-8
+ dmdg = 0
+ eigbinv = 1.1
+ laigsd = 6.1219753e-16
+ k2we = 5e-5
+ ijthsfwd = 0.01
+ tvoff = -0.00058332606
+ dsub = 0.5
+ dtox = 3.91e-10
+ xjbvd = 1
+ dvt0 = 3.48
+ dvt1 = 0.5088
+ dvt2 = -0.25
+ xjbvs = 1
+ lk2we = 0.0
+ eta0 = 0.11700471
+ alpha0 = 1.223e-8
+ alpha1 = 0.01
+ etab = -0.15063456
+ ijthsrev = 0.01
+ cigbacc = 0.245
+ ku0we = -0.0007
+ beta0 = 13.32
+ leta0 = 2.2591389e-9
+ letab = 4.3496496e-9
+ tnoimod = 0
+ ppclm = -3.5647768e-15
+ dlcig = 2.5e-9
+ cigbinv = 0.006
+ bgidl = 1834800000.0
+ ppdiblc2 = 0
+ toxref = 3e-9
+ version = 4.5
+ dmcgt = 0
+ tcjsw = 9.34e-5
+ tempmod = 0
+ ags = 1.2522222
+ cjd = 0.001270624
+ cit = -0.0077632099
+ cjs = 0.001270624
+ clc = 1e-7
+ cle = 0.6
+ bvd = 8.2
+ bvs = 8.2
+ dlc = 4.0349e-9
+ k3b = 2.1176
+ dwb = 0
+ dwc = 0
+ dwg = 0
+ dwj = 0
+ aigbacc = 0.012071
+ bigsd = 0.0003327
+ pkvth0we = 0.0
+ la0 = -3.4726683e-8
+ ltvoff = 1.026653e-10
+ jsd = 1.5e-7
+ jss = 1.5e-7
+ lat = 0.0010711306999999998
+ kt1 = -0.31430817
+ kt2 = -0.12562663
+ lk2 = 5.9641473e-9
+ wvoff = 3.3909703e-9
+ llc = 0
+ lln = 1
+ lu0 = 5.2721728e-10
+ mjd = 0.335
+ mjs = 0.335
+ lua = 9.0470184e-17
+ lub = -1.3836274e-26
+ luc = 2.7216576e-18
+ lud = 0
+ lwc = 0
+ lwl = 0
+ lwn = 1
+ njd = 1.02
+ njs = 1.02
+ pa0 = 1.4761752e-15
+ nsd = 1e+20
+ pbd = 0.75
+ pat = -5.6834015e-11
+ wvsat = -0.010288162
+ pbs = 0.75
+ pk2 = -2.7720832e-16
+ aigbinv = 0.009974
+ wvth0 = 2.2903735900000003e-9
+ pu0 = -6.1923224e-17
+ vfbsdoff = 0.01
+ prt = 0
+ pua = -4.2432063e-24
+ pub = -6.6397485e-33
+ puc = -1.7176927e-24
+ pud = 0
+ waigc = -4.0606639e-11
+ rsh = 15.2
+ tcj = 0.000832
+ ua1 = 2.1566906e-9
+ ub1 = -3.7269546e-18
+ pvfbsdoff = 0
+ uc1 = -1.7258848e-10
+ keta = 0.15497942
+ lku0we = 1.8e-11
+ tpb = 0.0016
+ wa0 = -1.421534e-7
+ epsrox = 3.9
+ ute = -1
+ wat = 0.002804707
+ web = 6628.3
+ wec = -16935.0
+ wk2 = 1.0175701e-8
+ wlc = 0
+ wln = 1
+ wu0 = 1.2726735e-9
+ xgl = -8.2e-9
+ xgw = 0
+ wua = 4.3503521e-18
+ wub = 1.8649442e-25
+ wuc = 4.6446086e-17
+ wud = 0
+ lketa = -7.3399177e-9
+ wwc = 0
+ wwl = 0
+ wwn = 1
+ paramchk = 1
+ jswd = 3.69e-13
+ jsws = 3.69e-13
+ lcit = 4.894380299999999e-10
+ xpart = 1
+ rdsmod = 0
+ kt1l = 0
+ igbmod = 1
+ egidl = 0.001
+ pscbe1 = 926400000.0
+ pscbe2 = 1e-20
+ lint = 0
+ poxedge = 1
+ pbswgd = 0.8
+ pbswgs = 0.8
+ lkt1 = 2.1163929e-9
+ lkt2 = 2.3369169e-9
+ lmax = 4.5e-8
+ lmin = 3.6e-8
+ ijthdfwd = 0.01
+ igcmod = 1
+ binunit = 2
+ lpe0 = 6.44e-8
+ lpeb = 0
+ minv = -0.33
+ lua1 = -7.3362164e-17
+ lub1 = 1.3390478e-25
+ luc1 = 1.4382206e-17
+ ndep = 1e+18
+ lwlc = 0
+ ijthdrev = 0.01
+ moin = 5.5538
+ nigc = 2.291
+ paigsd = -6.9790518e-23
+ lpdiblc2 = 0
+ pvoff = -1.14138231e-16
+ cdscb = 0
+ cdscd = 0
+ pvsat = 4.8577866e-10
+ noff = 2.2684
+ wk2we = 0.0
+ noia = 2.86e+42
+ noib = 2.5e+24
+ noic = 31000000000.0
+ pvth0 = -9.090969999999989e-18
+ jtsswgd = 1.75e-7
+ jtsswgs = 1.75e-7
+ permod = 1
+ drout = 0.56
+ paigc = 8.520035e-19
+ voffl = 0
+ ntox = 1.0
+ pcit = -1.8487562e-17
+ pclm = 0.41497396
+ weta0 = -1.051677e-9
+ wetab = 1.1541057e-8
+ lpclm = 5.9549575e-9
+ lkvth0we = 3e-12
+ phin = 0.15
+ voffcv = -0.125
+ wpemod = 1
+ pkt1 = -1.6740714e-15
+ pkt2 = -7.0509572e-16
+ cgidl = 1
+ acnqsmod = 0
+ njtsswg = 6.489
+ rbdb = 50
+ pua1 = 3.2441676e-23
+ prwb = 0
+ pub1 = -5.4663004e-32
+ prwg = 0
+ puc1 = -1.3788915e-24
+ xtsswgd = 0.32
+ xtsswgs = 0.32
+ pbswd = 0.9
+ rbpb = 50
+ rbpd = 50
+ pbsws = 0.9
+ rbps = 50
+ rbodymod = 0
+ rbsb = 50
+ pvag = 2.1
+ ckappad = 0.6
+ ckappas = 0.6
+ rdsw = 200
+ pdiblc1 = 0
+ pdiblc2 = 0.0014658889
+ pdiblcb = 0
+ tpbswg = 0.001
+ pdits = 0
+ cigsd = 0.013281
+ dvt0w = 0
+ dvt1w = 0
+ dvt2w = 0
+ bigbacc = 0.0054401
+ ptvoff = -3.9364956e-17
+ pk2we = 0.0
+ wpdiblc2 = 1.4741467e-10
+ rshg = 14.1
+ dvtp0 = 6e-7
+ dvtp1 = 0.5224
+ waigsd = 1.9730654e-12
+ kvth0we = -0.00022
+ diomod = 1
+ tnoia = 0
+ lintnoi = -5e-9
+ bigbinv = 0.00149
+ pditsd = 0
+ pditsl = 0
+ vtsswgd = 1.1
+ peta0 = -1.4493621999999998e-16
+ vtsswgs = 1.1
+ cjswgd = 1.7086399999999997e-10
+ pku0we = 0.0
+ cjswgs = 1.7086399999999997e-10
+ petab = -4.6421536e-16
+ wketa = -5.7187654e-8
+ tpbsw = 0.0025
+ tnom = 25
+ cjswd = 4.8144e-11
+ cjsws = 4.8144e-11
+ mjswd = 0.01
+ mjsws = 0.01
+ agidl = 3.2166e-9
+ tvfbsdoff = 0.1
+ toxe = 2.67e-9
+ toxm = 2.67e-9
+ wkvth0we = 0.0
+ mjswgd = 0.95
+ mjswgs = 0.95
+ wtvfbsdoff = 0
+ tcjswg = 0.00128
+ trnqsmod = 0
+ ltvfbsdoff = 0
+ wags = 2.5054667e-7
+ wcit = 2.9651259e-10
+ scref = 1e-6
+ voff = -0.12231559
+ pigcd = 2.572
+ acde = 0.5
+ aigsd = 0.0063632271
+ nfactor = 1
+ rgatemod = 0
+ wvfbsdoff = 0
+ lvfbsdoff = 0
+ tnjtsswg = 1
+ vsat = 151791.98
+ wint = 0
+ lvoff = -2.7499629e-9
+ vth0 = -0.31308607
+ fprout = 200
+ wkt1 = 3.6624982e-8
+ wkt2 = 1.5199615e-8
+ wmax = 2.674e-7
+ xrcrg1 = 12
+ xrcrg2 = 1
+ aigc = 0.0069354083
+ wmin = 1.08e-7
+ lvsat = -0.0028713534000000002
+ lvth0 = -1.0812769e-9
+ ptvfbsdoff = 0
+ delta = 0.018814
+ laigc = -2.0078906e-11
+ wtvoff = 8.5517561e-10
+ wua1 = -6.7415611e-16
+ wub1 = 1.1717873e-24
+ wuc1 = 2.6781086e-17
+ rnoia = 0
+ rnoib = 0
+ a0 = 0.69140412
+ a1 = 0
+ a2 = 1
+ nigbacc = 10
+ b0 = 0
+ b1 = 0
+ at = -30917.36
+ cf = 8.17e-11
+ ef = 1.15
+ k1 = 0.30425
+ k2 = -0.06369048
+ k3 = -2.5823
+ em = 20000000.0
+ bigc = 0.0012521
+ ll = 0
+ lw = 0
+ u0 = -0.0027875803
+ w0 = 0
+ wwlc = 0
+ ua = -2.1984191e-9
+ ub = 1.2906289e-18
+ uc = -1.4486626e-10
+ ud = 0
+ wl = 0
+ wr = 1
+ xj = 1.1e-7
+ xl = 4e-9
+ ww = 0
+ xw = 8.600000000000001e-9
+ pketa = 2.3263506e-15
+ ngate = 1.7e+20
+ ngcon = 1
+ capmod = 2
+ wpclm = 8.9861524e-8
+ cdsc = 0
+ cgbo = 0
+ cgdl = 3.0105e-11
+ cgdo = 2.6482e-11
+ wku0we = 1.5e-11
+ xtid = 3
+ xtis = 3
+ gbmin = 1e-12
+ nigbinv = 2.171
+ cgsl = 3.0105e-11
+ cgso = 2.6482e-11
+ cigc = 0.15259
+ jswgd = 3.69e-13
+ mobmod = 0
+ jswgs = 3.69e-13
+ )


