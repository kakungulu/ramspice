.model nch_ss_1 nmos (
+ level = 49
+ cjsw = 2.142574e-10
+ drout = 0.0
+ tpbsw = 0.001554306
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ cjswg = 3.507574e-10
+ pnfactor = 0.0
+ mjswg = 0.43879
+ wnfactor = 0.0
+ tnom = 25.0
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ wvoff = -6.32688e-10
+ pscbe1 = 200000030.0
+ pscbe2 = 1e-6
+ toxm = 4.08e-9
+ version = 3.24
+ pbsw = 0.6882682
+ pclm = 0.8000001
+ weta0 = 0
+ wvsat = 0.0
+ nqsmod = 0
+ lnfactor = 4.5192e-8
+ tpbswg = 0.001554306
+ wvth0 = 5.9653440000000004e-9
+ noimod = 2
+ ags = 0.02
+ keta = 0.009263485
+ cit = -0.00010000001
+ a0 = 0.3700794
+ a1 = 0.0
+ a2 = 0.99
+ b0 = 0.0
+ b1 = 0.0
+ dlc = 3e-9
+ dsub = 0.0
+ k3b = 0.0
+ at = 20000.0
+ cf = 0
+ cj = 0.001050279
+ ef = 0.874
+ k1 = 0.5142301
+ k2 = 0.022028564
+ k3 = 0.0
+ em = 30000000.0
+ dwb = 0.0
+ dwg = 0.0
+ js = 3.5e-7
+ ll = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ u0 = 0.04039571
+ pb = 0.6882682
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ dvt0 = 0.0
+ ua = -6.12274e-10
+ dvt1 = 0.0
+ ub = 2.3135539e-18
+ xpart = 1
+ dvt2 = 0.0
+ uc = 1.0876087e-10
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -1.3989464e-8
+ ww = 0.0
+ xw = -9.94224e-9
+ voff = -0.14328952
+ capmod = 3
+ ldif = 9e-8
+ pbswg = 0.6882682
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ jsw = 1.45e-12
+ kt1 = -0.2240464
+ lk2 = 3.6153600000000002e-9
+ kt2 = -0.030266136
+ lvoff = -9.038400000000001e-10
+ eta0 = 5e-5
+ llc = -0.039
+ lln = -1
+ pvag = 0.0
+ etab = -5e-5
+ lu0 = -4.5192000000000003e-10
+ vsat = 86384.65
+ beta0 = 11.59263
+ nch = 3.9e+17
+ wint = 3e-9
+ lwl = 0.0
+ lwn = 1.0
+ vth0 = 0.45508482
+ leta0 = 9.680916984722288e-19
+ mobmod = 1
+ nlx = 0.0
+ rdsw = 170.0
+ lint = 1e-8
+ wmax = 0.000900001
+ lvth0 = 2.621136e-9
+ pu0 = 0.0
+ wmin = 1.0009942240000001e-5
+ prt = 0
+ lmax = 2.0001e-5
+ delta = 0.01
+ lmin = 9.993989464000001e-6
+ rsh = 6.8
+ tcj = 0.001040287
+ ua1 = 1.224e-9
+ ub1 = -1.1209314e-18
+ uc1 = 1.1643822e-11
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ tpb = 0.001554306
+ tox = 4.14010536e-9
+ ute = -1.5799998
+ wln = 1.0
+ wu0 = 0.0
+ nfactor = 1.0
+ hdif = 2e-7
+ wwl = 0.0
+ wwn = 1
+ xti = 3
+ mjsw = 0.2003879
+ tcjswg = 0.000645489
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0006999999
+ pdiblcb = 0.01
+ tcjsw = 0.000645489
+ cdsc = 0.0
+ pvoff = -9.038400000000001e-16
+ cgdo = 3.48175e-10
+ binunit = 2
+ cgso = 3.48175e-10
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 4.148964422023837e-25
+ pvth0 = 2.71152e-15
+ )

.model nch_ss_2 nmos (
+ level = 49
+ wmax = 0.000900001
+ wmin = 1.0009942240000001e-5
+ lkt2 = -4.553491e-12
+ lmax = 9.993989464000001e-6
+ lmin = 1.193989464e-6
+ la0 = -3.496093e-7
+ jsw = 1.45e-12
+ kt1 = -0.2240468
+ lk1 = 1.4908844e-8
+ kt2 = -0.03026568
+ lk2 = -7.49802e-9
+ llc = -0.039
+ lln = -1
+ lketa = -4.320781e-8
+ lu0 = 2.8398890000000003e-9
+ lua = -4.643216e-16
+ lub = 7.375677e-25
+ luc = 3.898355e-17
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ xpart = 1
+ pnfactor = 0.0
+ nlx = 0.0
+ hdif = 2e-7
+ wnfactor = 0.0
+ capmod = 3
+ lub1 = 4.527317e-28
+ luc1 = 7.827772e-20
+ nfactor = 1.0
+ pu0 = 0.0
+ mjsw = 0.2003879
+ prt = 0
+ pbswg = 0.6882682
+ lute = -5.743953e-11
+ lvoff = -1.1375168e-8
+ rsh = 6.8
+ tcj = 0.001040287
+ ua1 = 1.224e-9
+ ub1 = -1.1209769e-18
+ uc1 = 1.1635963e-11
+ mobmod = 1
+ beta0 = 11.59263
+ tpb = 0.001554306
+ tox = 4.14010536e-9
+ lnfactor = 4.5192e-8
+ leta0 = 9.680916984722288e-19
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0003968181
+ cdsc = 0.0
+ pdiblcb = 0.01
+ lpscbe1 = 262.58185
+ ute = -1.5799941
+ lvsat = -0.006562638
+ cgdo = 3.48175e-10
+ wln = 1.0
+ lvth0 = 6.3234006e-8
+ wu0 = 0.0
+ wwl = 0.0
+ wwn = 1
+ cgso = 3.48175e-10
+ xti = 3
+ delta = 0.01
+ lpdiblc2 = 3.0196912e-9
+ binunit = 2
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ cjsw = 2.142574e-10
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ tnom = 25.0
+ tcjswg = 0.000645489
+ a0 = 0.4051808
+ a1 = 0.0
+ a2 = 0.99
+ b0 = 0.0
+ b1 = 0.0
+ at = 20000.0
+ cf = 0
+ cj = 0.001050279
+ ef = 0.874
+ k1 = 0.5127332
+ k2 = 0.023144367
+ k3 = 0.0
+ em = 30000000.0
+ toxm = 4.08e-9
+ js = 3.5e-7
+ ll = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ u0 = 0.040065210000000004
+ pb = 0.6882682
+ w0 = 0.0
+ pbsw = 0.6882682
+ rd = 0
+ pclm = 0.7736172
+ rs = 0
+ ua = -5.656554e-10
+ ub = 2.2395009e-18
+ uc = 1.0484686e-10
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -1.3989464e-8
+ ww = 0.0
+ xw = -9.94224e-9
+ tcjsw = 0.000645489
+ version = 3.24
+ pvoff = -9.038400000000001e-16
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 4.148964422023837e-25
+ pvth0 = 2.71152e-15
+ keta = 0.013601619
+ drout = 0.0
+ tpbsw = 0.001554306
+ dsub = 0.0
+ cjswg = 3.507574e-10
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ mjswg = 0.43879
+ pscbe1 = 173636400.0
+ pscbe2 = 1e-6
+ lcit = 2.6652053e-10
+ wvoff = -6.32688e-10
+ voff = -0.14223822
+ ldif = 9e-8
+ ags = 0.02
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ weta0 = 0
+ nqsmod = 0
+ eta0 = 5e-5
+ tpbswg = 0.001554306
+ pvag = 0.0
+ etab = -5e-5
+ cit = -0.00012675911
+ noimod = 2
+ wvsat = 0.0
+ vsat = 87043.55
+ wint = 3e-9
+ dlc = 3e-9
+ lpclm = 2.6277317e-7
+ wvth0 = 5.9653440000000004e-9
+ vth0 = 0.44899922
+ k3b = 0.0
+ rdsw = 170.0
+ dwb = 0.0
+ dwg = 0.0
+ lint = 1e-8
+ )

.model nch_ss_3 nmos (
+ level = 49
+ beta0 = 11.59263
+ leta0 = 3.8114280968091696e-11
+ letab = -3.811428e-11
+ lvsat = -0.0007622857
+ version = 3.24
+ lvth0 = 6.563892999999999e-9
+ delta = 0.01
+ keta = -0.015927497
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ dsub = 0.0
+ pnfactor = 0.0
+ lags = -3.044698e-8
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ tcjswg = 0.000645489
+ wnfactor = 0.0
+ lcit = 3.0262734e-10
+ voff = -0.16483012
+ ldif = 9e-8
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ eta0 = 1.7142866e-5
+ pvag = 0.0
+ etab = -1.7142866e-5
+ vsat = 82043.24
+ tcjsw = 0.000645489
+ lnfactor = 4.5192e-8
+ wint = 3e-9
+ vth0 = 0.49785271999999997
+ rdsw = 170.0
+ pvoff = -9.038400000000001e-16
+ lint = 1e-8
+ wmax = 0.000900001
+ wmin = 1.0009942240000001e-5
+ cdscb = 0.0
+ cdscd = 0.0
+ lkt1 = 5.782678e-9
+ lkt2 = 1.5570838e-9
+ peta0 = 4.148964422023837e-25
+ lmax = 1.193989464e-6
+ lpdiblc2 = 1.525682e-9
+ lmin = 4.93989464e-7
+ pvth0 = 2.71152e-15
+ ags = 0.0462474
+ drout = 0.0
+ tpbsw = 0.001554306
+ cit = -0.00015788565
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ dlc = 3e-9
+ cjswg = 3.507574e-10
+ k3b = 0.0
+ pscbe1 = 400000100.0
+ pscbe2 = 1e-6
+ mjswg = 0.43879
+ dwb = 0.0
+ dwg = 0.0
+ hdif = 2e-7
+ lua1 = -3.0446746e-18
+ lub1 = -1.2004175e-24
+ luc1 = -6.517273e-17
+ wvoff = -6.32688e-10
+ mjsw = 0.2003879
+ nqsmod = 0
+ tpbswg = 0.001554306
+ noimod = 2
+ nfactor = 1.0
+ lute = -2.6630502e-7
+ weta0 = 0
+ la0 = 4.581426e-7
+ wvsat = 0.0
+ jsw = 1.45e-12
+ kt1 = -0.2290285
+ lk1 = -7.214246e-9
+ kt2 = -0.031611919
+ lk2 = 5.318511e-9
+ lpclm = 1.5245718e-7
+ wvth0 = 5.9653440000000004e-9
+ a0 = -0.2911571
+ a1 = 0.0
+ a2 = 0.99
+ b0 = 0.0
+ b1 = 0.0
+ llc = -0.039
+ cdsc = 0.0
+ lln = -1
+ lu0 = 5.886878999999999e-10
+ at = 20000.0
+ cf = 0
+ cj = 0.001050279
+ ef = 0.874
+ k1 = 0.5318048
+ k2 = 0.012095633000000001
+ k3 = 0.0
+ em = 30000000.0
+ lua = 7.982966e-17
+ lub = -1.5630905e-25
+ luc = -9.669895e-18
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ js = 3.5e-7
+ cgdo = 3.48175e-10
+ ll = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0016847569
+ u0 = 0.0420059
+ pb = 0.6882682
+ w0 = 0.0
+ rd = 0
+ nlx = 0.0
+ rs = 0
+ pdiblcb = 0.01
+ ua = -1.0347512e-9
+ ub = 3.0100842e-18
+ uc = 1.4678947e-10
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -1.3989464e-8
+ ww = 0.0
+ xw = -9.94224e-9
+ cgso = 3.48175e-10
+ pu0 = 0.0
+ prt = 0
+ cjsw = 2.142574e-10
+ binunit = 2
+ rsh = 6.8
+ tcj = 0.001040287
+ ua1 = 1.2266247e-9
+ ub1 = -8.574386e-20
+ uc1 = 6.788683e-11
+ lketa = -8.954029e-9
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ tpb = 0.001554306
+ tox = 4.14010536e-9
+ capmod = 3
+ xpart = 1
+ ute = -1.3504703
+ tnom = 25.0
+ wln = 1.0
+ wu0 = 0.0
+ pbswg = 0.6882682
+ wwl = 0.0
+ wwn = 1
+ xti = 3
+ toxm = 4.08e-9
+ mobmod = 1
+ lvoff = 1.4831418000000001e-8
+ pbsw = 0.6882682
+ pclm = 0.8687172
+ )

.model nch_ss_4 nmos (
+ level = 49
+ lua1 = 8.039099e-19
+ lub1 = 3.824101e-25
+ luc1 = 2.9606131e-17
+ mjsw = 0.2003879
+ lute = 7.030476e-8
+ ags = -0.019916179
+ tcjsw = 0.000645489
+ nfactor = 1.0
+ cdsc = 0.0
+ cit = 0.000271889
+ pvoff = -9.038400000000001e-16
+ dlc = 3e-9
+ cgdo = 3.48175e-10
+ k3b = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cgso = 3.48175e-10
+ peta0 = 4.148964422023837e-25
+ pdiblc1 = 1e-6
+ pdiblc2 = -0.00593541
+ pdiblcb = 0.01
+ pvth0 = 2.71152e-15
+ drout = 0.0
+ alpha0 = 0.0
+ cjsw = 2.142574e-10
+ alpha1 = 0.448150714
+ tpbsw = 0.001554306
+ la0 = 7.545271e-8
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ pscbe1 = 400000000.0
+ pscbe2 = 1e-6
+ binunit = 2
+ jsw = 1.45e-12
+ kt1 = -0.22715
+ lk1 = 4.899558e-8
+ kt2 = -0.029537767
+ lk2 = -1.9725976e-8
+ cjswg = 3.507574e-10
+ pnfactor = 0.0
+ llc = -0.039
+ lln = -1
+ mjswg = 0.43879
+ lu0 = 7.998789e-10
+ wnfactor = 0.0
+ lua = -1.0530929e-18
+ lub = 5.559478e-27
+ luc = 4.133919e-18
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ tnom = 25.0
+ nqsmod = 0
+ tpbswg = 0.001554306
+ wvoff = -6.32688e-10
+ nlx = 0.0
+ noimod = 2
+ toxm = 4.08e-9
+ pu0 = 0.0
+ weta0 = 0
+ pbsw = 0.6882682
+ pclm = 1.1076791
+ prt = 0
+ wvsat = 0.0
+ lnfactor = 4.5192e-8
+ lpclm = 4.253467e-8
+ wvth0 = 5.9653440000000004e-9
+ rsh = 6.8
+ tcj = 0.001040287
+ ua1 = 1.2182583e-9
+ ub1 = -3.526674e-18
+ uc1 = -1.381542e-10
+ tpb = 0.001554306
+ tox = 4.14010536e-9
+ ute = -2.0822308
+ version = 3.24
+ wln = 1.0
+ wu0 = 0.0
+ lpdiblc2 = 5.030957e-9
+ wwl = 0.0
+ wwn = 1
+ xti = 3
+ keta = -0.04182327
+ capmod = 3
+ dsub = 0.0
+ lketa = 2.9580252e-9
+ xpart = 1
+ lags = -1.1735286e-11
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ lcit = 1.0493098e-10
+ voff = -0.12726132
+ pbswg = 0.6882682
+ mobmod = 1
+ ldif = 9e-8
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ lvoff = -2.4502018000000002e-9
+ eta0 = -0.0002937502
+ pvag = 0.0
+ etab = 0.0013875004
+ beta0 = 11.59263
+ vsat = 80823.6
+ wint = 3e-9
+ leta0 = 1.811250609680917e-10
+ vth0 = 0.49375982
+ letab = -6.842502e-10
+ rdsw = 170.0
+ lvsat = -0.00020125005
+ lint = 1e-8
+ lvth0 = 8.446637e-9
+ wmax = 0.000900001
+ wmin = 1.0009942240000001e-5
+ lkt1 = 4.918561e-9
+ lkt2 = 6.029743e-10
+ delta = 0.01
+ lmax = 4.93989464e-7
+ a0 = 0.5407774
+ a1 = 0.0
+ a2 = 0.99
+ b0 = 0.0
+ b1 = 0.0
+ lmin = 1.8e-7
+ at = 20000.0
+ cf = 0
+ cj = 0.001050279
+ ef = 0.874
+ k1 = 0.4096095
+ k2 = 0.06654018
+ k3 = 0.0
+ em = 30000000.0
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ js = 3.5e-7
+ ll = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ u0 = 0.04154679
+ pb = 0.6882682
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ua = -8.589192e-10
+ ub = 2.6581962e-18
+ uc = 1.1678118e-10
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -1.3989464e-8
+ ww = 0.0
+ xw = -9.94224e-9
+ tcjswg = 0.000645489
+ hdif = 2e-7
+ )

.model nch_ss_5 nmos (
+ level = 49
+ pu0 = 0.0
+ pscbe1 = 200000030.0
+ pscbe2 = 1e-6
+ tpbsw = 0.001554306
+ prt = 0
+ dsub = 0.0
+ cjswg = 3.507574e-10
+ rsh = 6.8
+ tcj = 0.001040287
+ ua1 = 1.224e-9
+ ub1 = -1.0684574e-18
+ a0 = 0.3702259
+ a1 = 0.0
+ a2 = 0.99
+ uc1 = 2.4230474e-11
+ b0 = 0.0
+ b1 = 0.0
+ mjswg = 0.43879
+ nqsmod = 0
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ tpbswg = 0.001554306
+ at = 20000.0
+ cf = 0
+ cj = 0.001050279
+ ef = 0.874
+ k1 = 0.5102321
+ k2 = 0.023322214
+ k3 = 0.0
+ tpb = 0.001554306
+ noimod = 2
+ em = 30000000.0
+ tox = 4.14010536e-9
+ js = 3.5e-7
+ wa0 = -1.4643313e-9
+ ll = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ wvoff = 2.5803440000000005e-10
+ u0 = 0.04122822
+ pb = 0.6882682
+ w0 = 0.0
+ rd = 0
+ ute = -1.5803809
+ rs = 0
+ ua = -5.885942e-10
+ ub = 2.3329335e-18
+ uc = 1.1057788e-10
+ voff = -0.14337861999999998
+ wk1 = 3.995606e-8
+ wk2 = -1.2928737e-8
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -1.3989464e-8
+ ww = 0.0
+ ldif = 9e-8
+ xw = -9.94224e-9
+ wln = 1.0
+ wu0 = -8.320099e-9
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ puc1 = -1.4905616e-28
+ weta0 = 0
+ wua = -2.3665659e-16
+ wub = -1.936796e-25
+ wuc = -1.815927e-17
+ wwl = 0.0
+ wwn = 1
+ eta0 = 5e-5
+ xti = 3
+ wvsat = 0.0
+ pvag = 0.0
+ etab = -5e-5
+ vsat = 86384.65
+ wvth0 = 6.652955400000001e-9
+ wint = 3e-9
+ vth0 = 0.45501602
+ rdsw = 170.0
+ wkt1 = -8.215166e-9
+ wkt2 = 1.6245854e-9
+ lint = 1e-8
+ wmax = 1.0009942240000001e-5
+ wmin = 1.20994224e-6
+ lmax = 2.0001e-5
+ lmin = 9.993989464000001e-6
+ capmod = 3
+ xpart = 1
+ wub1 = -5.244247e-25
+ pnfactor = 0.0
+ wuc1 = -1.257911e-16
+ wnfactor = 0.0
+ hdif = 2e-7
+ mobmod = 1
+ wute = 3.808433e-9
+ pbswg = 0.6882682
+ mjsw = 0.2003879
+ lvoff = -9.038400000000001e-10
+ beta0 = 11.59263
+ lnfactor = 4.5192e-8
+ leta0 = 9.680916984722288e-19
+ cdsc = 0.0
+ nfactor = 1.0
+ lvth0 = 2.621136e-9
+ cgdo = 3.48175e-10
+ cgso = 3.48175e-10
+ delta = 0.01
+ dvt0w = 0.0
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0006999999
+ dvt1w = 0.0
+ dvt2w = 0.0
+ pdiblcb = 0.01
+ cjsw = 2.142574e-10
+ tcjswg = 0.000645489
+ ags = 0.02
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ cit = -0.00010000001
+ binunit = 2
+ dlc = 3e-9
+ tnom = 25.0
+ k3b = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ toxm = 4.08e-9
+ pbsw = 0.6882682
+ pclm = 0.8000001
+ tcjsw = 0.000645489
+ pvoff = -9.038400000000001e-16
+ jsw = 1.45e-12
+ kt1 = -0.2232244
+ kt2 = -0.030428693
+ lk2 = 3.6153600000000002e-9
+ llc = -0.039
+ lln = -1
+ lu0 = -4.5192000000000003e-10
+ cdscb = 0.0
+ cdscd = 0.0
+ nch = 3.9e+17
+ peta0 = 4.148964422023837e-25
+ lwl = 0.0
+ lwn = 1.0
+ nlx = 0.0
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ version = 3.24
+ wketa = -1.0935369e-8
+ pvth0 = 2.71152e-15
+ keta = 0.010357677
+ drout = 0.0
+ )

.model nch_ss_6 nmos (
+ level = 49
+ nfactor = 1.0
+ cgso = 3.48175e-10
+ capmod = 3
+ cjsw = 2.142574e-10
+ lketa = -4.518989e-8
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0003968181
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ pdiblcb = 0.01
+ lpscbe1 = 262.58185
+ xpart = 1
+ mobmod = 1
+ tnom = 25.0
+ pbswg = 0.6882682
+ binunit = 2
+ toxm = 4.08e-9
+ lvoff = -1.1709891999999999e-8
+ a0 = 0.40626
+ a1 = 0.0
+ a2 = 0.99
+ b0 = 0.0
+ b1 = 0.0
+ pbsw = 0.6882682
+ pclm = 0.7755287
+ at = 20000.0
+ cf = 0
+ cj = 0.001050279
+ ef = 0.874
+ k1 = 0.508509
+ beta0 = 11.59263
+ k2 = 0.02454095
+ k3 = 0.0
+ em = 30000000.0
+ js = 3.5e-7
+ ll = 0.0
+ leta0 = 9.680916984722288e-19
+ mj = 0.3595262
+ lw = 0.0
+ u0 = 0.04092259
+ pb = 0.6882682
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ags = 0.02
+ ua = -5.377125e-10
+ ub = 2.2537915e-18
+ uc = 1.0657759e-10
+ lvsat = -0.006753025
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -1.3989464e-8
+ ww = 0.0
+ xw = -9.94224e-9
+ lvth0 = 6.3327226e-8
+ cit = -0.00012675911
+ ppclm = 1.9027247e-13
+ delta = 0.01
+ dlc = 3e-9
+ k3b = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ tcjswg = 0.000645489
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ pkt1 = 4.710912e-15
+ pkt2 = -4.130377e-15
+ keta = 0.014894814
+ version = 3.24
+ dsub = 0.0
+ pnfactor = 0.0
+ la0 = -3.588995e-7
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ wnfactor = 0.0
+ jsw = 1.45e-12
+ lk1 = 1.7161611e-8
+ kt1 = -0.2231775
+ lk2 = -8.523252e-9
+ kt2 = -0.030469729
+ pketa = 1.9809019e-14
+ llc = -0.039
+ lln = -1
+ lu0 = 2.5921712e-9
+ lcit = 2.6652053e-10
+ voff = -0.14229371999999998
+ lua = -5.067804e-16
+ lub = 7.882536e-25
+ luc = 3.984287e-17
+ nch = 3.9e+17
+ ldif = 9e-8
+ lwl = 0.0
+ lwn = 1.0
+ wpclm = -1.9103656e-8
+ kt1l = 0.0
+ pa0 = 9.284546e-14
+ prwb = 0.0
+ prwg = 0.0
+ pub1 = 4.176128e-31
+ nlx = 0.0
+ puc1 = 7.417578e-23
+ eta0 = 5e-5
+ pk1 = -2.2514154e-14
+ pk2 = 1.0246181e-14
+ pvag = 0.0
+ etab = -5e-5
+ tcjsw = 0.000645489
+ pu0 = 2.4756895e-15
+ vsat = 87062.66
+ lnfactor = 4.5192e-8
+ wint = 3e-9
+ pute = -5.708167e-14
+ prt = 0
+ pua = 4.243342e-22
+ pub = -5.065558e-31
+ puc = -8.588134e-24
+ vth0 = 0.44892112
+ rdsw = 170.0
+ pvoff = 2.441401e-15
+ wkt1 = -8.688151e-9
+ wkt2 = 2.0392819e-9
+ rsh = 6.8
+ lint = 1e-8
+ tcj = 0.001040287
+ ua1 = 1.224e-9
+ ub1 = -1.0643074e-18
+ uc1 = 2.4967807e-11
+ wmax = 1.0009942240000001e-5
+ wmin = 1.20994224e-6
+ cdscb = 0.0
+ cdscd = 0.0
+ tpb = 0.001554306
+ peta0 = 4.148964422023837e-25
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ tox = 4.14010536e-9
+ lkt1 = -4.674615e-10
+ lkt2 = 4.087321e-10
+ wa0 = -1.0786144e-8
+ lpdiblc2 = 3.0196912e-9
+ lmax = 9.993989464000001e-6
+ pvsat = 1.9027204e-9
+ ute = -1.5809486
+ pscbe1 = 173636400.0
+ pscbe2 = 1e-6
+ wk1 = 4.221652e-8
+ wk2 = -1.3957471e-8
+ lmin = 1.193989464e-6
+ wketa = -1.292423e-8
+ pvth0 = 1.7798325e-15
+ wln = 1.0
+ drout = 0.0
+ wu0 = -8.568663e-9
+ tpbsw = 0.001554306
+ wua = -2.7926046e-16
+ wub = -1.4282058e-25
+ wuc = -1.7297008e-17
+ wwl = 0.0
+ wwn = 1
+ xti = 3
+ nqsmod = 0
+ tpbswg = 0.001554306
+ cjswg = 3.507574e-10
+ noimod = 2
+ wub1 = -5.663537e-25
+ wuc1 = -1.3323848e-16
+ mjswg = 0.43879
+ hdif = 2e-7
+ wvoff = -7.783409999999999e-11
+ lub1 = -4.133362e-26
+ luc1 = -7.343755e-18
+ wute = 9.539526e-9
+ mjsw = 0.2003879
+ weta0 = 0
+ lute = 5.654154e-9
+ wvsat = -0.00019104627
+ lpclm = 2.4373449e-7
+ wvth0 = 6.7464942e-9
+ cdsc = 0.0
+ cgdo = 3.48175e-10
+ )

.model nch_ss_7 nmos (
+ level = 49
+ beta0 = 11.59263
+ pvag = 0.0
+ etab = -1.7142869e-5
+ vsat = 81898.23
+ leta0 = 3.8114280968091696e-11
+ wint = 3e-9
+ pute = 4.357466e-13
+ letab = -3.811428e-11
+ vth0 = 0.49852362
+ lvsat = -0.0007622865
+ rdsw = 170.0
+ lvth0 = 5.788268e-9
+ wkt1 = -3.681822e-9
+ wkt2 = -1.3190541e-9
+ lint = 1e-8
+ wmax = 1.0009942240000001e-5
+ la0 = 4.645035e-7
+ ppclm = 7.258032e-15
+ wmin = 1.20994224e-6
+ jsw = 1.45e-12
+ lk1 = -1.1179709e-8
+ kt1 = -0.2286601
+ lk2 = 7.0464250000000005e-9
+ kt2 = -0.031479932
+ delta = 0.01
+ tcjswg = 0.000645489
+ lkt1 = 5.892387e-9
+ lkt2 = 1.5805686e-9
+ llc = -0.039
+ lln = -1
+ lmax = 1.193989464e-6
+ lu0 = 5.085513000000001e-10
+ lmin = 4.93989464e-7
+ lua = 6.148926e-17
+ lub = -1.2783527e-25
+ luc = -6.505068e-18
+ nch = 3.9e+17
+ dvt0w = 0.0
+ lwl = 0.0
+ lwn = 1.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ pa0 = -6.357063e-14
+ nlx = 0.0
+ pk1 = 3.963084e-14
+ pk2 = -1.7268767e-14
+ pu0 = 8.008865e-16
+ prt = 0
+ pua = 1.8329395e-22
+ pub = -2.8456703e-31
+ puc = -3.16293e-23
+ wua1 = -3.55913e-18
+ wub1 = -1.6132161e-24
+ wuc1 = -1.8047248e-16
+ hdif = 2e-7
+ rsh = 6.8
+ pketa = 9.843987e-15
+ tcj = 0.001040287
+ ua1 = 1.2269809e-9
+ ub1 = 7.567455e-20
+ lua1 = -3.457781e-18
+ uc1 = 8.594492e-11
+ lub1 = -1.3637128e-24
+ luc1 = -7.807721e-17
+ wute = -4.153124e-7
+ mjsw = 0.2003879
+ tpb = 0.001554306
+ tox = 4.14010536e-9
+ wa0 = 1.2405528e-7
+ wpclm = 1.3866737e-7
+ ute = -1.3089141
+ lute = -3.0990586e-7
+ wk1 = -1.1356744e-8
+ wk2 = 9.762311e-9
+ wln = 1.0
+ tcjsw = 0.000645489
+ wu0 = -7.124867e-9
+ wua = -7.146715e-17
+ wub = -3.341902e-25
+ wuc = 2.5660584e-18
+ wwl = 0.0
+ wwn = 1
+ xti = 3
+ cdsc = 0.0
+ pvoff = -3.917654e-15
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ cgdo = 3.48175e-10
+ a0 = -0.3035701
+ a1 = 0.0
+ a2 = 0.99
+ b0 = 0.0
+ b1 = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 4.148964422023837e-25
+ at = 20000.0
+ cf = 0
+ cj = 0.001050279
+ pscbe1 = 400000100.0
+ pscbe2 = 1e-6
+ ef = 0.874
+ k1 = 0.5329412
+ k2 = 0.011118815
+ k3 = 0.0
+ em = 30000000.0
+ cgso = 3.48175e-10
+ js = 3.5e-7
+ ll = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ u0 = 0.04271881
+ pb = 0.6882682
+ nfactor = 1.0
+ w0 = 0.0
+ rd = 0
+ wketa = -4.333682e-9
+ rs = 0
+ ua = -1.0276002e-9
+ ub = 3.0435232e-18
+ uc = 1.4653272e-10
+ pvth0 = 1.0463117999999999e-14
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -1.3989464e-8
+ ww = 0.0
+ xw = -9.94224e-9
+ drout = 0.0
+ tpbsw = 0.001554306
+ nqsmod = 0
+ cjsw = 2.142574e-10
+ tpbswg = 0.001554306
+ noimod = 2
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ cjswg = 3.507574e-10
+ pnfactor = 0.0
+ mjswg = 0.43879
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0017737894
+ pdiblcb = 0.01
+ wnfactor = 0.0
+ tnom = 25.0
+ wvoff = 5.40411e-9
+ pags = 4.128623e-14
+ toxm = 4.08e-9
+ weta0 = 0
+ ppdiblc2 = 1.0321563e-15
+ binunit = 2
+ pbsw = 0.6882682
+ pclm = 0.8548421
+ wvsat = 0.0014492224
+ wpdiblc2 = -8.897895e-10
+ lpclm = 1.5173094e-7
+ wvth0 = -7.390919999999996e-10
+ lnfactor = 4.5192e-8
+ capmod = 3
+ lpdiblc2 = 1.4224044e-9
+ pkt1 = -1.0964308e-15
+ pkt2 = -2.3470743e-16
+ keta = -0.01549387
+ lketa = -9.939018e-9
+ mobmod = 1
+ wags = -3.559157e-8
+ dsub = 0.0
+ version = 3.24
+ xpart = 1
+ ags = 0.04980868
+ lags = -3.457808e-8
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ cit = -0.00015788565
+ pbswg = 0.6882682
+ lcit = 3.0262734e-10
+ voff = -0.16543412
+ ldif = 9e-8
+ dlc = 3e-9
+ k3b = 0.0
+ kt1l = 0.0
+ lvoff = 1.5132981999999998e-8
+ pua1 = 4.128591e-24
+ prwb = 0.0
+ prwg = 0.0
+ pub1 = 1.6319734e-30
+ puc1 = 1.2896722e-22
+ dwb = 0.0
+ dwg = 0.0
+ eta0 = 1.7142869e-5
+ )

.model nch_ss_8 nmos (
+ level = 49
+ pketa = -2.7027957e-15
+ tnom = 25.0
+ pdiblc1 = 1e-6
+ pdiblc2 = -0.006119013
+ pdiblcb = 0.01
+ pags = -1.0838496e-14
+ toxm = 4.08e-9
+ wpclm = 6.656068e-8
+ pcit = 1.4220811e-17
+ pbsw = 0.6882682
+ pclm = 1.1010191
+ tcjsw = 0.000645489
+ binunit = 2
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ pvoff = -1.8792550000000002e-15
+ pscbe1 = 400000000.0
+ pscbe2 = 1e-6
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = -1.3821213851035578e-18
+ petab = 1.6959704e-18
+ pvsat = 1.5350395e-12
+ wketa = 2.2941933e-8
+ nqsmod = 0
+ pvth0 = 7.220458e-15
+ tpbswg = 0.001554306
+ drout = 0.0
+ noimod = 2
+ pkt1 = -1.7512235e-15
+ pkt2 = 7.382567e-17
+ keta = -0.04411884
+ tpbsw = 0.001554306
+ wags = 7.772305e-8
+ dsub = 0.0
+ cjswg = 3.507574e-10
+ mjswg = 0.43879
+ lags = 1.0727657e-9
+ wcit = -3.0914837e-11
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ version = 3.24
+ wvoff = 9.728084e-10
+ lcit = 1.0350804e-10
+ voff = -0.12742202
+ ldif = 9e-8
+ weta0 = 3.0046217e-12
+ kt1l = 0.0
+ pua1 = -1.0901051e-24
+ prwb = 0.0
+ prwg = 0.0
+ pub1 = -4.238914e-31
+ puc1 = -2.7204607e-23
+ wetab = -3.686654e-12
+ wvsat = 0.0014459029
+ eta0 = -0.00029405078
+ pvag = 0.0
+ etab = 0.0013878694
+ lpclm = 3.848953e-8
+ wvth0 = 6.3101676e-9
+ vsat = 80678.92
+ wint = 3e-9
+ pute = -1.178615e-13
+ vth0 = 0.49372532
+ rdsw = 170.0
+ capmod = 3
+ wkt1 = -2.2583577e-9
+ wkt2 = -1.9897783e-9
+ lint = 1e-8
+ ags = -0.027693154
+ wmax = 1.0009942240000001e-5
+ wmin = 1.20994224e-6
+ lkt1 = 5.093789e-9
+ lkt2 = 5.955873e-10
+ lmax = 4.93989464e-7
+ cit = 0.00027498236
+ lmin = 1.8e-7
+ dlc = 3e-9
+ mobmod = 1
+ k3b = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ a0 = 0.5262308
+ a1 = 0.0
+ a2 = 0.99
+ lketa = 3.228467e-9
+ b0 = 0.0
+ b1 = 0.0
+ at = 20000.0
+ cf = 0
+ cj = 0.001050279
+ ef = 0.874
+ k1 = 0.4007356
+ k2 = 0.07041932
+ k3 = 0.0
+ em = 30000000.0
+ xpart = 1
+ js = 3.5e-7
+ ll = 0.0
+ pnfactor = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ u0 = 0.04203316
+ wua1 = 7.785862e-18
+ pb = 0.6882682
+ wub1 = 2.8560549e-24
+ w0 = 0.0
+ wuc1 = 1.5903152e-16
+ rd = 0
+ rs = 0
+ ua = -9.017296e-10
+ ub = 2.7527719e-18
+ uc = 1.2291169e-10
+ wnfactor = 0.0
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -1.3989464e-8
+ ww = 0.0
+ xw = -9.94224e-9
+ hdif = 2e-7
+ lua1 = 9.129858e-19
+ lub1 = 4.248247e-25
+ la0 = 8.279508e-8
+ luc1 = 3.232822e-17
+ pbswg = 0.6882682
+ wute = 7.881835e-7
+ mjsw = 0.2003879
+ jsw = 1.45e-12
+ lk1 = 4.963488e-8
+ kt1 = -0.226924
+ lk2 = -2.0231804000000002e-8
+ kt2 = -0.029338669
+ llc = -0.039
+ lvoff = -2.3526017e-9
+ lln = -1
+ lu0 = 8.239492e-10
+ ppdiblc2 = -2.2121929e-16
+ lute = 8.209799e-8
+ lua = 3.588764e-18
+ lub = 5.910339e-27
+ luc = 4.360599e-18
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ wpdiblc2 = 1.8349379e-9
+ beta0 = 11.59263
+ pa0 = -7.337964e-14
+ lnfactor = 4.5192e-8
+ nlx = 0.0
+ leta0 = 1.812633409680917e-10
+ letab = -6.844199e-10
+ pk1 = -6.389182e-15
+ pk2 = 5.055259e-15
+ lvsat = -0.00020140363
+ cdsc = 0.0
+ pu0 = -2.4055863e-16
+ lvth0 = 7.995472e-9
+ prt = 0
+ pua = -4.639069e-23
+ pub = -3.506499e-33
+ puc = -2.2654354e-24
+ cgdo = 3.48175e-10
+ tcjswg = 0.000645489
+ ppclm = 4.042711e-14
+ delta = 0.01
+ cgso = 3.48175e-10
+ rsh = 6.8
+ tcj = 0.001040287
+ lpdiblc2 = 5.053093e-9
+ ua1 = 1.2174792e-9
+ ub1 = -3.81245e-18
+ uc1 = -1.540669e-10
+ tpb = 0.001554306
+ tox = 4.14010536e-9
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ wa0 = 1.4537927e-7
+ nfactor = 1.0
+ ute = -2.1610963
+ cjsw = 2.142574e-10
+ wk1 = 8.868675e-8
+ wk2 = -3.876818e-8
+ wln = 1.0
+ wu0 = -4.860856e-9
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ wua = 4.278473e-16
+ wub = -9.451913e-25
+ wuc = -6.126842e-17
+ wwl = 0.0
+ wwn = 1
+ xti = 3
+ )

.model nch_ss_9 nmos (
+ level = 49
+ cjswg = 3.507574e-10
+ mjswg = 0.43879
+ wub1 = -7.675553e-27
+ wuc1 = -1.4706552e-17
+ hdif = 2e-7
+ wvoff = -1.499257e-9
+ ags = 0.02
+ wute = 3.836007e-8
+ mjsw = 0.2003879
+ weta0 = 0
+ cit = -0.00010000004
+ wvsat = 0.0
+ dlc = 3e-9
+ k3b = 0.0
+ wvth0 = 1.7022350000000006e-9
+ dwb = 0.0
+ dwg = 0.0
+ capmod = 3
+ cdsc = 0.0
+ cgdo = 3.48175e-10
+ cgso = 3.48175e-10
+ mobmod = 1
+ jsw = 1.45e-12
+ kt1 = -0.2313184
+ lk2 = 3.6153600000000002e-9
+ kt2 = -0.029076951
+ llc = -0.039
+ lln = -1
+ lu0 = -4.5192000000000003e-10
+ cjsw = 2.142574e-10
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ nlx = 0.0
+ nfactor = 1.0
+ xpart = 1
+ pu0 = 0.0
+ prt = 0
+ tnom = 25.0
+ pbswg = 0.6882682
+ rsh = 6.8
+ tcj = 0.001040287
+ ua1 = 1.224e-9
+ pdiblc1 = 1e-6
+ toxm = 4.08e-9
+ pdiblc2 = 0.0007000003
+ ub1 = -1.5012456e-18
+ lvoff = -9.038400000000001e-10
+ uc1 = -6.880516e-11
+ pdiblcb = 0.01
+ pbsw = 0.6882682
+ tpb = 0.001554306
+ pclm = 0.8000001
+ tox = 4.14010536e-9
+ beta0 = 11.59263
+ wa0 = 7.667051e-8
+ leta0 = 9.680916984722288e-19
+ ute = -1.6093186
+ wk1 = -2.074723e-8
+ wk2 = 4.920634e-9
+ tcjswg = 0.000645489
+ wln = 1.0
+ wu0 = 1.0362965e-9
+ lvth0 = 2.621136e-9
+ binunit = 2
+ wua = 1.4309126e-16
+ wub = -1.5411778e-25
+ wuc = -1.4141237e-17
+ wwl = 0.0
+ wwn = 1
+ xti = 3
+ delta = 0.01
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ keta = 0.0010152902
+ dsub = 0.0
+ pnfactor = 0.0
+ wnfactor = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ a0 = 0.3047864
+ a1 = 0.0
+ a2 = 0.99
+ b0 = 0.0
+ b1 = 0.0
+ voff = -0.14190692
+ version = 3.24
+ at = 20000.0
+ cf = 0
+ cj = 0.001050279
+ ldif = 9e-8
+ ef = 0.874
+ k1 = 0.5610723
+ k2 = 0.0083729917
+ k3 = 0.0
+ em = 30000000.0
+ kt1l = 0.0
+ js = 3.5e-7
+ prwb = 0.0
+ ll = 0.0
+ prwg = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ u0 = 0.03339204
+ pb = 0.6882682
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ua = -9.066409e-10
+ ub = 2.2997995e-18
+ uc = 1.072127e-10
+ eta0 = 5e-5
+ wl = 0.0
+ tcjsw = 0.000645489
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -1.3989464e-8
+ ww = 0.0
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ xw = -9.94224e-9
+ pvag = 0.0
+ etab = -5e-5
+ lnfactor = 4.5192e-8
+ vsat = 86384.65
+ wint = 3e-9
+ pscbe1 = 200000030.0
+ pscbe2 = 1e-6
+ vth0 = 0.45916242
+ pvoff = -9.038400000000001e-16
+ rdsw = 170.0
+ wkt1 = 1.4490446e-9
+ wkt2 = 1.0605161e-11
+ lint = 1e-8
+ wmax = 1.20994224e-6
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 4.148964422023837e-25
+ wmin = 5.0994224e-7
+ nqsmod = 0
+ tpbswg = 0.001554306
+ noimod = 2
+ lmax = 2.0001e-5
+ wketa = 2.1944087e-10
+ pvth0 = 2.71152e-15
+ lmin = 9.993989464000001e-6
+ drout = 0.0
+ tpbsw = 0.001554306
+ )

.model nch_ss_10 nmos (
+ level = 49
+ lute = -1.2190513e-8
+ nqsmod = 0
+ tpbswg = 0.001554306
+ noimod = 2
+ cdsc = 0.0
+ cgdo = 3.48175e-10
+ nfactor = 1.0
+ lketa = -2.8027248e-8
+ cgso = 3.48175e-10
+ xpart = 1
+ cjsw = 2.142574e-10
+ pbswg = 0.6882682
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0003968185
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ pdiblcb = 0.01
+ lpscbe1 = 262.58185
+ lvoff = -4.506062e-9
+ capmod = 3
+ beta0 = 11.59263
+ tnom = 25.0
+ leta0 = 9.680916984722288e-19
+ binunit = 2
+ lvsat = -0.006201102
+ toxm = 4.08e-9
+ lvth0 = 6.8541616e-8
+ pcit = 4.302753e-19
+ pbsw = 0.6882682
+ pclm = 0.7699873
+ ppclm = 1.243718e-13
+ mobmod = 1
+ delta = 0.01
+ ags = 0.02
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ cit = -0.00012672294
+ dlc = 3e-9
+ k3b = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ pnfactor = 0.0
+ pkt1 = 7.833639e-15
+ pkt2 = 9.747044e-16
+ keta = 0.00382927
+ wnfactor = 0.0
+ pketa = -6.831802e-16
+ version = 3.24
+ dsub = 0.0
+ wpclm = -1.2487239e-8
+ wcit = -4.317371e-14
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ la0 = -1.9725388e-7
+ tcjsw = 0.000645489
+ jsw = 1.45e-12
+ tcjswg = 0.000645489
+ lk1 = 1.0512358e-8
+ kt1 = -0.2310088
+ lk2 = -1.7946909999999996e-9
+ kt2 = -0.028688708
+ lcit = 2.6616018e-10
+ llc = -0.039
+ lln = -1
+ voff = -0.14154522
+ lu0 = 3.253832e-9
+ lnfactor = 4.5192e-8
+ ldif = 9e-8
+ lua = -1.9124487e-16
+ lub = 4.117038e-25
+ luc = 4.038815e-17
+ nch = 3.9e+17
+ pvoff = -6.159972e-15
+ lwl = 0.0
+ lwn = 1.0
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ pub1 = -1.8996434e-32
+ puc1 = 1.3569954e-23
+ pa0 = -1.0015934e-13
+ nlx = 0.0
+ eta0 = 5e-5
+ pk1 = -1.457495e-14
+ pk2 = 2.2122807e-15
+ pvag = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ etab = -5e-5
+ peta0 = 4.148964422023837e-25
+ vsat = 87007.25
+ wint = 3e-9
+ pu0 = 1.6856667e-15
+ pute = -3.577514e-14
+ pvsat = 1.2437262e-9
+ vth0 = 0.45254382
+ prt = 0
+ pua = 4.758471e-23
+ pub = -5.695533e-32
+ puc = -9.239189e-24
+ lpdiblc2 = 3.0196912e-9
+ wketa = 2.8803285e-10
+ rdsw = 170.0
+ pvth0 = -4.446152000000001e-15
+ wkt1 = 6.625341e-10
+ wkt2 = -8.725676e-11
+ drout = 0.0
+ lint = 1e-8
+ rsh = 6.8
+ tpbsw = 0.001554306
+ wmax = 1.20994224e-6
+ tcj = 0.001040287
+ ua1 = 1.224e-9
+ ub1 = -1.5338095e-18
+ uc1 = -7.316409e-11
+ wmin = 5.0994224e-7
+ lkt1 = -3.0828107e-9
+ lkt2 = -3.866881e-9
+ tpb = 0.001554306
+ tox = 4.14010536e-9
+ cjswg = 3.507574e-10
+ lmax = 9.993989464000001e-6
+ wa0 = 8.672666e-8
+ lmin = 1.193989464e-6
+ ute = -1.6080947
+ mjswg = 0.43879
+ wk1 = -1.9283881e-8
+ wk2 = 4.698517e-9
+ wln = 1.0
+ wu0 = 8.670528e-10
+ wvoff = -9.715325e-10
+ wua = 1.3831368e-16
+ wub = -1.4839938e-25
+ wuc = -1.3213606e-17
+ wwl = 0.0
+ wwn = 1
+ xti = 3
+ a0 = 0.324591
+ a1 = 0.0
+ a2 = 0.99
+ b0 = 0.0
+ b1 = 0.0
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ wub1 = -5.768295e-27
+ wuc1 = -1.6068998e-17
+ weta0 = 0
+ at = 20000.0
+ cf = 0
+ cj = 0.001050279
+ ef = 0.874
+ k1 = 0.5600169
+ k2 = 0.008916168700000001
+ k3 = 0.0
+ em = 30000000.0
+ hdif = 2e-7
+ wvsat = -0.00012487893
+ js = 3.5e-7
+ pscbe1 = 173636400.0
+ pscbe2 = 1e-6
+ ll = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ u0 = 0.033019980000000004
+ pb = 0.6882682
+ lub1 = 3.243357e-25
+ lpclm = 2.9892766e-7
+ wvth0 = 2.4208780000000006e-9
+ luc1 = 4.341489e-17
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ wute = 4.195195e-8
+ ua = -8.874397e-10
+ ub = 2.2584638e-18
+ uc = 1.0315766e-10
+ mjsw = 0.2003879
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -1.3989464e-8
+ ww = 0.0
+ xw = -9.94224e-9
+ )

.model nch_ss_11 nmos (
+ level = 49
+ lvoff = 1.025939e-8
+ wcit = 5.431231e-13
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ ags = 0.02
+ beta0 = 11.59263
+ leta0 = 3.8114300968091695e-11
+ lcit = 3.0283653e-10
+ cit = -0.0001583405
+ letab = -3.81143e-11
+ voff = -0.15427401999999998
+ ldif = 9e-8
+ lvsat = -0.0007659488
+ dlc = 3e-9
+ kt1l = 0.0
+ mobmod = 1
+ prwb = 0.0
+ lvth0 = 1.2730886999999999e-8
+ prwg = 0.0
+ pub1 = -5.874811e-31
+ puc1 = -3.67348e-23
+ a0 = -0.1914371
+ a1 = 0.0
+ a2 = 0.99
+ k3b = 0.0
+ b0 = 0.0
+ b1 = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ eta0 = 1.7142847e-5
+ at = 20000.0
+ cf = 0
+ cj = 0.001050279
+ ef = 0.874
+ k1 = 0.5552615
+ ppclm = 7.308824e-14
+ k2 = 0.010775519
+ k3 = 0.0
+ em = 30000000.0
+ pvag = 0.0
+ etab = -1.7142847e-5
+ delta = 0.01
+ js = 3.5e-7
+ vsat = 82321.77
+ ll = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ u0 = 0.03400418
+ pb = 0.6882682
+ wint = 3e-9
+ pute = -2.0303331e-13
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ua = -1.3333591e-9
+ ub = 2.969086e-18
+ uc = 1.6160392e-10
+ vth0 = 0.50065652
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -1.3989464e-8
+ ww = 0.0
+ xw = -9.94224e-9
+ rdsw = 170.0
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ wkt1 = 1.1898274e-8
+ wkt2 = 2.0987987e-9
+ lint = 1e-8
+ wmax = 1.20994224e-6
+ la0 = 4.013388e-7
+ wmin = 5.0994224e-7
+ lkt1 = 9.329063e-9
+ lkt2 = 2.691467e-9
+ jsw = 1.45e-12
+ lk1 = 1.6028618e-8
+ kt1 = -0.2417087
+ lk2 = -3.9515360000000006e-9
+ kt2 = -0.03434246
+ lmax = 1.193989464e-6
+ llc = -0.039
+ lln = -1
+ lu0 = 2.1121620999999997e-9
+ lmin = 4.93989464e-7
+ lua = 3.260216e-16
+ lub = -4.12618e-25
+ luc = -2.7409531e-17
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ pketa = 1.4501565e-15
+ pa0 = 1.1848049e-14
+ nlx = 0.0
+ pk1 = 7.144098e-15
+ pk2 = -4.137203e-15
+ pu0 = -1.1138246e-15
+ wpclm = 3.172275e-8
+ wub1 = 4.843047e-25
+ prt = 0
+ wuc1 = 2.7297169e-17
+ pua = -1.3255767e-22
+ pub = 5.546348e-32
+ puc = -6.669366e-24
+ tcjswg = 0.000645489
+ hdif = 2e-7
+ tcjsw = 0.000645489
+ rsh = 6.8
+ lub1 = 4.951269e-25
+ luc1 = 6.070172e-17
+ tcj = 0.001040287
+ ua1 = 1.224e-9
+ ub1 = -1.6810433e-18
+ uc1 = -8.806652e-11
+ wute = 1.8614003e-7
+ mjsw = 0.2003879
+ pvoff = 1.9014135e-15
+ tpb = 0.001554306
+ tox = 4.14010536e-9
+ wa0 = -9.831444e-9
+ lute = 2.2508574e-7
+ ute = -1.8126432
+ wk1 = -3.80072e-8
+ wk2 = 1.0172209e-8
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 4.148964422023837e-25
+ wln = 1.0
+ wu0 = 3.280407e-9
+ wua = 2.9360883e-16
+ pvsat = 4.380818e-12
+ wub = -2.4531215e-25
+ wuc = -1.542897e-17
+ wwl = 0.0
+ wwn = 1
+ cdsc = 0.0
+ wketa = -1.5510503e-9
+ pvth0 = 2.1736318e-15
+ xti = 3
+ drout = 0.0
+ cgdo = 3.48175e-10
+ tpbsw = 0.001554306
+ cgso = 3.48175e-10
+ cjswg = 3.507574e-10
+ nfactor = 1.0
+ mjswg = 0.43879
+ pnfactor = 0.0
+ cjsw = 2.142574e-10
+ wnfactor = 0.0
+ wvoff = -7.921003e-9
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ weta0 = 0
+ pscbe1 = 400000100.0
+ pscbe2 = 1e-6
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0011219129
+ pdiblcb = 0.01
+ wvsat = 0.0009435224
+ ppdiblc2 = 1.2928064e-16
+ tnom = 25.0
+ lpclm = 9.659676e-8
+ wvth0 = -3.2858339999999996e-9
+ wpdiblc2 = -1.1144895e-10
+ lnfactor = 4.5192e-8
+ nqsmod = 0
+ tpbswg = 0.001554306
+ toxm = 4.08e-9
+ noimod = 2
+ pcit = -2.4980728e-19
+ binunit = 2
+ pbsw = 0.6882682
+ pclm = 0.9444105
+ lpdiblc2 = 2.1785818e-9
+ lketa = -2.9090079e-9
+ xpart = 1
+ pkt1 = -5.199821e-15
+ pkt2 = -1.5611203e-15
+ keta = -0.017824383
+ pbswg = 0.6882682
+ dsub = 0.0
+ capmod = 3
+ version = 3.24
+ )

.model nch_ss_12 nmos (
+ level = 49
+ tpb = 0.001554306
+ tox = 4.14010536e-9
+ wa0 = 1.7605426e-7
+ pketa = -7.367843e-16
+ cjsw = 2.142574e-10
+ nfactor = 1.0
+ ute = -1.2073984
+ wk1 = -1.7855582e-8
+ wk2 = 1.6966123e-9
+ tcjswg = 0.000645489
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ wln = 1.0
+ wu0 = -4.268465e-11
+ wpclm = 1.9327061e-7
+ wua = -1.9101984e-17
+ wub = -5.11281e-26
+ wuc = -9.012729e-18
+ wwl = 0.0
+ wwn = 1
+ xti = 3
+ tcjsw = 0.000645489
+ tnom = 25.0
+ pdiblc1 = 1e-6
+ pdiblc2 = -0.00401322
+ pags = 1.8981756e-15
+ pdiblcb = 0.01
+ pvoff = -3.1245874000000002e-15
+ toxm = 4.08e-9
+ pcit = -1.4232223e-17
+ pbsw = 0.6882682
+ pclm = 0.9948969
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = -1.1371990585103558e-17
+ petab = 1.3954016e-17
+ binunit = 2
+ pvsat = 1.606088e-11
+ wketa = 3.203169e-9
+ pvth0 = 5.427536e-15
+ drout = 0.0
+ tpbsw = 0.001554306
+ a0 = 0.5005398
+ a1 = 0.0
+ a2 = 0.99
+ b0 = 0.0
+ b1 = 0.0
+ at = 20000.0
+ cf = 0
+ cj = 0.001050279
+ ef = 0.874
+ k1 = 0.489967
+ k2 = 0.036529204
+ k3 = 0.0
+ em = 30000000.0
+ js = 3.5e-7
+ cjswg = 3.507574e-10
+ ll = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ u0 = 0.03799784
+ pb = 0.6882682
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ua = -5.274002e-10
+ ub = 2.0039751e-18
+ uc = 7.914647e-11
+ mjswg = 0.43879
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -1.3989464e-8
+ ww = 0.0
+ xw = -9.94224e-9
+ pkt1 = 2.3961372e-15
+ pkt2 = 8.832021e-16
+ keta = -0.027587207
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ wvoff = 3.005086e-9
+ wags = -4.12647e-9
+ dsub = 0.0
+ pscbe1 = 400000000.0
+ pscbe2 = 1e-6
+ weta0 = 2.4721704e-11
+ lags = -9.594464e-9
+ wetab = -3.0334849e-11
+ wcit = 3.093965e-11
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ wvsat = 0.000918131
+ version = 3.24
+ nqsmod = 0
+ lpclm = 7.337301e-8
+ wvth0 = -1.0359539e-8
+ tpbswg = 0.001554306
+ noimod = 2
+ lcit = 1.2733804e-10
+ voff = -0.12912402
+ ldif = 9e-8
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ pub1 = 1.6165291e-31
+ puc1 = 2.0250814e-23
+ eta0 = -0.00031223928
+ pvag = 0.0
+ etab = 0.0014101875
+ vsat = 81120.94
+ wint = 3e-9
+ pute = 4.383575e-14
+ vth0 = 0.50768662
+ rdsw = 170.0
+ wkt1 = -4.614678e-9
+ wkt2 = -3.214946e-9
+ lint = 1e-8
+ wmax = 1.20994224e-6
+ ags = 0.04085753
+ lketa = 1.5818911e-9
+ wmin = 5.0994224e-7
+ lkt1 = 1.6202869e-9
+ lkt2 = -8.228257e-11
+ lmax = 4.93989464e-7
+ xpart = 1
+ cit = 0.00022317801
+ lmin = 1.8e-7
+ pnfactor = 0.0
+ dlc = 3e-9
+ wnfactor = 0.0
+ k3b = 0.0
+ capmod = 3
+ dwb = 0.0
+ dwg = 0.0
+ pbswg = 0.6882682
+ lvoff = -1.3096095e-9
+ wub1 = -1.1442477e-24
+ wuc1 = -9.658459e-17
+ ppdiblc2 = 3.905237e-16
+ hdif = 2e-7
+ beta0 = 11.59263
+ wpdiblc2 = -6.793707e-10
+ lub1 = -6.558089e-26
+ leta0 = 1.8963006096809171e-10
+ luc1 = -7.416688e-18
+ wute = -3.505318e-7
+ mobmod = 1
+ la0 = 8.302936e-8
+ letab = -6.946862e-10
+ lnfactor = 4.5192e-8
+ mjsw = 0.2003879
+ lvsat = -0.00021356932
+ jsw = 1.45e-12
+ lk1 = 4.606408e-8
+ kt1 = -0.2249505
+ lk2 = -1.5798233e-8
+ kt2 = -0.028312566
+ lvth0 = 9.497081e-9
+ llc = -0.039
+ lln = -1
+ lute = -5.332685e-8
+ lu0 = 2.7507449999999995e-10
+ lua = -4.471944e-17
+ lub = 3.1333025e-26
+ luc = 1.0520902e-17
+ ppclm = -1.2237712e-15
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ delta = 0.01
+ pa0 = -7.365936e-14
+ nlx = 0.0
+ lpdiblc2 = 4.540744e-9
+ cdsc = 0.0
+ pk1 = -2.1256446e-15
+ pk2 = -2.3842633e-16
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ pu0 = 4.147977e-16
+ cgdo = 3.48175e-10
+ prt = 0
+ pua = 1.1289303e-23
+ pub = -3.386118e-32
+ puc = -9.620837e-24
+ cgso = 3.48175e-10
+ rsh = 6.8
+ tcj = 0.001040287
+ ua1 = 1.224e-9
+ ub1 = -4.621132e-19
+ uc1 = 6.001696e-11
+ )

.model nch_ss_13 nmos (
+ level = 49
+ drout = 0.0
+ wkt1 = 5.128653e-9
+ wkt2 = 3.532295e-9
+ tpbsw = 0.001554306
+ lint = 1e-8
+ wmax = 5.0994224e-7
+ wmin = 2.2e-7
+ cjswg = 3.507574e-10
+ lmax = 2.0001e-5
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ mjswg = 0.43879
+ lmin = 9.993989464000001e-6
+ pscbe1 = 200000030.0
+ pscbe2 = 1e-6
+ wvoff = -2.3603662000000002e-9
+ weta0 = 0
+ nqsmod = 0
+ wub1 = -4.432931e-26
+ wuc1 = -1.7086574e-17
+ tpbswg = 0.001554306
+ wvsat = 0.0
+ noimod = 2
+ hdif = 2e-7
+ wvth0 = -9.490401e-9
+ ags = 0.02
+ wute = 2.5547985e-8
+ mjsw = 0.2003879
+ cit = -9.999998e-5
+ dlc = 3e-9
+ k3b = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ cdsc = 0.0
+ cgdo = 3.48175e-10
+ cgso = 3.48175e-10
+ xpart = 1
+ jsw = 1.45e-12
+ capmod = 3
+ kt1 = -0.238767
+ lk2 = 3.6153600000000002e-9
+ kt2 = -0.03620588
+ llc = -0.039
+ cjsw = 2.142574e-10
+ lln = -1
+ a0 = 0.352982
+ a1 = 0.0
+ a2 = 0.99
+ lu0 = -4.5192000000000003e-10
+ b0 = 0.0
+ b1 = 0.0
+ pbswg = 0.6882682
+ nch = 3.9e+17
+ at = 20000.0
+ cf = 0
+ cj = 0.001050279
+ lwl = 0.0
+ lwn = 1.0
+ ef = 0.874
+ k1 = 0.5220979
+ k2 = 0.023773289
+ k3 = 0.0
+ em = 30000000.0
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ nfactor = 1.0
+ js = 3.5e-7
+ ll = 0.0
+ nlx = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ lvoff = -9.038400000000001e-10
+ u0 = 0.03352974
+ pb = 0.6882682
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ua = -5.860608e-10
+ ub = 1.7266676e-18
+ uc = 7.252202e-11
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -1.3989464e-8
+ ww = 0.0
+ xw = -9.94224e-9
+ mobmod = 1
+ beta0 = 11.59263
+ pu0 = 0.0
+ tnom = 25.0
+ leta0 = 9.680916984722288e-19
+ prt = 0
+ toxm = 4.08e-9
+ rsh = 6.8
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0006999999
+ lvth0 = 2.621136e-9
+ tcj = 0.001040287
+ ua1 = 1.224e-9
+ ub1 = -1.4270478e-18
+ uc1 = -6.39873e-11
+ pdiblcb = 0.01
+ pbsw = 0.6882682
+ pclm = 0.7999999
+ tpb = 0.001554306
+ tox = 4.14010536e-9
+ delta = 0.01
+ wa0 = 5.286186e-8
+ ute = -1.5833832
+ wk1 = -1.4938487e-9
+ wk2 = -2.6871128e-9
+ dvt0w = 0.0
+ dvt1w = 0.0
+ wln = 1.0
+ dvt2w = 0.0
+ wu0 = 9.682726e-10
+ binunit = 2
+ wua = -1.5275344e-17
+ wub = 1.2900942e-25
+ wuc = 2.9959555e-18
+ wwl = 0.0
+ wwn = 1
+ xti = 3
+ pnfactor = 0.0
+ keta = 0.002064252
+ tcjswg = 0.000645489
+ wnfactor = 0.0
+ dsub = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ tcjsw = 0.000645489
+ lnfactor = 4.5192e-8
+ voff = -0.14016372
+ version = 3.24
+ pvoff = -9.038400000000001e-16
+ ldif = 9e-8
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ eta0 = 5e-5
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 4.148964422023837e-25
+ pvag = 0.0
+ etab = -5e-5
+ vsat = 86384.63
+ wint = 3e-9
+ vth0 = 0.48181952
+ wketa = -2.9874625e-10
+ pvth0 = 2.71152e-15
+ rdsw = 170.0
+ )

.model nch_ss_14 nmos (
+ level = 49
+ la0 = -2.4964379e-7
+ pcit = 1.5653096e-18
+ pbsw = 0.6882682
+ pclm = 0.7606163
+ jsw = 1.45e-12
+ lk1 = -6.331243e-8
+ kt1 = -0.2407974
+ lk2 = 2.4414092e-8
+ kt2 = -0.03589625
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0003968183
+ pdiblcb = 0.01
+ lpscbe1 = 262.58182
+ llc = -0.039
+ lln = -1
+ lu0 = 9.442635e-9
+ lpdiblc2 = 3.0196909e-9
+ lua = -1.2876533e-16
+ lub = 7.836163e-25
+ luc = 7.064626e-17
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ pa0 = -7.427873e-14
+ nlx = 0.0
+ pk1 = 2.1894499e-14
+ pk2 = -1.0734859e-14
+ lketa = -3.0377027e-8
+ binunit = 2
+ pu0 = -1.3716021e-15
+ capmod = 3
+ prt = 0
+ pua = 1.6719826e-23
+ pub = -2.4068014e-31
+ xpart = 1
+ puc = -2.4186704e-23
+ pkt1 = -3.679308e-15
+ pkt2 = 5.879336e-16
+ rsh = 6.8
+ keta = 0.005114151
+ tcj = 0.001040287
+ ua1 = 1.224e-9
+ ub1 = -1.4513121e-18
+ uc1 = -6.991786e-11
+ pbswg = 0.6882682
+ tpb = 0.001554306
+ tox = 4.14010536e-9
+ dsub = 0.0
+ wa0 = 6.031956e-8
+ lvoff = -2.0631212000000003e-8
+ mobmod = 1
+ ute = -1.5785241
+ wk1 = -3.692092e-9
+ wk2 = -1.6093152e-9
+ wcit = -1.5715551e-13
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ wln = 1.0
+ beta0 = 11.59263
+ wu0 = 1.1059835e-9
+ wua = -1.6954039e-17
+ wub = 1.5317406e-25
+ wuc = 5.42434e-18
+ leta0 = 9.680916984722288e-19
+ wwl = 0.0
+ wwn = 1
+ lcit = 2.6386249e-10
+ xti = 3
+ voff = -0.13818312
+ lvsat = -0.005267757
+ ldif = 9e-8
+ lvth0 = 5.8899376e-8
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ pub1 = 2.1839324e-32
+ puc1 = 5.837128e-24
+ version = 3.24
+ ppclm = 7.826515e-14
+ eta0 = 5e-5
+ delta = 0.01
+ pvag = 0.0
+ etab = -5e-5
+ vsat = 86913.52
+ wint = 3e-9
+ pute = -1.7889165e-14
+ vth0 = 0.47616912
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ rdsw = 170.0
+ wkt1 = 5.498062e-9
+ wkt2 = 3.473265e-9
+ lint = 1e-8
+ wmax = 5.0994224e-7
+ wmin = 2.2e-7
+ lkt1 = 2.0222748e-8
+ lkt2 = -3.0839447e-9
+ lmax = 9.993989464000001e-6
+ tcjswg = 0.000645489
+ lmin = 1.193989464e-6
+ pketa = 4.776125e-16
+ wpclm = -7.857923e-9
+ wub1 = -4.652201e-26
+ wuc1 = -1.7672629e-17
+ tcjsw = 0.000645489
+ hdif = 2e-7
+ lub1 = 2.4167225e-25
+ a0 = 0.3780467
+ a1 = 0.0
+ a2 = 0.99
+ luc1 = 5.906839e-17
+ b0 = 0.0
+ b1 = 0.0
+ wute = 2.7344081e-8
+ mjsw = 0.2003879
+ at = 20000.0
+ pvoff = 1.8058529e-15
+ cf = 0
+ cj = 0.001050279
+ ef = 0.874
+ k1 = 0.5284545
+ k2 = 0.021685062
+ k3 = 0.0
+ em = 30000000.0
+ js = 3.5e-7
+ ll = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ u0 = 0.03253632
+ pb = 0.6882682
+ w0 = 0.0
+ rd = 0
+ lute = -4.839696e-8
+ rs = 0
+ ua = -5.731325e-10
+ ub = 1.6479914e-18
+ uc = 6.542903e-11
+ cdscb = 0.0
+ cdscd = 0.0
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -1.3989464e-8
+ ww = 0.0
+ peta0 = 4.148964422023837e-25
+ xw = -9.94224e-9
+ pvsat = 7.826533e-10
+ wketa = -3.466991e-10
+ pvth0 = 3.1711749999999997e-16
+ cdsc = 0.0
+ drout = 0.0
+ tpbsw = 0.001554306
+ cgdo = 3.48175e-10
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ cgso = 3.48175e-10
+ cjswg = 3.507574e-10
+ pscbe1 = 173636400.0
+ pscbe2 = 1e-6
+ mjswg = 0.43879
+ ags = 0.02
+ pnfactor = 0.0
+ wnfactor = 0.0
+ wvoff = -2.6324233e-9
+ cjsw = 2.142574e-10
+ cit = -0.00012649217
+ nqsmod = 0
+ dlc = 3e-9
+ tpbswg = 0.001554306
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ noimod = 2
+ k3b = 0.0
+ weta0 = 0
+ dwb = 0.0
+ dwg = 0.0
+ wvsat = -7.857954e-5
+ nfactor = 1.0
+ lpclm = 3.92261e-7
+ wvth0 = -9.25e-9
+ tnom = 25.0
+ lnfactor = 4.5192e-8
+ toxm = 4.08e-9
+ )

.model nch_ss_15 nmos (
+ level = 49
+ wub1 = -1.0574451e-25
+ wuc1 = -4.040928e-17
+ ppdiblc2 = 4.703685e-16
+ beta0 = 11.59263
+ hdif = 2e-7
+ wpdiblc2 = -4.054901e-10
+ leta0 = 3.8114280968091696e-11
+ lub1 = -8.773805e-25
+ luc1 = -7.886598e-17
+ letab = -3.811428e-11
+ lnfactor = 4.5192e-8
+ wute = 1.9757099e-8
+ lvsat = -0.0007893788
+ mjsw = 0.2003879
+ lvth0 = 1.1480395e-8
+ lute = -1.6751561e-7
+ ppclm = 4.863229e-14
+ delta = 0.01
+ lpdiblc2 = 1.4881204e-9
+ dvt0w = 0.0
+ cdsc = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ cgdo = 3.48175e-10
+ tcjswg = 0.000645489
+ cgso = 3.48175e-10
+ pketa = 3.1429577e-15
+ cjsw = 2.142574e-10
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ wpclm = 1.7687656e-8
+ tcjsw = 0.000645489
+ tnom = 25.0
+ nfactor = 1.0
+ pvoff = -2.2875942e-15
+ toxm = 4.08e-9
+ ags = 0.02
+ pcit = -9.088336e-19
+ pbsw = 0.6882682
+ pclm = 0.9728217
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 4.148964422023837e-25
+ pvsat = 1.5955267e-11
+ cit = -0.00016124053
+ wketa = -2.6444102e-9
+ pvth0 = 2.7913746499999998e-15
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0017171376
+ dlc = 3e-9
+ drout = 0.0
+ pdiblcb = 0.01
+ k3b = 0.0
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ tpbsw = 0.001554306
+ dwb = 0.0
+ dwg = 0.0
+ pscbe1 = 400000100.0
+ pscbe2 = 1e-6
+ cjswg = 3.507574e-10
+ mjswg = 0.43879
+ binunit = 2
+ pkt1 = -1.1651986e-14
+ pkt2 = -1.4582807e-15
+ keta = -0.015611105
+ nqsmod = 0
+ wvoff = 8.9641e-10
+ tpbswg = 0.001554306
+ la0 = 2.7901473e-7
+ noimod = 2
+ jsw = 1.45e-12
+ dsub = 0.0
+ lk1 = 6.936774e-8
+ kt1 = -0.2426658
+ lk2 = -2.7913247000000003e-8
+ kt2 = -0.04069558
+ llc = -0.039
+ lln = -1
+ weta0 = 0
+ lu0 = -2.1965306e-9
+ lua = 6.135559e-17
+ lub = -2.9489129e-25
+ luc = -2.7169401e-17
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ wvsat = 0.0005823669
+ wcit = 1.975718e-12
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ pa0 = 7.227613e-14
+ nlx = 0.0
+ lpclm = 1.4610272e-7
+ wvth0 = -1.138298e-8
+ pk1 = -1.920543e-14
+ pk2 = 7.699883e-15
+ lcit = 3.0417063e-10
+ voff = -0.17212312
+ pu0 = 1.0146696e-15
+ ldif = 9e-8
+ prt = 0
+ pua = -1.8126578e-24
+ pub = -2.6935e-33
+ puc = -6.78799e-24
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ pub1 = 9.053745e-32
+ puc1 = 3.221165e-23
+ eta0 = 1.7142866e-5
+ rsh = 6.8
+ pvag = 0.0
+ etab = -1.7142866e-5
+ tcj = 0.001040287
+ ua1 = 1.224e-9
+ ub1 = -4.866116e-19
+ uc1 = 4.899104e-11
+ vsat = 83052.85
+ version = 3.24
+ a0 = -0.07769345
+ wint = 3e-9
+ a1 = 0.0
+ a2 = 0.99
+ pute = -9.088265e-15
+ b0 = 0.0
+ b1 = 0.0
+ tpb = 0.001554306
+ vth0 = 0.51704752
+ tox = 4.14010536e-9
+ at = 20000.0
+ cf = 0
+ cj = 0.001050279
+ ef = 0.874
+ k1 = 0.4140751
+ k2 = 0.06679484
+ k3 = 0.0
+ rdsw = 170.0
+ wa0 = -6.602082e-8
+ em = 30000000.0
+ js = 3.5e-7
+ wkt1 = 1.2371058e-8
+ wkt2 = 5.237243e-9
+ ute = -1.4758356
+ ll = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ lint = 1e-8
+ u0 = 0.04257008
+ pb = 0.6882682
+ wk1 = 3.173889e-8
+ wk2 = -1.7501334e-8
+ w0 = 0.0
+ rd = 0
+ wmax = 5.0994224e-7
+ lketa = -6.33573e-9
+ capmod = 3
+ rs = 0
+ ua = -7.370299e-10
+ ub = 2.5777392e-18
+ uc = 1.4975288e-10
+ wln = 1.0
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -1.3989464e-8
+ ww = 0.0
+ wmin = 2.2e-7
+ wu0 = -9.511471e-10
+ xw = -9.94224e-9
+ lkt1 = 2.2390124e-8
+ wua = -9.777621e-19
+ lkt2 = 2.4832894e-9
+ wub = -5.19868e-26
+ wuc = -9.57455e-18
+ xpart = 1
+ wwl = 0.0
+ wwn = 1
+ lmax = 1.193989464e-6
+ xti = 3
+ lmin = 4.93989464e-7
+ pnfactor = 0.0
+ wnfactor = 0.0
+ pbswg = 0.6882682
+ mobmod = 1
+ lvoff = 1.8739164e-8
+ )

.model nch_ss_16 nmos (
+ level = 49
+ at = 20000.0
+ cf = 0
+ cj = 0.001050279
+ ef = 0.874
+ k1 = 0.4942783
+ k2 = 0.030748973
+ k3 = 0.0
+ em = 30000000.0
+ pketa = -1.9609824e-16
+ pkt1 = 3.435378e-15
+ pkt2 = -8.505888e-17
+ wnfactor = 0.0
+ keta = -0.030443965
+ js = 3.5e-7
+ ll = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ ags = 0.0548038
+ u0 = 0.03529582
+ pb = 0.6882682
+ w0 = 0.0
+ binunit = 2
+ rd = 0
+ rs = 0
+ ua = -6.614348e-10
+ ub = 2.1301375e-18
+ uc = 1.2526492e-10
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ wags = -1.1015922e-8
+ xl = -1.3989464e-8
+ ww = 0.0
+ dsub = 0.0
+ xw = -9.94224e-9
+ wpclm = 1.2379924e-7
+ cit = 0.00029138371
+ lags = -1.6009743e-8
+ dlc = 3e-9
+ wcit = -2.7539906e-12
+ ppdiblc2 = -1.1422951e-16
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ tcjsw = 0.000645489
+ k3b = 0.0
+ wpdiblc2 = 8.65375e-10
+ dwb = 0.0
+ dwg = 0.0
+ lnfactor = 4.5192e-8
+ lcit = 9.596344e-11
+ pvoff = -1.4007737000000002e-15
+ voff = -0.12095291999999999
+ ldif = 9e-8
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ pub1 = -3.181536e-32
+ puc1 = -1.1609298e-23
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 4.148964422023837e-25
+ eta0 = -0.00026219533
+ pvag = 0.0
+ etab = 0.0013487812
+ pvsat = 1.2452966e-11
+ la0 = 1.1871046e-7
+ vsat = 81785.22
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ wint = 3e-9
+ pute = -6.731688e-15
+ wketa = 4.614407e-9
+ lpdiblc2 = 5.562512e-9
+ pvth0 = 1.6693625999999999e-15
+ jsw = 1.45e-12
+ vth0 = 0.50482072
+ lk1 = 3.247429e-8
+ kt1 = -0.1929406
+ lk2 = -1.1332151999999999e-8
+ kt2 = -0.03937921
+ drout = 0.0
+ rdsw = 170.0
+ llc = -0.039
+ lln = -1
+ tpbsw = 0.001554306
+ pscbe1 = 400000000.0
+ pscbe2 = 1e-6
+ lu0 = 1.1496252e-9
+ version = 3.24
+ wkt1 = -2.0427562e-8
+ wkt2 = 2.2519782e-9
+ lint = 1e-8
+ lua = 2.6581833e-17
+ lub = -8.899446e-26
+ luc = -1.5904941e-17
+ nch = 3.9e+17
+ wmax = 5.0994224e-7
+ lwl = 0.0
+ lwn = 1.0
+ wmin = 2.2e-7
+ pa0 = -9.128582e-14
+ nlx = 0.0
+ cjswg = 3.507574e-10
+ lkt1 = -4.834396e-10
+ lkt2 = 1.8777602e-9
+ mjswg = 0.43879
+ pk1 = 4.587708e-15
+ pk2 = -2.4446703e-15
+ lmax = 4.93989464e-7
+ nqsmod = 0
+ tpbswg = 0.001554306
+ lmin = 1.8e-7
+ noimod = 2
+ pu0 = -1.7230291e-17
+ prt = 0
+ pua = -2.3933522e-23
+ pub = 2.5580594e-32
+ puc = 3.433529e-24
+ wvoff = -1.031461e-9
+ rsh = 6.8
+ tcj = 0.001040287
+ ua1 = 1.224e-9
+ ub1 = -3.1027764e-18
+ uc1 = -2.4653823e-10
+ weta0 = 0
+ tpb = 0.001554306
+ wub1 = 1.602399e-25
+ wuc1 = 5.485366e-17
+ tox = 4.14010536e-9
+ wvsat = 0.0005899806
+ wa0 = 2.8954867e-7
+ hdif = 2e-7
+ lpclm = 7.125815e-8
+ wvth0 = -8.94382e-9
+ ute = -1.9466008
+ wk1 = -1.9985334e-8
+ wk2 = 4.552045e-9
+ lub1 = 3.260553e-25
+ luc1 = 5.707747e-17
+ wute = 1.4634106e-8
+ wln = 1.0
+ mjsw = 0.2003879
+ wu0 = 1.2921135e-9
+ wua = 4.711108e-17
+ wub = -1.1345223e-25
+ wuc = -3.179524e-17
+ wwl = 0.0
+ wwn = 1
+ xti = 3
+ lute = 4.90364e-8
+ cdsc = 0.0
+ capmod = 3
+ cgdo = 3.48175e-10
+ lketa = 4.87385e-10
+ cgso = 3.48175e-10
+ xpart = 1
+ mobmod = 1
+ cjsw = 2.142574e-10
+ pbswg = 0.6882682
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ lvoff = -4.7991109999999995e-9
+ beta0 = 11.59263
+ leta0 = 1.666098409680917e-10
+ tnom = 25.0
+ letab = -6.664392e-10
+ lvsat = -0.00020626588
+ pags = 5.067323e-15
+ lvth0 = 1.7104719e-8
+ toxm = 4.08e-9
+ nfactor = 1.0
+ pcit = 1.266836e-18
+ ppclm = -1.7902992e-16
+ pbsw = 0.6882682
+ pclm = 1.1355271
+ delta = 0.01
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ tcjswg = 0.000645489
+ pdiblc1 = 1e-6
+ pdiblc2 = -0.007140237
+ pdiblcb = 0.01
+ a0 = 0.270794
+ a1 = 0.0
+ a2 = 0.99
+ b0 = 0.0
+ b1 = 0.0
+ pnfactor = 0.0
+ )

.model nch_ff_1 nmos (
+ level = 49
+ cjsw = 1.93852e-10
+ drout = 0.0
+ tpbsw = 0.001554306
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ cjswg = 3.17352e-10
+ pnfactor = 0.0
+ mjswg = 0.43879
+ wnfactor = 0.0
+ tnom = 25.0
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ wvoff = 6.32688e-10
+ pscbe1 = 200000030.0
+ pscbe2 = 1e-6
+ toxm = 4.08e-9
+ version = 3.24
+ pbsw = 0.6882682
+ pclm = 0.8000001
+ weta0 = 0
+ wvsat = 0.0
+ nqsmod = 0
+ lnfactor = -4.5192e-8
+ tpbswg = 0.001554306
+ wvth0 = -5.9653440000000004e-9
+ noimod = 2
+ ags = 0.02
+ keta = 0.009263485
+ cit = -0.00010000001
+ a0 = 0.3700794
+ a1 = 0.0
+ a2 = 0.99
+ b0 = 0.0
+ b1 = 0.0
+ dlc = 3e-9
+ dsub = 0.0
+ k3b = 0.0
+ at = 20000.0
+ cf = 0
+ cj = 0.0009502527
+ ef = 0.874
+ k1 = 0.5142301
+ k2 = 0.007567123999999999
+ k3 = 0.0
+ em = 30000000.0
+ dwb = 0.0
+ dwg = 0.0
+ js = 3.5e-7
+ ll = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ u0 = 0.04401107
+ pb = 0.6882682
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ dvt0 = 0.0
+ ua = -6.12274e-10
+ dvt1 = 0.0
+ ub = 2.3135539e-18
+ xpart = 1
+ dvt2 = 0.0
+ uc = 1.0876087e-10
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -2.6010536e-8
+ ww = 0.0
+ xw = 9.94224e-9
+ voff = -0.13786648
+ capmod = 3
+ ldif = 9e-8
+ pbswg = 0.6882682
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ jsw = 1.45e-12
+ kt1 = -0.2240464
+ lk2 = -3.6153600000000002e-9
+ kt2 = -0.030266136
+ lvoff = 9.038400000000001e-10
+ eta0 = 5e-5
+ llc = -0.039
+ lln = -1
+ pvag = 0.0
+ etab = -5e-5
+ lu0 = 4.5192000000000003e-10
+ vsat = 93615.37
+ beta0 = 11.59263
+ nch = 3.9e+17
+ wint = 3e-9
+ lwl = 0.0
+ lwn = 1.0
+ vth0 = 0.41802738
+ leta0 = 3.163440009680917e-10
+ mobmod = 1
+ nlx = 0.0
+ rdsw = 170.0
+ lint = 1e-8
+ wmax = 0.000900001
+ lvth0 = -2.621136e-9
+ pu0 = 0.0
+ wmin = 9.99005776e-6
+ prt = 0
+ lmax = 2.0001e-5
+ delta = 0.01
+ lmin = 1.0006010536e-5
+ rsh = 6.8
+ tcj = 0.001040287
+ ua1 = 1.224e-9
+ ub1 = -1.1209314e-18
+ uc1 = 1.1643822e-11
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ tpb = 0.001554306
+ tox = 4.01989464e-9
+ ute = -1.5799998
+ wln = 1.0
+ wu0 = 0.0
+ nfactor = 1.0
+ hdif = 2e-7
+ wwl = 0.0
+ wwn = 1
+ xti = 3
+ mjsw = 0.2003879
+ tcjswg = 0.000645489
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0006999999
+ pdiblcb = 0.01
+ tcjsw = 0.000645489
+ cdsc = 0.0
+ pvoff = 9.038400000000001e-16
+ cgdo = 3.84825e-10
+ binunit = 2
+ cgso = 3.84825e-10
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 1.3557600041489644e-16
+ pvth0 = -2.71152e-15
+ )

.model nch_ff_2 nmos (
+ level = 49
+ wmax = 0.000900001
+ wmin = 9.99005776e-6
+ lkt2 = -4.553491e-12
+ lmax = 1.0006010536e-5
+ lmin = 1.2060105359999999e-6
+ la0 = -3.496093e-7
+ jsw = 1.45e-12
+ kt1 = -0.2240468
+ lk1 = 1.4908844e-8
+ kt2 = -0.03026568
+ lk2 = -1.472874e-8
+ llc = -0.039
+ lln = -1
+ lketa = -4.320781e-8
+ lu0 = 3.743729e-9
+ lua = -4.643216e-16
+ lub = 7.375677e-25
+ luc = 3.898355e-17
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ xpart = 1
+ pnfactor = 0.0
+ nlx = 0.0
+ hdif = 2e-7
+ wnfactor = 0.0
+ capmod = 3
+ lub1 = 4.527317e-28
+ luc1 = 7.827772e-20
+ nfactor = 1.0
+ pu0 = 0.0
+ mjsw = 0.2003879
+ prt = 0
+ pbswg = 0.6882682
+ lute = -5.743953e-11
+ lvoff = -9.567488e-9
+ rsh = 6.8
+ tcj = 0.001040287
+ ua1 = 1.224e-9
+ ub1 = -1.1209769e-18
+ uc1 = 1.1635963e-11
+ mobmod = 1
+ beta0 = 11.59263
+ tpb = 0.001554306
+ tox = 4.01989464e-9
+ lnfactor = -4.5192e-8
+ leta0 = 3.163440009680917e-10
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0003968181
+ cdsc = 0.0
+ pdiblcb = 0.01
+ lpscbe1 = 262.58185
+ ute = -1.5799941
+ lvsat = -0.006562638
+ cgdo = 3.84825e-10
+ wln = 1.0
+ lvth0 = 5.799173400000001e-8
+ wu0 = 0.0
+ wwl = 0.0
+ wwn = 1
+ cgso = 3.84825e-10
+ xti = 3
+ delta = 0.01
+ lpdiblc2 = 3.0196912e-9
+ binunit = 2
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ cjsw = 1.93852e-10
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ tnom = 25.0
+ tcjswg = 0.000645489
+ a0 = 0.4051808
+ a1 = 0.0
+ a2 = 0.99
+ b0 = 0.0
+ b1 = 0.0
+ at = 20000.0
+ cf = 0
+ cj = 0.0009502527
+ ef = 0.874
+ k1 = 0.5127332
+ k2 = 0.008682927
+ k3 = 0.0
+ em = 30000000.0
+ toxm = 4.08e-9
+ js = 3.5e-7
+ ll = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ u0 = 0.04368057
+ pb = 0.6882682
+ w0 = 0.0
+ pbsw = 0.6882682
+ rd = 0
+ pclm = 0.7736172
+ rs = 0
+ ua = -5.656554e-10
+ ub = 2.2395009e-18
+ uc = 1.0484686e-10
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -2.6010536e-8
+ ww = 0.0
+ xw = 9.94224e-9
+ tcjsw = 0.000645489
+ version = 3.24
+ pvoff = 9.038400000000001e-16
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 1.3557600041489644e-16
+ pvth0 = -2.71152e-15
+ keta = 0.013601619
+ drout = 0.0
+ tpbsw = 0.001554306
+ dsub = 0.0
+ cjswg = 3.17352e-10
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ mjswg = 0.43879
+ pscbe1 = 173636400.0
+ pscbe2 = 1e-6
+ lcit = 2.6652053e-10
+ wvoff = 6.32688e-10
+ voff = -0.13681518
+ ldif = 9e-8
+ ags = 0.02
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ weta0 = 0
+ nqsmod = 0
+ eta0 = 5e-5
+ tpbswg = 0.001554306
+ pvag = 0.0
+ etab = -5e-5
+ cit = -0.00012675911
+ noimod = 2
+ wvsat = 0.0
+ vsat = 94274.27
+ wint = 3e-9
+ dlc = 3e-9
+ lpclm = 2.6277317e-7
+ wvth0 = -5.9653440000000004e-9
+ vth0 = 0.41194178
+ k3b = 0.0
+ rdsw = 170.0
+ dwb = 0.0
+ dwg = 0.0
+ lint = 1e-8
+ )

.model nch_ff_3 nmos (
+ level = 49
+ beta0 = 11.59263
+ leta0 = 3.544582809680917e-10
+ letab = -3.811428e-11
+ lvsat = -0.0007622857
+ version = 3.24
+ lvth0 = 1.3216209999999997e-9
+ delta = 0.01
+ keta = -0.015927497
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ dsub = 0.0
+ pnfactor = 0.0
+ lags = -3.044698e-8
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ tcjswg = 0.000645489
+ wnfactor = 0.0
+ lcit = 3.0262734e-10
+ voff = -0.15940708
+ ldif = 9e-8
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ eta0 = 1.7142866e-5
+ pvag = 0.0
+ etab = -1.7142866e-5
+ vsat = 89273.96
+ tcjsw = 0.000645489
+ lnfactor = -4.5192e-8
+ wint = 3e-9
+ vth0 = 0.46079528
+ rdsw = 170.0
+ pvoff = 9.038400000000001e-16
+ lint = 1e-8
+ wmax = 0.000900001
+ wmin = 9.99005776e-6
+ cdscb = 0.0
+ cdscd = 0.0
+ lkt1 = 5.782678e-9
+ lkt2 = 1.5570838e-9
+ peta0 = 1.3557600041489644e-16
+ lmax = 1.2060105359999999e-6
+ lpdiblc2 = 1.525682e-9
+ lmin = 5.06010536e-7
+ pvth0 = -2.71152e-15
+ ags = 0.0462474
+ drout = 0.0
+ tpbsw = 0.001554306
+ cit = -0.00015788565
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ dlc = 3e-9
+ cjswg = 3.17352e-10
+ k3b = 0.0
+ pscbe1 = 400000100.0
+ pscbe2 = 1e-6
+ mjswg = 0.43879
+ dwb = 0.0
+ dwg = 0.0
+ hdif = 2e-7
+ lua1 = -3.0446746e-18
+ lub1 = -1.2004175e-24
+ luc1 = -6.517273e-17
+ wvoff = 6.32688e-10
+ mjsw = 0.2003879
+ nqsmod = 0
+ tpbswg = 0.001554306
+ noimod = 2
+ nfactor = 1.0
+ lute = -2.6630502e-7
+ weta0 = 0
+ la0 = 4.581426e-7
+ wvsat = 0.0
+ jsw = 1.45e-12
+ kt1 = -0.2290285
+ lk1 = -7.214246e-9
+ kt2 = -0.031611919
+ lk2 = -1.9122090000000005e-9
+ lpclm = 1.5245718e-7
+ wvth0 = -5.9653440000000004e-9
+ a0 = -0.2911571
+ a1 = 0.0
+ a2 = 0.99
+ b0 = 0.0
+ b1 = 0.0
+ llc = -0.039
+ cdsc = 0.0
+ lln = -1
+ lu0 = 1.4925279e-9
+ at = 20000.0
+ cf = 0
+ cj = 0.0009502527
+ ef = 0.874
+ k1 = 0.5318048
+ k2 = -0.002365807
+ k3 = 0.0
+ em = 30000000.0
+ lua = 7.982966e-17
+ lub = -1.5630905e-25
+ luc = -9.669895e-18
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ js = 3.5e-7
+ cgdo = 3.84825e-10
+ ll = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0016847569
+ u0 = 0.04562126
+ pb = 0.6882682
+ w0 = 0.0
+ rd = 0
+ nlx = 0.0
+ rs = 0
+ pdiblcb = 0.01
+ ua = -1.0347512e-9
+ ub = 3.0100842e-18
+ uc = 1.4678947e-10
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -2.6010536e-8
+ ww = 0.0
+ xw = 9.94224e-9
+ cgso = 3.84825e-10
+ pu0 = 0.0
+ prt = 0
+ cjsw = 1.93852e-10
+ binunit = 2
+ rsh = 6.8
+ tcj = 0.001040287
+ ua1 = 1.2266247e-9
+ ub1 = -8.574386e-20
+ uc1 = 6.788683e-11
+ lketa = -8.954029e-9
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ tpb = 0.001554306
+ tox = 4.01989464e-9
+ capmod = 3
+ xpart = 1
+ ute = -1.3504703
+ tnom = 25.0
+ wln = 1.0
+ wu0 = 0.0
+ pbswg = 0.6882682
+ wwl = 0.0
+ wwn = 1
+ xti = 3
+ toxm = 4.08e-9
+ mobmod = 1
+ lvoff = 1.6639098000000002e-8
+ pbsw = 0.6882682
+ pclm = 0.8687172
+ )

.model nch_ff_4 nmos (
+ level = 49
+ lua1 = 8.039099e-19
+ lub1 = 3.824101e-25
+ luc1 = 2.9606131e-17
+ mjsw = 0.2003879
+ lute = 7.030476e-8
+ ags = -0.019916179
+ tcjsw = 0.000645489
+ nfactor = 1.0
+ cdsc = 0.0
+ cit = 0.000271889
+ pvoff = 9.038400000000001e-16
+ dlc = 3e-9
+ cgdo = 3.84825e-10
+ k3b = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cgso = 3.84825e-10
+ peta0 = 1.3557600041489644e-16
+ pdiblc1 = 1e-6
+ pdiblc2 = -0.00593541
+ pdiblcb = 0.01
+ pvth0 = -2.71152e-15
+ drout = 0.0
+ alpha0 = 0.0
+ cjsw = 1.93852e-10
+ alpha1 = 0.448150714
+ tpbsw = 0.001554306
+ la0 = 7.545271e-8
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ pscbe1 = 400000000.0
+ pscbe2 = 1e-6
+ binunit = 2
+ jsw = 1.45e-12
+ kt1 = -0.22715
+ lk1 = 4.899558e-8
+ kt2 = -0.029537767
+ lk2 = -2.6956696000000003e-8
+ cjswg = 3.17352e-10
+ pnfactor = 0.0
+ llc = -0.039
+ lln = -1
+ mjswg = 0.43879
+ lu0 = 1.7037189e-9
+ wnfactor = 0.0
+ lua = -1.0530929e-18
+ lub = 5.559478e-27
+ luc = 4.133919e-18
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ tnom = 25.0
+ nqsmod = 0
+ tpbswg = 0.001554306
+ wvoff = 6.32688e-10
+ nlx = 0.0
+ noimod = 2
+ toxm = 4.08e-9
+ pu0 = 0.0
+ weta0 = 0
+ pbsw = 0.6882682
+ pclm = 1.1076791
+ prt = 0
+ wvsat = 0.0
+ lnfactor = -4.5192e-8
+ lpclm = 4.253467e-8
+ wvth0 = -5.9653440000000004e-9
+ rsh = 6.8
+ tcj = 0.001040287
+ ua1 = 1.2182583e-9
+ ub1 = -3.526674e-18
+ uc1 = -1.381542e-10
+ tpb = 0.001554306
+ tox = 4.01989464e-9
+ ute = -2.0822308
+ version = 3.24
+ wln = 1.0
+ wu0 = 0.0
+ lpdiblc2 = 5.030957e-9
+ wwl = 0.0
+ wwn = 1
+ xti = 3
+ keta = -0.04182327
+ capmod = 3
+ dsub = 0.0
+ lketa = 2.9580252e-9
+ xpart = 1
+ lags = -1.1735286e-11
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ lcit = 1.0493098e-10
+ voff = -0.12183828000000001
+ pbswg = 0.6882682
+ mobmod = 1
+ ldif = 9e-8
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ lvoff = -6.425217999999999e-10
+ eta0 = -0.0002937502
+ pvag = 0.0
+ etab = 0.0013875004
+ beta0 = 11.59263
+ vsat = 88054.32
+ wint = 3e-9
+ leta0 = 4.974690609680917e-10
+ vth0 = 0.45670238
+ letab = -6.842502e-10
+ rdsw = 170.0
+ lvsat = -0.00020125005
+ lint = 1e-8
+ lvth0 = 3.2043650000000002e-9
+ wmax = 0.000900001
+ wmin = 9.99005776e-6
+ lkt1 = 4.918561e-9
+ lkt2 = 6.029743e-10
+ delta = 0.01
+ lmax = 5.06010536e-7
+ a0 = 0.5407774
+ a1 = 0.0
+ a2 = 0.99
+ b0 = 0.0
+ b1 = 0.0
+ lmin = 1.8e-7
+ at = 20000.0
+ cf = 0
+ cj = 0.0009502527
+ ef = 0.874
+ k1 = 0.4096095
+ k2 = 0.05207874
+ k3 = 0.0
+ em = 30000000.0
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ js = 3.5e-7
+ ll = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ u0 = 0.04516215
+ pb = 0.6882682
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ua = -8.589192e-10
+ ub = 2.6581962e-18
+ uc = 1.1678118e-10
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -2.6010536e-8
+ ww = 0.0
+ xw = 9.94224e-9
+ tcjswg = 0.000645489
+ hdif = 2e-7
+ )

.model nch_ff_5 nmos (
+ level = 49
+ pu0 = 0.0
+ pscbe1 = 200000030.0
+ pscbe2 = 1e-6
+ tpbsw = 0.001554306
+ prt = 0
+ dsub = 0.0
+ cjswg = 3.17352e-10
+ rsh = 6.8
+ tcj = 0.001040287
+ ua1 = 1.224e-9
+ ub1 = -1.0684574e-18
+ a0 = 0.3702259
+ a1 = 0.0
+ a2 = 0.99
+ uc1 = 2.4230474e-11
+ b0 = 0.0
+ b1 = 0.0
+ mjswg = 0.43879
+ nqsmod = 0
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ tpbswg = 0.001554306
+ at = 20000.0
+ cf = 0
+ cj = 0.0009502527
+ ef = 0.874
+ k1 = 0.5102321
+ k2 = 0.008860774000000002
+ k3 = 0.0
+ tpb = 0.001554306
+ noimod = 2
+ em = 30000000.0
+ tox = 4.01989464e-9
+ js = 3.5e-7
+ wa0 = -1.4643313e-9
+ ll = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ wvoff = 1.5234104e-9
+ u0 = 0.04484358
+ pb = 0.6882682
+ w0 = 0.0
+ rd = 0
+ ute = -1.5803809
+ rs = 0
+ ua = -5.885942e-10
+ ub = 2.3329335e-18
+ uc = 1.1057788e-10
+ voff = -0.13795558
+ wk1 = 3.995606e-8
+ wk2 = -1.2928737e-8
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -2.6010536e-8
+ ww = 0.0
+ ldif = 9e-8
+ xw = 9.94224e-9
+ wln = 1.0
+ wu0 = -8.320099e-9
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ puc1 = -1.4905616e-28
+ weta0 = 0
+ wua = -2.3665659e-16
+ wub = -1.936796e-25
+ wuc = -1.815927e-17
+ wwl = 0.0
+ wwn = 1
+ eta0 = 5e-5
+ xti = 3
+ wvsat = 0.0
+ pvag = 0.0
+ etab = -5e-5
+ vsat = 93615.37
+ wvth0 = -5.2777326e-9
+ wint = 3e-9
+ vth0 = 0.41795858
+ rdsw = 170.0
+ wkt1 = -8.215166e-9
+ wkt2 = 1.6245854e-9
+ lint = 1e-8
+ wmax = 9.99005776e-6
+ wmin = 1.19005776e-6
+ lmax = 2.0001e-5
+ lmin = 1.0006010536e-5
+ capmod = 3
+ xpart = 1
+ wub1 = -5.244247e-25
+ pnfactor = 0.0
+ wuc1 = -1.257911e-16
+ wnfactor = 0.0
+ hdif = 2e-7
+ mobmod = 1
+ wute = 3.808433e-9
+ pbswg = 0.6882682
+ mjsw = 0.2003879
+ lvoff = 9.038400000000001e-10
+ beta0 = 11.59263
+ lnfactor = -4.5192e-8
+ leta0 = 3.163440009680917e-10
+ cdsc = 0.0
+ nfactor = 1.0
+ lvth0 = -2.621136e-9
+ cgdo = 3.84825e-10
+ cgso = 3.84825e-10
+ delta = 0.01
+ dvt0w = 0.0
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0006999999
+ dvt1w = 0.0
+ dvt2w = 0.0
+ pdiblcb = 0.01
+ cjsw = 1.93852e-10
+ tcjswg = 0.000645489
+ ags = 0.02
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ cit = -0.00010000001
+ binunit = 2
+ dlc = 3e-9
+ tnom = 25.0
+ k3b = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ toxm = 4.08e-9
+ pbsw = 0.6882682
+ pclm = 0.8000001
+ tcjsw = 0.000645489
+ pvoff = 9.038400000000001e-16
+ jsw = 1.45e-12
+ kt1 = -0.2232244
+ kt2 = -0.030428693
+ lk2 = -3.6153600000000002e-9
+ llc = -0.039
+ lln = -1
+ lu0 = 4.5192000000000003e-10
+ cdscb = 0.0
+ cdscd = 0.0
+ nch = 3.9e+17
+ peta0 = 1.3557600041489644e-16
+ lwl = 0.0
+ lwn = 1.0
+ nlx = 0.0
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ version = 3.24
+ wketa = -1.0935369e-8
+ pvth0 = -2.71152e-15
+ keta = 0.010357677
+ drout = 0.0
+ )

.model nch_ff_6 nmos (
+ level = 49
+ nfactor = 1.0
+ cgso = 3.84825e-10
+ capmod = 3
+ cjsw = 1.93852e-10
+ lketa = -4.518989e-8
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0003968181
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ pdiblcb = 0.01
+ lpscbe1 = 262.58185
+ xpart = 1
+ mobmod = 1
+ tnom = 25.0
+ pbswg = 0.6882682
+ binunit = 2
+ toxm = 4.08e-9
+ lvoff = -9.902212e-9
+ a0 = 0.40626
+ a1 = 0.0
+ a2 = 0.99
+ b0 = 0.0
+ b1 = 0.0
+ pbsw = 0.6882682
+ pclm = 0.7755287
+ at = 20000.0
+ cf = 0
+ cj = 0.0009502527
+ ef = 0.874
+ k1 = 0.508509
+ beta0 = 11.59263
+ k2 = 0.01007951
+ k3 = 0.0
+ em = 30000000.0
+ js = 3.5e-7
+ ll = 0.0
+ leta0 = 3.163440009680917e-10
+ mj = 0.3595262
+ lw = 0.0
+ u0 = 0.04453795
+ pb = 0.6882682
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ags = 0.02
+ ua = -5.377125e-10
+ ub = 2.2537915e-18
+ uc = 1.0657759e-10
+ lvsat = -0.006753025
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -2.6010536e-8
+ ww = 0.0
+ xw = 9.94224e-9
+ lvth0 = 5.8084954e-8
+ cit = -0.00012675911
+ ppclm = 1.9027247e-13
+ delta = 0.01
+ dlc = 3e-9
+ k3b = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ tcjswg = 0.000645489
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ pkt1 = 4.710912e-15
+ pkt2 = -4.130377e-15
+ keta = 0.014894814
+ version = 3.24
+ dsub = 0.0
+ pnfactor = 0.0
+ la0 = -3.588995e-7
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ wnfactor = 0.0
+ jsw = 1.45e-12
+ lk1 = 1.7161611e-8
+ kt1 = -0.2231775
+ lk2 = -1.5753972e-8
+ kt2 = -0.030469729
+ pketa = 1.9809019e-14
+ llc = -0.039
+ lln = -1
+ lu0 = 3.4960111999999998e-9
+ lcit = 2.6652053e-10
+ voff = -0.13687068
+ lua = -5.067804e-16
+ lub = 7.882536e-25
+ luc = 3.984287e-17
+ nch = 3.9e+17
+ ldif = 9e-8
+ lwl = 0.0
+ lwn = 1.0
+ wpclm = -1.9103656e-8
+ kt1l = 0.0
+ pa0 = 9.284546e-14
+ prwb = 0.0
+ prwg = 0.0
+ pub1 = 4.176128e-31
+ nlx = 0.0
+ puc1 = 7.417578e-23
+ eta0 = 5e-5
+ pk1 = -2.2514154e-14
+ pk2 = 1.0246181e-14
+ pvag = 0.0
+ etab = -5e-5
+ tcjsw = 0.000645489
+ pu0 = 2.4756895e-15
+ vsat = 94293.38
+ lnfactor = -4.5192e-8
+ wint = 3e-9
+ pute = -5.708167e-14
+ prt = 0
+ pua = 4.243342e-22
+ pub = -5.065558e-31
+ puc = -8.588134e-24
+ vth0 = 0.41186368
+ rdsw = 170.0
+ pvoff = 4.249081000000001e-15
+ wkt1 = -8.688151e-9
+ wkt2 = 2.0392819e-9
+ rsh = 6.8
+ lint = 1e-8
+ tcj = 0.001040287
+ ua1 = 1.224e-9
+ ub1 = -1.0643074e-18
+ uc1 = 2.4967807e-11
+ wmax = 9.99005776e-6
+ wmin = 1.19005776e-6
+ cdscb = 0.0
+ cdscd = 0.0
+ tpb = 0.001554306
+ peta0 = 1.3557600041489644e-16
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ tox = 4.01989464e-9
+ lkt1 = -4.674615e-10
+ lkt2 = 4.087321e-10
+ wa0 = -1.0786144e-8
+ lpdiblc2 = 3.0196912e-9
+ lmax = 1.0006010536e-5
+ pvsat = 1.9027204e-9
+ ute = -1.5809486
+ pscbe1 = 173636400.0
+ pscbe2 = 1e-6
+ wk1 = 4.221652e-8
+ wk2 = -1.3957471e-8
+ lmin = 1.2060105359999999e-6
+ wketa = -1.292423e-8
+ pvth0 = -3.6432075e-15
+ wln = 1.0
+ drout = 0.0
+ wu0 = -8.568663e-9
+ tpbsw = 0.001554306
+ wua = -2.7926046e-16
+ wub = -1.4282058e-25
+ wuc = -1.7297008e-17
+ wwl = 0.0
+ wwn = 1
+ xti = 3
+ nqsmod = 0
+ tpbswg = 0.001554306
+ cjswg = 3.17352e-10
+ noimod = 2
+ wub1 = -5.663537e-25
+ wuc1 = -1.3323848e-16
+ mjswg = 0.43879
+ hdif = 2e-7
+ wvoff = 1.1875419e-9
+ lub1 = -4.133362e-26
+ luc1 = -7.343755e-18
+ wute = 9.539526e-9
+ mjsw = 0.2003879
+ weta0 = 0
+ lute = 5.654154e-9
+ wvsat = -0.00019104627
+ lpclm = 2.4373449e-7
+ wvth0 = -5.184193800000001e-9
+ cdsc = 0.0
+ cgdo = 3.84825e-10
+ )

.model nch_ff_7 nmos (
+ level = 49
+ beta0 = 11.59263
+ pvag = 0.0
+ etab = -1.7142869e-5
+ vsat = 89128.95
+ leta0 = 3.544582809680917e-10
+ wint = 3e-9
+ pute = 4.357466e-13
+ letab = -3.811428e-11
+ vth0 = 0.46146618
+ lvsat = -0.0007622865
+ rdsw = 170.0
+ lvth0 = 5.459959999999999e-10
+ wkt1 = -3.681822e-9
+ wkt2 = -1.3190541e-9
+ lint = 1e-8
+ wmax = 9.99005776e-6
+ la0 = 4.645035e-7
+ ppclm = 7.258032e-15
+ wmin = 1.19005776e-6
+ jsw = 1.45e-12
+ lk1 = -1.1179709e-8
+ kt1 = -0.2286601
+ lk2 = -1.8429500000000034e-10
+ kt2 = -0.031479932
+ delta = 0.01
+ tcjswg = 0.000645489
+ lkt1 = 5.892387e-9
+ lkt2 = 1.5805686e-9
+ llc = -0.039
+ lln = -1
+ lmax = 1.2060105359999999e-6
+ lu0 = 1.4123913000000001e-9
+ lmin = 5.06010536e-7
+ lua = 6.148926e-17
+ lub = -1.2783527e-25
+ luc = -6.505068e-18
+ nch = 3.9e+17
+ dvt0w = 0.0
+ lwl = 0.0
+ lwn = 1.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ pa0 = -6.357063e-14
+ nlx = 0.0
+ pk1 = 3.963084e-14
+ pk2 = -1.7268767e-14
+ pu0 = 8.008865e-16
+ prt = 0
+ pua = 1.8329395e-22
+ pub = -2.8456703e-31
+ puc = -3.16293e-23
+ wua1 = -3.55913e-18
+ wub1 = -1.6132161e-24
+ wuc1 = -1.8047248e-16
+ hdif = 2e-7
+ rsh = 6.8
+ pketa = 9.843987e-15
+ tcj = 0.001040287
+ ua1 = 1.2269809e-9
+ ub1 = 7.567455e-20
+ lua1 = -3.457781e-18
+ uc1 = 8.594492e-11
+ lub1 = -1.3637128e-24
+ luc1 = -7.807721e-17
+ wute = -4.153124e-7
+ mjsw = 0.2003879
+ tpb = 0.001554306
+ tox = 4.01989464e-9
+ wa0 = 1.2405528e-7
+ wpclm = 1.3866737e-7
+ ute = -1.3089141
+ lute = -3.0990586e-7
+ wk1 = -1.1356744e-8
+ wk2 = 9.762311e-9
+ wln = 1.0
+ tcjsw = 0.000645489
+ wu0 = -7.124867e-9
+ wua = -7.146715e-17
+ wub = -3.341902e-25
+ wuc = 2.5660584e-18
+ wwl = 0.0
+ wwn = 1
+ xti = 3
+ cdsc = 0.0
+ pvoff = -2.109974e-15
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ cgdo = 3.84825e-10
+ a0 = -0.3035701
+ a1 = 0.0
+ a2 = 0.99
+ b0 = 0.0
+ b1 = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 1.3557600041489644e-16
+ at = 20000.0
+ cf = 0
+ cj = 0.0009502527
+ pscbe1 = 400000100.0
+ pscbe2 = 1e-6
+ ef = 0.874
+ k1 = 0.5329412
+ k2 = -0.0033426250000000005
+ k3 = 0.0
+ em = 30000000.0
+ cgso = 3.84825e-10
+ js = 3.5e-7
+ ll = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ u0 = 0.04633417
+ pb = 0.6882682
+ nfactor = 1.0
+ w0 = 0.0
+ rd = 0
+ wketa = -4.333682e-9
+ rs = 0
+ ua = -1.0276002e-9
+ ub = 3.0435232e-18
+ uc = 1.4653272e-10
+ pvth0 = 5.040078e-15
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -2.6010536e-8
+ ww = 0.0
+ xw = 9.94224e-9
+ drout = 0.0
+ tpbsw = 0.001554306
+ nqsmod = 0
+ cjsw = 1.93852e-10
+ tpbswg = 0.001554306
+ noimod = 2
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ cjswg = 3.17352e-10
+ pnfactor = 0.0
+ mjswg = 0.43879
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0017737894
+ pdiblcb = 0.01
+ wnfactor = 0.0
+ tnom = 25.0
+ wvoff = 6.6694859999999994e-9
+ pags = 4.128623e-14
+ toxm = 4.08e-9
+ weta0 = 0
+ ppdiblc2 = 1.0321563e-15
+ binunit = 2
+ pbsw = 0.6882682
+ pclm = 0.8548421
+ wvsat = 0.0014492224
+ wpdiblc2 = -8.897895e-10
+ lpclm = 1.5173094e-7
+ wvth0 = -1.266978e-8
+ lnfactor = -4.5192e-8
+ capmod = 3
+ lpdiblc2 = 1.4224044e-9
+ pkt1 = -1.0964308e-15
+ pkt2 = -2.3470743e-16
+ keta = -0.01549387
+ lketa = -9.939018e-9
+ mobmod = 1
+ wags = -3.559157e-8
+ dsub = 0.0
+ version = 3.24
+ xpart = 1
+ ags = 0.04980868
+ lags = -3.457808e-8
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ cit = -0.00015788565
+ pbswg = 0.6882682
+ lcit = 3.0262734e-10
+ voff = -0.16001108
+ ldif = 9e-8
+ dlc = 3e-9
+ k3b = 0.0
+ kt1l = 0.0
+ lvoff = 1.6940662e-8
+ pua1 = 4.128591e-24
+ prwb = 0.0
+ prwg = 0.0
+ pub1 = 1.6319734e-30
+ puc1 = 1.2896722e-22
+ dwb = 0.0
+ dwg = 0.0
+ eta0 = 1.7142869e-5
+ )

.model nch_ff_8 nmos (
+ level = 49
+ pketa = -2.7027957e-15
+ tnom = 25.0
+ pdiblc1 = 1e-6
+ pdiblc2 = -0.006119013
+ pdiblcb = 0.01
+ pags = -1.0838496e-14
+ toxm = 4.08e-9
+ wpclm = 6.656068e-8
+ pcit = 1.4220811e-17
+ pbsw = 0.6882682
+ pclm = 1.1010191
+ tcjsw = 0.000645489
+ binunit = 2
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ pvoff = -7.157499999999998e-17
+ pscbe1 = 400000000.0
+ pscbe2 = 1e-6
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 1.3419387861489644e-16
+ petab = 1.6959704e-18
+ pvsat = 1.5350395e-12
+ wketa = 2.2941933e-8
+ nqsmod = 0
+ pvth0 = 1.797418e-15
+ tpbswg = 0.001554306
+ drout = 0.0
+ noimod = 2
+ pkt1 = -1.7512235e-15
+ pkt2 = 7.382567e-17
+ keta = -0.04411884
+ tpbsw = 0.001554306
+ wags = 7.772305e-8
+ dsub = 0.0
+ cjswg = 3.17352e-10
+ mjswg = 0.43879
+ lags = 1.0727657e-9
+ wcit = -3.0914837e-11
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ version = 3.24
+ wvoff = 2.2381844e-9
+ lcit = 1.0350804e-10
+ voff = -0.12199898
+ ldif = 9e-8
+ weta0 = 3.0046217e-12
+ kt1l = 0.0
+ pua1 = -1.0901051e-24
+ prwb = 0.0
+ prwg = 0.0
+ pub1 = -4.238914e-31
+ puc1 = -2.7204607e-23
+ wetab = -3.686654e-12
+ wvsat = 0.0014459029
+ eta0 = -0.00029405078
+ pvag = 0.0
+ etab = 0.0013878694
+ lpclm = 3.848953e-8
+ wvth0 = -5.6205204000000005e-9
+ vsat = 87909.64
+ wint = 3e-9
+ pute = -1.178615e-13
+ vth0 = 0.45666788
+ rdsw = 170.0
+ capmod = 3
+ wkt1 = -2.2583577e-9
+ wkt2 = -1.9897783e-9
+ lint = 1e-8
+ ags = -0.027693154
+ wmax = 9.99005776e-6
+ wmin = 1.19005776e-6
+ lkt1 = 5.093789e-9
+ lkt2 = 5.955873e-10
+ lmax = 5.06010536e-7
+ cit = 0.00027498236
+ lmin = 1.8e-7
+ dlc = 3e-9
+ mobmod = 1
+ k3b = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ a0 = 0.5262308
+ a1 = 0.0
+ a2 = 0.99
+ lketa = 3.228467e-9
+ b0 = 0.0
+ b1 = 0.0
+ at = 20000.0
+ cf = 0
+ cj = 0.0009502527
+ ef = 0.874
+ k1 = 0.4007356
+ k2 = 0.055957879999999995
+ k3 = 0.0
+ em = 30000000.0
+ xpart = 1
+ js = 3.5e-7
+ ll = 0.0
+ pnfactor = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ u0 = 0.04564852
+ wua1 = 7.785862e-18
+ pb = 0.6882682
+ wub1 = 2.8560549e-24
+ w0 = 0.0
+ wuc1 = 1.5903152e-16
+ rd = 0
+ rs = 0
+ ua = -9.017296e-10
+ ub = 2.7527719e-18
+ uc = 1.2291169e-10
+ wnfactor = 0.0
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -2.6010536e-8
+ ww = 0.0
+ xw = 9.94224e-9
+ hdif = 2e-7
+ lua1 = 9.129858e-19
+ lub1 = 4.248247e-25
+ la0 = 8.279508e-8
+ luc1 = 3.232822e-17
+ pbswg = 0.6882682
+ wute = 7.881835e-7
+ mjsw = 0.2003879
+ jsw = 1.45e-12
+ lk1 = 4.963488e-8
+ kt1 = -0.226924
+ lk2 = -2.7462524e-8
+ kt2 = -0.029338669
+ llc = -0.039
+ lvoff = -5.449216999999999e-10
+ lln = -1
+ lu0 = 1.7277892e-9
+ ppdiblc2 = -2.2121929e-16
+ lute = 8.209799e-8
+ lua = 3.588764e-18
+ lub = 5.910339e-27
+ luc = 4.360599e-18
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ wpdiblc2 = 1.8349379e-9
+ beta0 = 11.59263
+ pa0 = -7.337964e-14
+ lnfactor = -4.5192e-8
+ nlx = 0.0
+ leta0 = 4.976073409680917e-10
+ letab = -6.844199e-10
+ pk1 = -6.389182e-15
+ pk2 = 5.055259e-15
+ lvsat = -0.00020140363
+ cdsc = 0.0
+ pu0 = -2.4055863e-16
+ lvth0 = 2.7532000000000004e-9
+ prt = 0
+ pua = -4.639069e-23
+ pub = -3.506499e-33
+ puc = -2.2654354e-24
+ cgdo = 3.84825e-10
+ tcjswg = 0.000645489
+ ppclm = 4.042711e-14
+ delta = 0.01
+ cgso = 3.84825e-10
+ rsh = 6.8
+ tcj = 0.001040287
+ lpdiblc2 = 5.053093e-9
+ ua1 = 1.2174792e-9
+ ub1 = -3.81245e-18
+ uc1 = -1.540669e-10
+ tpb = 0.001554306
+ tox = 4.01989464e-9
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ wa0 = 1.4537927e-7
+ nfactor = 1.0
+ ute = -2.1610963
+ cjsw = 1.93852e-10
+ wk1 = 8.868675e-8
+ wk2 = -3.876818e-8
+ wln = 1.0
+ wu0 = -4.860856e-9
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ wua = 4.278473e-16
+ wub = -9.451913e-25
+ wuc = -6.126842e-17
+ wwl = 0.0
+ wwn = 1
+ xti = 3
+ )

.model nch_ff_9 nmos (
+ level = 49
+ cjswg = 3.17352e-10
+ mjswg = 0.43879
+ wub1 = -7.675553e-27
+ wuc1 = -1.4706552e-17
+ hdif = 2e-7
+ wvoff = -2.3388100000000003e-10
+ ags = 0.02
+ wute = 3.836007e-8
+ mjsw = 0.2003879
+ weta0 = 0
+ cit = -0.00010000004
+ wvsat = 0.0
+ dlc = 3e-9
+ k3b = 0.0
+ wvth0 = -1.0228453e-8
+ dwb = 0.0
+ dwg = 0.0
+ capmod = 3
+ cdsc = 0.0
+ cgdo = 3.84825e-10
+ cgso = 3.84825e-10
+ mobmod = 1
+ jsw = 1.45e-12
+ kt1 = -0.2313184
+ lk2 = -3.6153600000000002e-9
+ kt2 = -0.029076951
+ llc = -0.039
+ lln = -1
+ lu0 = 4.5192000000000003e-10
+ cjsw = 1.93852e-10
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ nlx = 0.0
+ nfactor = 1.0
+ xpart = 1
+ pu0 = 0.0
+ prt = 0
+ tnom = 25.0
+ pbswg = 0.6882682
+ rsh = 6.8
+ tcj = 0.001040287
+ ua1 = 1.224e-9
+ pdiblc1 = 1e-6
+ toxm = 4.08e-9
+ pdiblc2 = 0.0007000003
+ ub1 = -1.5012456e-18
+ lvoff = 9.038400000000001e-10
+ uc1 = -6.880516e-11
+ pdiblcb = 0.01
+ pbsw = 0.6882682
+ tpb = 0.001554306
+ pclm = 0.8000001
+ tox = 4.01989464e-9
+ beta0 = 11.59263
+ wa0 = 7.667051e-8
+ leta0 = 3.163440009680917e-10
+ ute = -1.6093186
+ wk1 = -2.074723e-8
+ wk2 = 4.920634e-9
+ tcjswg = 0.000645489
+ wln = 1.0
+ wu0 = 1.0362965e-9
+ lvth0 = -2.621136e-9
+ binunit = 2
+ wua = 1.4309126e-16
+ wub = -1.5411778e-25
+ wuc = -1.4141237e-17
+ wwl = 0.0
+ wwn = 1
+ xti = 3
+ delta = 0.01
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ keta = 0.0010152902
+ dsub = 0.0
+ pnfactor = 0.0
+ wnfactor = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ a0 = 0.3047864
+ a1 = 0.0
+ a2 = 0.99
+ b0 = 0.0
+ b1 = 0.0
+ voff = -0.13648388
+ version = 3.24
+ at = 20000.0
+ cf = 0
+ cj = 0.0009502527
+ ldif = 9e-8
+ ef = 0.874
+ k1 = 0.5610723
+ k2 = -0.0060884483
+ k3 = 0.0
+ em = 30000000.0
+ kt1l = 0.0
+ js = 3.5e-7
+ prwb = 0.0
+ ll = 0.0
+ prwg = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ u0 = 0.037007399999999996
+ pb = 0.6882682
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ua = -9.066409e-10
+ ub = 2.2997995e-18
+ uc = 1.072127e-10
+ eta0 = 5e-5
+ wl = 0.0
+ tcjsw = 0.000645489
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -2.6010536e-8
+ ww = 0.0
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ xw = 9.94224e-9
+ pvag = 0.0
+ etab = -5e-5
+ lnfactor = -4.5192e-8
+ vsat = 93615.37
+ wint = 3e-9
+ pscbe1 = 200000030.0
+ pscbe2 = 1e-6
+ vth0 = 0.42210498
+ pvoff = 9.038400000000001e-16
+ rdsw = 170.0
+ wkt1 = 1.4490446e-9
+ wkt2 = 1.0605161e-11
+ lint = 1e-8
+ wmax = 1.19005776e-6
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 1.3557600041489644e-16
+ wmin = 4.9005776e-7
+ nqsmod = 0
+ tpbswg = 0.001554306
+ noimod = 2
+ lmax = 2.0001e-5
+ wketa = 2.1944087e-10
+ pvth0 = -2.71152e-15
+ lmin = 1.0006010536e-5
+ drout = 0.0
+ tpbsw = 0.001554306
+ )

.model nch_ff_10 nmos (
+ level = 49
+ lute = -1.2190513e-8
+ nqsmod = 0
+ tpbswg = 0.001554306
+ noimod = 2
+ cdsc = 0.0
+ cgdo = 3.84825e-10
+ nfactor = 1.0
+ lketa = -2.8027248e-8
+ cgso = 3.84825e-10
+ xpart = 1
+ cjsw = 1.93852e-10
+ pbswg = 0.6882682
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0003968185
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ pdiblcb = 0.01
+ lpscbe1 = 262.58185
+ lvoff = -2.6983819999999998e-9
+ capmod = 3
+ beta0 = 11.59263
+ tnom = 25.0
+ leta0 = 3.163440009680917e-10
+ binunit = 2
+ lvsat = -0.006201102
+ toxm = 4.08e-9
+ lvth0 = 6.329934400000001e-8
+ pcit = 4.302753e-19
+ pbsw = 0.6882682
+ pclm = 0.7699873
+ ppclm = 1.243718e-13
+ mobmod = 1
+ delta = 0.01
+ ags = 0.02
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ cit = -0.00012672294
+ dlc = 3e-9
+ k3b = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ pnfactor = 0.0
+ pkt1 = 7.833639e-15
+ pkt2 = 9.747044e-16
+ keta = 0.00382927
+ wnfactor = 0.0
+ pketa = -6.831802e-16
+ version = 3.24
+ dsub = 0.0
+ wpclm = -1.2487239e-8
+ wcit = -4.317371e-14
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ la0 = -1.9725388e-7
+ tcjsw = 0.000645489
+ jsw = 1.45e-12
+ tcjswg = 0.000645489
+ lk1 = 1.0512358e-8
+ kt1 = -0.2310088
+ lk2 = -9.025411e-9
+ kt2 = -0.028688708
+ lcit = 2.6616018e-10
+ llc = -0.039
+ lln = -1
+ voff = -0.13612218
+ lu0 = 4.157672e-9
+ lnfactor = -4.5192e-8
+ ldif = 9e-8
+ lua = -1.9124487e-16
+ lub = 4.117038e-25
+ luc = 4.038815e-17
+ nch = 3.9e+17
+ pvoff = -4.352292e-15
+ lwl = 0.0
+ lwn = 1.0
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ pub1 = -1.8996434e-32
+ puc1 = 1.3569954e-23
+ pa0 = -1.0015934e-13
+ nlx = 0.0
+ eta0 = 5e-5
+ pk1 = -1.457495e-14
+ pk2 = 2.2122807e-15
+ pvag = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ etab = -5e-5
+ peta0 = 1.3557600041489644e-16
+ vsat = 94237.97
+ wint = 3e-9
+ pu0 = 1.6856667e-15
+ pute = -3.577514e-14
+ pvsat = 1.2437262e-9
+ vth0 = 0.41548638
+ prt = 0
+ pua = 4.758471e-23
+ pub = -5.695533e-32
+ puc = -9.239189e-24
+ lpdiblc2 = 3.0196912e-9
+ wketa = 2.8803285e-10
+ rdsw = 170.0
+ pvth0 = -9.869192e-15
+ wkt1 = 6.625341e-10
+ wkt2 = -8.725676e-11
+ drout = 0.0
+ lint = 1e-8
+ rsh = 6.8
+ tpbsw = 0.001554306
+ wmax = 1.19005776e-6
+ tcj = 0.001040287
+ ua1 = 1.224e-9
+ ub1 = -1.5338095e-18
+ uc1 = -7.316409e-11
+ wmin = 4.9005776e-7
+ lkt1 = -3.0828107e-9
+ lkt2 = -3.866881e-9
+ tpb = 0.001554306
+ tox = 4.01989464e-9
+ cjswg = 3.17352e-10
+ lmax = 1.0006010536e-5
+ wa0 = 8.672666e-8
+ lmin = 1.2060105359999999e-6
+ ute = -1.6080947
+ mjswg = 0.43879
+ wk1 = -1.9283881e-8
+ wk2 = 4.698517e-9
+ wln = 1.0
+ wu0 = 8.670528e-10
+ wvoff = 2.938435e-10
+ wua = 1.3831368e-16
+ wub = -1.4839938e-25
+ wuc = -1.3213606e-17
+ wwl = 0.0
+ wwn = 1
+ xti = 3
+ a0 = 0.324591
+ a1 = 0.0
+ a2 = 0.99
+ b0 = 0.0
+ b1 = 0.0
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ wub1 = -5.768295e-27
+ wuc1 = -1.6068998e-17
+ weta0 = 0
+ at = 20000.0
+ cf = 0
+ cj = 0.0009502527
+ ef = 0.874
+ k1 = 0.5600169
+ k2 = -0.005545271300000001
+ k3 = 0.0
+ em = 30000000.0
+ hdif = 2e-7
+ wvsat = -0.00012487893
+ js = 3.5e-7
+ pscbe1 = 173636400.0
+ pscbe2 = 1e-6
+ ll = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ u0 = 0.03663534
+ pb = 0.6882682
+ lub1 = 3.243357e-25
+ lpclm = 2.9892766e-7
+ wvth0 = -9.50981e-9
+ luc1 = 4.341489e-17
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ wute = 4.195195e-8
+ ua = -8.874397e-10
+ ub = 2.2584638e-18
+ uc = 1.0315766e-10
+ mjsw = 0.2003879
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -2.6010536e-8
+ ww = 0.0
+ xw = 9.94224e-9
+ )

.model nch_ff_11 nmos (
+ level = 49
+ lvoff = 1.2067069999999999e-8
+ wcit = 5.431231e-13
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ ags = 0.02
+ beta0 = 11.59263
+ leta0 = 3.544583009680917e-10
+ lcit = 3.0283653e-10
+ cit = -0.0001583405
+ letab = -3.81143e-11
+ voff = -0.14885098
+ ldif = 9e-8
+ lvsat = -0.0007659488
+ dlc = 3e-9
+ kt1l = 0.0
+ mobmod = 1
+ prwb = 0.0
+ lvth0 = 7.488615e-9
+ prwg = 0.0
+ pub1 = -5.874811e-31
+ puc1 = -3.67348e-23
+ a0 = -0.1914371
+ a1 = 0.0
+ a2 = 0.99
+ k3b = 0.0
+ b0 = 0.0
+ b1 = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ eta0 = 1.7142847e-5
+ at = 20000.0
+ cf = 0
+ cj = 0.0009502527
+ ef = 0.874
+ k1 = 0.5552615
+ ppclm = 7.308824e-14
+ k2 = -0.0036859210000000004
+ k3 = 0.0
+ em = 30000000.0
+ pvag = 0.0
+ etab = -1.7142847e-5
+ delta = 0.01
+ js = 3.5e-7
+ vsat = 89552.49
+ ll = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ u0 = 0.03761954
+ pb = 0.6882682
+ wint = 3e-9
+ pute = -2.0303331e-13
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ua = -1.3333591e-9
+ ub = 2.969086e-18
+ uc = 1.6160392e-10
+ vth0 = 0.46359908
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -2.6010536e-8
+ ww = 0.0
+ xw = 9.94224e-9
+ rdsw = 170.0
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ wkt1 = 1.1898274e-8
+ wkt2 = 2.0987987e-9
+ lint = 1e-8
+ wmax = 1.19005776e-6
+ la0 = 4.013388e-7
+ wmin = 4.9005776e-7
+ lkt1 = 9.329063e-9
+ lkt2 = 2.691467e-9
+ jsw = 1.45e-12
+ lk1 = 1.6028618e-8
+ kt1 = -0.2417087
+ lk2 = -1.1182256000000001e-8
+ kt2 = -0.03434246
+ lmax = 1.2060105359999999e-6
+ llc = -0.039
+ lln = -1
+ lu0 = 3.0160021e-9
+ lmin = 5.06010536e-7
+ lua = 3.260216e-16
+ lub = -4.12618e-25
+ luc = -2.7409531e-17
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ pketa = 1.4501565e-15
+ pa0 = 1.1848049e-14
+ nlx = 0.0
+ pk1 = 7.144098e-15
+ pk2 = -4.137203e-15
+ pu0 = -1.1138246e-15
+ wpclm = 3.172275e-8
+ wub1 = 4.843047e-25
+ prt = 0
+ wuc1 = 2.7297169e-17
+ pua = -1.3255767e-22
+ pub = 5.546348e-32
+ puc = -6.669366e-24
+ tcjswg = 0.000645489
+ hdif = 2e-7
+ tcjsw = 0.000645489
+ rsh = 6.8
+ lub1 = 4.951269e-25
+ luc1 = 6.070172e-17
+ tcj = 0.001040287
+ ua1 = 1.224e-9
+ ub1 = -1.6810433e-18
+ uc1 = -8.806652e-11
+ wute = 1.8614003e-7
+ mjsw = 0.2003879
+ pvoff = 3.7090935e-15
+ tpb = 0.001554306
+ tox = 4.01989464e-9
+ wa0 = -9.831444e-9
+ lute = 2.2508574e-7
+ ute = -1.8126432
+ wk1 = -3.80072e-8
+ wk2 = 1.0172209e-8
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 1.3557600041489644e-16
+ wln = 1.0
+ wu0 = 3.280407e-9
+ wua = 2.9360883e-16
+ pvsat = 4.380818e-12
+ wub = -2.4531215e-25
+ wuc = -1.542897e-17
+ wwl = 0.0
+ wwn = 1
+ cdsc = 0.0
+ wketa = -1.5510503e-9
+ pvth0 = -3.2494082e-15
+ xti = 3
+ drout = 0.0
+ cgdo = 3.84825e-10
+ tpbsw = 0.001554306
+ cgso = 3.84825e-10
+ cjswg = 3.17352e-10
+ nfactor = 1.0
+ mjswg = 0.43879
+ pnfactor = 0.0
+ cjsw = 1.93852e-10
+ wnfactor = 0.0
+ wvoff = -6.655627e-9
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ weta0 = 0
+ pscbe1 = 400000100.0
+ pscbe2 = 1e-6
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0011219129
+ pdiblcb = 0.01
+ wvsat = 0.0009435224
+ ppdiblc2 = 1.2928064e-16
+ tnom = 25.0
+ lpclm = 9.659676e-8
+ wvth0 = -1.5216522e-8
+ wpdiblc2 = -1.1144895e-10
+ lnfactor = -4.5192e-8
+ nqsmod = 0
+ tpbswg = 0.001554306
+ toxm = 4.08e-9
+ noimod = 2
+ pcit = -2.4980728e-19
+ binunit = 2
+ pbsw = 0.6882682
+ pclm = 0.9444105
+ lpdiblc2 = 2.1785818e-9
+ lketa = -2.9090079e-9
+ xpart = 1
+ pkt1 = -5.199821e-15
+ pkt2 = -1.5611203e-15
+ keta = -0.017824383
+ pbswg = 0.6882682
+ dsub = 0.0
+ capmod = 3
+ version = 3.24
+ )

.model nch_ff_12 nmos (
+ level = 49
+ tpb = 0.001554306
+ tox = 4.01989464e-9
+ wa0 = 1.7605426e-7
+ pketa = -7.367843e-16
+ cjsw = 1.93852e-10
+ nfactor = 1.0
+ ute = -1.2073984
+ wk1 = -1.7855582e-8
+ wk2 = 1.6966123e-9
+ tcjswg = 0.000645489
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ wln = 1.0
+ wu0 = -4.268465e-11
+ wpclm = 1.9327061e-7
+ wua = -1.9101984e-17
+ wub = -5.11281e-26
+ wuc = -9.012729e-18
+ wwl = 0.0
+ wwn = 1
+ xti = 3
+ tcjsw = 0.000645489
+ tnom = 25.0
+ pdiblc1 = 1e-6
+ pdiblc2 = -0.00401322
+ pags = 1.8981756e-15
+ pdiblcb = 0.01
+ pvoff = -1.3169074e-15
+ toxm = 4.08e-9
+ pcit = -1.4232223e-17
+ pbsw = 0.6882682
+ pclm = 0.9948969
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 1.2420400941489644e-16
+ petab = 1.3954016e-17
+ binunit = 2
+ pvsat = 1.606088e-11
+ wketa = 3.203169e-9
+ pvth0 = 4.495999999999906e-18
+ drout = 0.0
+ tpbsw = 0.001554306
+ a0 = 0.5005398
+ a1 = 0.0
+ a2 = 0.99
+ b0 = 0.0
+ b1 = 0.0
+ at = 20000.0
+ cf = 0
+ cj = 0.0009502527
+ ef = 0.874
+ k1 = 0.489967
+ k2 = 0.022067764
+ k3 = 0.0
+ em = 30000000.0
+ js = 3.5e-7
+ cjswg = 3.17352e-10
+ ll = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ u0 = 0.041613199999999996
+ pb = 0.6882682
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ua = -5.274002e-10
+ ub = 2.0039751e-18
+ uc = 7.914647e-11
+ mjswg = 0.43879
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -2.6010536e-8
+ ww = 0.0
+ xw = 9.94224e-9
+ pkt1 = 2.3961372e-15
+ pkt2 = 8.832021e-16
+ keta = -0.027587207
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ wvoff = 4.2704619999999996e-9
+ wags = -4.12647e-9
+ dsub = 0.0
+ pscbe1 = 400000000.0
+ pscbe2 = 1e-6
+ weta0 = 2.4721704e-11
+ lags = -9.594464e-9
+ wetab = -3.0334849e-11
+ wcit = 3.093965e-11
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ wvsat = 0.000918131
+ version = 3.24
+ nqsmod = 0
+ lpclm = 7.337301e-8
+ wvth0 = -2.2290227000000003e-8
+ tpbswg = 0.001554306
+ noimod = 2
+ lcit = 1.2733804e-10
+ voff = -0.12370098000000002
+ ldif = 9e-8
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ pub1 = 1.6165291e-31
+ puc1 = 2.0250814e-23
+ eta0 = -0.00031223928
+ pvag = 0.0
+ etab = 0.0014101875
+ vsat = 88351.66
+ wint = 3e-9
+ pute = 4.383575e-14
+ vth0 = 0.47062918
+ rdsw = 170.0
+ wkt1 = -4.614678e-9
+ wkt2 = -3.214946e-9
+ lint = 1e-8
+ wmax = 1.19005776e-6
+ ags = 0.04085753
+ lketa = 1.5818911e-9
+ wmin = 4.9005776e-7
+ lkt1 = 1.6202869e-9
+ lkt2 = -8.228257e-11
+ lmax = 5.06010536e-7
+ xpart = 1
+ cit = 0.00022317801
+ lmin = 1.8e-7
+ pnfactor = 0.0
+ dlc = 3e-9
+ wnfactor = 0.0
+ k3b = 0.0
+ capmod = 3
+ dwb = 0.0
+ dwg = 0.0
+ pbswg = 0.6882682
+ lvoff = 4.980705000000001e-10
+ wub1 = -1.1442477e-24
+ wuc1 = -9.658459e-17
+ ppdiblc2 = 3.905237e-16
+ hdif = 2e-7
+ beta0 = 11.59263
+ wpdiblc2 = -6.793707e-10
+ lub1 = -6.558089e-26
+ leta0 = 5.059740609680917e-10
+ luc1 = -7.416688e-18
+ wute = -3.505318e-7
+ mobmod = 1
+ la0 = 8.302936e-8
+ letab = -6.946862e-10
+ lnfactor = -4.5192e-8
+ mjsw = 0.2003879
+ lvsat = -0.00021356932
+ jsw = 1.45e-12
+ lk1 = 4.606408e-8
+ kt1 = -0.2249505
+ lk2 = -2.3028953000000002e-8
+ kt2 = -0.028312566
+ lvth0 = 4.254808999999999e-9
+ llc = -0.039
+ lln = -1
+ lute = -5.332685e-8
+ lu0 = 1.1789145e-9
+ lua = -4.471944e-17
+ lub = 3.1333025e-26
+ luc = 1.0520902e-17
+ ppclm = -1.2237712e-15
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ delta = 0.01
+ pa0 = -7.365936e-14
+ nlx = 0.0
+ lpdiblc2 = 4.540744e-9
+ cdsc = 0.0
+ pk1 = -2.1256446e-15
+ pk2 = -2.3842633e-16
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ pu0 = 4.147977e-16
+ cgdo = 3.84825e-10
+ prt = 0
+ pua = 1.1289303e-23
+ pub = -3.386118e-32
+ puc = -9.620837e-24
+ cgso = 3.84825e-10
+ rsh = 6.8
+ tcj = 0.001040287
+ ua1 = 1.224e-9
+ ub1 = -4.621132e-19
+ uc1 = 6.001696e-11
+ )

.model nch_ff_13 nmos (
+ level = 49
+ drout = 0.0
+ wkt1 = 5.128653e-9
+ wkt2 = 3.532295e-9
+ tpbsw = 0.001554306
+ lint = 1e-8
+ wmax = 4.9005776e-7
+ wmin = 2.2e-7
+ cjswg = 3.17352e-10
+ lmax = 2.0001e-5
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ mjswg = 0.43879
+ lmin = 1.0006010536e-5
+ pscbe1 = 200000030.0
+ pscbe2 = 1e-6
+ wvoff = -1.0949902e-9
+ weta0 = 0
+ nqsmod = 0
+ wub1 = -4.432931e-26
+ wuc1 = -1.7086574e-17
+ tpbswg = 0.001554306
+ wvsat = 0.0
+ noimod = 2
+ hdif = 2e-7
+ wvth0 = -2.1421089000000002e-8
+ ags = 0.02
+ wute = 2.5547985e-8
+ mjsw = 0.2003879
+ cit = -9.999998e-5
+ dlc = 3e-9
+ k3b = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ cdsc = 0.0
+ cgdo = 3.84825e-10
+ cgso = 3.84825e-10
+ xpart = 1
+ jsw = 1.45e-12
+ capmod = 3
+ kt1 = -0.238767
+ lk2 = -3.6153600000000002e-9
+ kt2 = -0.03620588
+ llc = -0.039
+ cjsw = 1.93852e-10
+ lln = -1
+ a0 = 0.352982
+ a1 = 0.0
+ a2 = 0.99
+ lu0 = 4.5192000000000003e-10
+ b0 = 0.0
+ b1 = 0.0
+ pbswg = 0.6882682
+ nch = 3.9e+17
+ at = 20000.0
+ cf = 0
+ cj = 0.0009502527
+ lwl = 0.0
+ lwn = 1.0
+ ef = 0.874
+ k1 = 0.5220979
+ k2 = 0.009311849
+ k3 = 0.0
+ em = 30000000.0
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ nfactor = 1.0
+ js = 3.5e-7
+ ll = 0.0
+ nlx = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ lvoff = 9.038400000000001e-10
+ u0 = 0.0371451
+ pb = 0.6882682
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ua = -5.860608e-10
+ ub = 1.7266676e-18
+ uc = 7.252202e-11
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -2.6010536e-8
+ ww = 0.0
+ xw = 9.94224e-9
+ mobmod = 1
+ beta0 = 11.59263
+ pu0 = 0.0
+ tnom = 25.0
+ leta0 = 3.163440009680917e-10
+ prt = 0
+ toxm = 4.08e-9
+ rsh = 6.8
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0006999999
+ lvth0 = -2.621136e-9
+ tcj = 0.001040287
+ ua1 = 1.224e-9
+ ub1 = -1.4270478e-18
+ uc1 = -6.39873e-11
+ pdiblcb = 0.01
+ pbsw = 0.6882682
+ pclm = 0.7999999
+ tpb = 0.001554306
+ tox = 4.01989464e-9
+ delta = 0.01
+ wa0 = 5.286186e-8
+ ute = -1.5833832
+ wk1 = -1.4938487e-9
+ wk2 = -2.6871128e-9
+ dvt0w = 0.0
+ dvt1w = 0.0
+ wln = 1.0
+ dvt2w = 0.0
+ wu0 = 9.682726e-10
+ binunit = 2
+ wua = -1.5275344e-17
+ wub = 1.2900942e-25
+ wuc = 2.9959555e-18
+ wwl = 0.0
+ wwn = 1
+ xti = 3
+ pnfactor = 0.0
+ keta = 0.002064252
+ tcjswg = 0.000645489
+ wnfactor = 0.0
+ dsub = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ tcjsw = 0.000645489
+ lnfactor = -4.5192e-8
+ voff = -0.13474068
+ version = 3.24
+ pvoff = 9.038400000000001e-16
+ ldif = 9e-8
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ eta0 = 5e-5
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 1.3557600041489644e-16
+ pvag = 0.0
+ etab = -5e-5
+ vsat = 93615.35
+ wint = 3e-9
+ vth0 = 0.44476208
+ wketa = -2.9874625e-10
+ pvth0 = -2.71152e-15
+ rdsw = 170.0
+ )

.model nch_ff_14 nmos (
+ level = 49
+ la0 = -2.4964379e-7
+ pcit = 1.5653096e-18
+ pbsw = 0.6882682
+ pclm = 0.7606163
+ jsw = 1.45e-12
+ lk1 = -6.331243e-8
+ kt1 = -0.2407974
+ lk2 = 1.7183372000000002e-8
+ kt2 = -0.03589625
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0003968183
+ pdiblcb = 0.01
+ lpscbe1 = 262.58182
+ llc = -0.039
+ lln = -1
+ lu0 = 1.0346475000000001e-8
+ lpdiblc2 = 3.0196909e-9
+ lua = -1.2876533e-16
+ lub = 7.836163e-25
+ luc = 7.064626e-17
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ pa0 = -7.427873e-14
+ nlx = 0.0
+ pk1 = 2.1894499e-14
+ pk2 = -1.0734859e-14
+ lketa = -3.0377027e-8
+ binunit = 2
+ pu0 = -1.3716021e-15
+ capmod = 3
+ prt = 0
+ pua = 1.6719826e-23
+ pub = -2.4068014e-31
+ xpart = 1
+ puc = -2.4186704e-23
+ pkt1 = -3.679308e-15
+ pkt2 = 5.879336e-16
+ rsh = 6.8
+ keta = 0.005114151
+ tcj = 0.001040287
+ ua1 = 1.224e-9
+ ub1 = -1.4513121e-18
+ uc1 = -6.991786e-11
+ pbswg = 0.6882682
+ tpb = 0.001554306
+ tox = 4.01989464e-9
+ dsub = 0.0
+ wa0 = 6.031956e-8
+ lvoff = -1.8823532e-8
+ mobmod = 1
+ ute = -1.5785241
+ wk1 = -3.692092e-9
+ wk2 = -1.6093152e-9
+ wcit = -1.5715551e-13
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ wln = 1.0
+ beta0 = 11.59263
+ wu0 = 1.1059835e-9
+ wua = -1.6954039e-17
+ wub = 1.5317406e-25
+ wuc = 5.42434e-18
+ leta0 = 3.163440009680917e-10
+ wwl = 0.0
+ wwn = 1
+ lcit = 2.6386249e-10
+ xti = 3
+ voff = -0.13276008
+ lvsat = -0.005267757
+ ldif = 9e-8
+ lvth0 = 5.3657104e-8
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ pub1 = 2.1839324e-32
+ puc1 = 5.837128e-24
+ version = 3.24
+ ppclm = 7.826515e-14
+ eta0 = 5e-5
+ delta = 0.01
+ pvag = 0.0
+ etab = -5e-5
+ vsat = 94144.24
+ wint = 3e-9
+ pute = -1.7889165e-14
+ vth0 = 0.43911168
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ rdsw = 170.0
+ wkt1 = 5.498062e-9
+ wkt2 = 3.473265e-9
+ lint = 1e-8
+ wmax = 4.9005776e-7
+ wmin = 2.2e-7
+ lkt1 = 2.0222748e-8
+ lkt2 = -3.0839447e-9
+ lmax = 1.0006010536e-5
+ tcjswg = 0.000645489
+ lmin = 1.2060105359999999e-6
+ pketa = 4.776125e-16
+ wpclm = -7.857923e-9
+ wub1 = -4.652201e-26
+ wuc1 = -1.7672629e-17
+ tcjsw = 0.000645489
+ hdif = 2e-7
+ lub1 = 2.4167225e-25
+ a0 = 0.3780467
+ a1 = 0.0
+ a2 = 0.99
+ luc1 = 5.906839e-17
+ b0 = 0.0
+ b1 = 0.0
+ wute = 2.7344081e-8
+ mjsw = 0.2003879
+ at = 20000.0
+ pvoff = 3.6135329e-15
+ cf = 0
+ cj = 0.0009502527
+ ef = 0.874
+ k1 = 0.5284545
+ k2 = 0.007223622
+ k3 = 0.0
+ em = 30000000.0
+ js = 3.5e-7
+ ll = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ u0 = 0.03615168
+ pb = 0.6882682
+ w0 = 0.0
+ rd = 0
+ lute = -4.839696e-8
+ rs = 0
+ ua = -5.731325e-10
+ ub = 1.6479914e-18
+ uc = 6.542903e-11
+ cdscb = 0.0
+ cdscd = 0.0
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -2.6010536e-8
+ ww = 0.0
+ peta0 = 1.3557600041489644e-16
+ xw = 9.94224e-9
+ pvsat = 7.826533e-10
+ wketa = -3.466991e-10
+ pvth0 = -5.1059225e-15
+ cdsc = 0.0
+ drout = 0.0
+ tpbsw = 0.001554306
+ cgdo = 3.84825e-10
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ cgso = 3.84825e-10
+ cjswg = 3.17352e-10
+ pscbe1 = 173636400.0
+ pscbe2 = 1e-6
+ mjswg = 0.43879
+ ags = 0.02
+ pnfactor = 0.0
+ wnfactor = 0.0
+ wvoff = -1.3670473000000001e-9
+ cjsw = 1.93852e-10
+ cit = -0.00012649217
+ nqsmod = 0
+ dlc = 3e-9
+ tpbswg = 0.001554306
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ noimod = 2
+ k3b = 0.0
+ weta0 = 0
+ dwb = 0.0
+ dwg = 0.0
+ wvsat = -7.857954e-5
+ nfactor = 1.0
+ lpclm = 3.92261e-7
+ wvth0 = -2.1180688000000003e-8
+ tnom = 25.0
+ lnfactor = -4.5192e-8
+ toxm = 4.08e-9
+ )

.model nch_ff_15 nmos (
+ level = 49
+ wub1 = -1.0574451e-25
+ wuc1 = -4.040928e-17
+ ppdiblc2 = 4.703685e-16
+ beta0 = 11.59263
+ hdif = 2e-7
+ wpdiblc2 = -4.054901e-10
+ leta0 = 3.544582809680917e-10
+ lub1 = -8.773805e-25
+ luc1 = -7.886598e-17
+ letab = -3.811428e-11
+ lnfactor = -4.5192e-8
+ wute = 1.9757099e-8
+ lvsat = -0.0007893788
+ mjsw = 0.2003879
+ lvth0 = 6.2381230000000005e-9
+ lute = -1.6751561e-7
+ ppclm = 4.863229e-14
+ delta = 0.01
+ lpdiblc2 = 1.4881204e-9
+ dvt0w = 0.0
+ cdsc = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ cgdo = 3.84825e-10
+ tcjswg = 0.000645489
+ cgso = 3.84825e-10
+ pketa = 3.1429577e-15
+ cjsw = 1.93852e-10
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ wpclm = 1.7687656e-8
+ tcjsw = 0.000645489
+ tnom = 25.0
+ nfactor = 1.0
+ pvoff = -4.799142e-16
+ toxm = 4.08e-9
+ ags = 0.02
+ pcit = -9.088336e-19
+ pbsw = 0.6882682
+ pclm = 0.9728217
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 1.3557600041489644e-16
+ pvsat = 1.5955267e-11
+ cit = -0.00016124053
+ wketa = -2.6444102e-9
+ pvth0 = -2.63166535e-15
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0017171376
+ dlc = 3e-9
+ drout = 0.0
+ pdiblcb = 0.01
+ k3b = 0.0
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ tpbsw = 0.001554306
+ dwb = 0.0
+ dwg = 0.0
+ pscbe1 = 400000100.0
+ pscbe2 = 1e-6
+ cjswg = 3.17352e-10
+ mjswg = 0.43879
+ binunit = 2
+ pkt1 = -1.1651986e-14
+ pkt2 = -1.4582807e-15
+ keta = -0.015611105
+ nqsmod = 0
+ wvoff = 2.1617860000000002e-9
+ tpbswg = 0.001554306
+ la0 = 2.7901473e-7
+ noimod = 2
+ jsw = 1.45e-12
+ dsub = 0.0
+ lk1 = 6.936774e-8
+ kt1 = -0.2426658
+ lk2 = -3.5143967e-8
+ kt2 = -0.04069558
+ llc = -0.039
+ lln = -1
+ weta0 = 0
+ lu0 = -1.2926906e-9
+ lua = 6.135559e-17
+ lub = -2.9489129e-25
+ luc = -2.7169401e-17
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ wvsat = 0.0005823669
+ wcit = 1.975718e-12
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ pa0 = 7.227613e-14
+ nlx = 0.0
+ lpclm = 1.4610272e-7
+ wvth0 = -2.3313668000000003e-8
+ pk1 = -1.920543e-14
+ pk2 = 7.699883e-15
+ lcit = 3.0417063e-10
+ voff = -0.16670008
+ pu0 = 1.0146696e-15
+ ldif = 9e-8
+ prt = 0
+ pua = -1.8126578e-24
+ pub = -2.6935e-33
+ puc = -6.78799e-24
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ pub1 = 9.053745e-32
+ puc1 = 3.221165e-23
+ eta0 = 1.7142866e-5
+ rsh = 6.8
+ pvag = 0.0
+ etab = -1.7142866e-5
+ tcj = 0.001040287
+ ua1 = 1.224e-9
+ ub1 = -4.866116e-19
+ uc1 = 4.899104e-11
+ vsat = 90283.57
+ version = 3.24
+ a0 = -0.07769345
+ wint = 3e-9
+ a1 = 0.0
+ a2 = 0.99
+ pute = -9.088265e-15
+ b0 = 0.0
+ b1 = 0.0
+ tpb = 0.001554306
+ vth0 = 0.47999008
+ tox = 4.01989464e-9
+ at = 20000.0
+ cf = 0
+ cj = 0.0009502527
+ ef = 0.874
+ k1 = 0.4140751
+ k2 = 0.052333399999999995
+ k3 = 0.0
+ rdsw = 170.0
+ wa0 = -6.602082e-8
+ em = 30000000.0
+ js = 3.5e-7
+ wkt1 = 1.2371058e-8
+ wkt2 = 5.237243e-9
+ ute = -1.4758356
+ ll = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ lint = 1e-8
+ u0 = 0.04618544
+ pb = 0.6882682
+ wk1 = 3.173889e-8
+ wk2 = -1.7501334e-8
+ w0 = 0.0
+ rd = 0
+ wmax = 4.9005776e-7
+ lketa = -6.33573e-9
+ capmod = 3
+ rs = 0
+ ua = -7.370299e-10
+ ub = 2.5777392e-18
+ uc = 1.4975288e-10
+ wln = 1.0
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -2.6010536e-8
+ ww = 0.0
+ wmin = 2.2e-7
+ wu0 = -9.511471e-10
+ xw = 9.94224e-9
+ lkt1 = 2.2390124e-8
+ wua = -9.777621e-19
+ lkt2 = 2.4832894e-9
+ wub = -5.19868e-26
+ wuc = -9.57455e-18
+ xpart = 1
+ wwl = 0.0
+ wwn = 1
+ lmax = 1.2060105359999999e-6
+ xti = 3
+ lmin = 5.06010536e-7
+ pnfactor = 0.0
+ wnfactor = 0.0
+ pbswg = 0.6882682
+ mobmod = 1
+ lvoff = 2.0546844000000002e-8
+ )

.model nch_ff_16 nmos (
+ level = 49
+ at = 20000.0
+ cf = 0
+ cj = 0.0009502527
+ ef = 0.874
+ k1 = 0.4942783
+ k2 = 0.016287533
+ k3 = 0.0
+ em = 30000000.0
+ pketa = -1.9609824e-16
+ pkt1 = 3.435378e-15
+ pkt2 = -8.505888e-17
+ wnfactor = 0.0
+ keta = -0.030443965
+ js = 3.5e-7
+ ll = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ ags = 0.0548038
+ u0 = 0.03891118
+ pb = 0.6882682
+ w0 = 0.0
+ binunit = 2
+ rd = 0
+ rs = 0
+ ua = -6.614348e-10
+ ub = 2.1301375e-18
+ uc = 1.2526492e-10
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ wags = -1.1015922e-8
+ xl = -2.6010536e-8
+ ww = 0.0
+ dsub = 0.0
+ xw = 9.94224e-9
+ wpclm = 1.2379924e-7
+ cit = 0.00029138371
+ lags = -1.6009743e-8
+ dlc = 3e-9
+ wcit = -2.7539906e-12
+ ppdiblc2 = -1.1422951e-16
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ tcjsw = 0.000645489
+ k3b = 0.0
+ wpdiblc2 = 8.65375e-10
+ dwb = 0.0
+ dwg = 0.0
+ lnfactor = -4.5192e-8
+ lcit = 9.596344e-11
+ pvoff = 4.069063000000001e-16
+ voff = -0.11552988
+ ldif = 9e-8
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ pub1 = -3.181536e-32
+ puc1 = -1.1609298e-23
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 1.3557600041489644e-16
+ eta0 = -0.00026219533
+ pvag = 0.0
+ etab = 0.0013487812
+ pvsat = 1.2452966e-11
+ la0 = 1.1871046e-7
+ vsat = 89015.94
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ wint = 3e-9
+ pute = -6.731688e-15
+ wketa = 4.614407e-9
+ lpdiblc2 = 5.562512e-9
+ pvth0 = -3.7536774e-15
+ jsw = 1.45e-12
+ vth0 = 0.46776328
+ lk1 = 3.247429e-8
+ kt1 = -0.1929406
+ lk2 = -1.8562871999999998e-8
+ kt2 = -0.03937921
+ drout = 0.0
+ rdsw = 170.0
+ llc = -0.039
+ lln = -1
+ tpbsw = 0.001554306
+ pscbe1 = 400000000.0
+ pscbe2 = 1e-6
+ lu0 = 2.0534652e-9
+ version = 3.24
+ wkt1 = -2.0427562e-8
+ wkt2 = 2.2519782e-9
+ lint = 1e-8
+ lua = 2.6581833e-17
+ lub = -8.899446e-26
+ luc = -1.5904941e-17
+ nch = 3.9e+17
+ wmax = 4.9005776e-7
+ lwl = 0.0
+ lwn = 1.0
+ wmin = 2.2e-7
+ pa0 = -9.128582e-14
+ nlx = 0.0
+ cjswg = 3.17352e-10
+ lkt1 = -4.834396e-10
+ lkt2 = 1.8777602e-9
+ mjswg = 0.43879
+ pk1 = 4.587708e-15
+ pk2 = -2.4446703e-15
+ lmax = 5.06010536e-7
+ nqsmod = 0
+ tpbswg = 0.001554306
+ lmin = 1.8e-7
+ noimod = 2
+ pu0 = -1.7230291e-17
+ prt = 0
+ pua = -2.3933522e-23
+ pub = 2.5580594e-32
+ puc = 3.433529e-24
+ wvoff = 2.33915e-10
+ rsh = 6.8
+ tcj = 0.001040287
+ ua1 = 1.224e-9
+ ub1 = -3.1027764e-18
+ uc1 = -2.4653823e-10
+ weta0 = 0
+ tpb = 0.001554306
+ wub1 = 1.602399e-25
+ wuc1 = 5.485366e-17
+ tox = 4.01989464e-9
+ wvsat = 0.0005899806
+ wa0 = 2.8954867e-7
+ hdif = 2e-7
+ lpclm = 7.125815e-8
+ wvth0 = -2.0874508000000002e-8
+ ute = -1.9466008
+ wk1 = -1.9985334e-8
+ wk2 = 4.552045e-9
+ lub1 = 3.260553e-25
+ luc1 = 5.707747e-17
+ wute = 1.4634106e-8
+ wln = 1.0
+ mjsw = 0.2003879
+ wu0 = 1.2921135e-9
+ wua = 4.711108e-17
+ wub = -1.1345223e-25
+ wuc = -3.179524e-17
+ wwl = 0.0
+ wwn = 1
+ xti = 3
+ lute = 4.90364e-8
+ cdsc = 0.0
+ capmod = 3
+ cgdo = 3.84825e-10
+ lketa = 4.87385e-10
+ cgso = 3.84825e-10
+ xpart = 1
+ mobmod = 1
+ cjsw = 1.93852e-10
+ pbswg = 0.6882682
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ lvoff = -2.9914309999999998e-9
+ beta0 = 11.59263
+ leta0 = 4.829538409680917e-10
+ tnom = 25.0
+ letab = -6.664392e-10
+ lvsat = -0.00020626588
+ pags = 5.067323e-15
+ lvth0 = 1.1862447e-8
+ toxm = 4.08e-9
+ nfactor = 1.0
+ pcit = 1.266836e-18
+ ppclm = -1.7902992e-16
+ pbsw = 0.6882682
+ pclm = 1.1355271
+ delta = 0.01
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ tcjswg = 0.000645489
+ pdiblc1 = 1e-6
+ pdiblc2 = -0.007140237
+ pdiblcb = 0.01
+ a0 = 0.270794
+ a1 = 0.0
+ a2 = 0.99
+ b0 = 0.0
+ b1 = 0.0
+ pnfactor = 0.0
+ )

.model nch_tt_1 nmos (
+ level = 49
+ cjsw = 2.040547e-10
+ drout = 0.0
+ tpbsw = 0.001554306
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ cjswg = 3.340547e-10
+ pnfactor = 0.0
+ mjswg = 0.43879
+ wnfactor = 0.0
+ tnom = 25.0
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ wvoff = 0.0
+ pscbe1 = 200000030.0
+ pscbe2 = 1e-6
+ toxm = 4.08e-9
+ version = 3.24
+ pbsw = 0.6882682
+ pclm = 0.8000001
+ weta0 = 0
+ wvsat = 0.0
+ nqsmod = 0
+ lnfactor = 0.0
+ tpbswg = 0.001554306
+ wvth0 = 0.0
+ noimod = 2
+ ags = 0.02
+ keta = 0.009263485
+ cit = -0.00010000001
+ a0 = 0.3700794
+ a1 = 0.0
+ a2 = 0.99
+ b0 = 0.0
+ b1 = 0.0
+ dlc = 3e-9
+ dsub = 0.0
+ k3b = 0.0
+ at = 20000.0
+ cf = 0
+ cj = 0.001000266
+ ef = 0.874
+ k1 = 0.5142301
+ k2 = 0.014797844
+ k3 = 0.0
+ em = 30000000.0
+ dwb = 0.0
+ dwg = 0.0
+ js = 3.5e-7
+ ll = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ u0 = 0.04220339
+ pb = 0.6882682
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ dvt0 = 0.0
+ ua = -6.12274e-10
+ dvt1 = 0.0
+ ub = 2.3135539e-18
+ xpart = 1
+ dvt2 = 0.0
+ uc = 1.0876087e-10
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ voff = -0.140578
+ capmod = 3
+ ldif = 9e-8
+ pbswg = 0.6882682
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ jsw = 1.45e-12
+ kt1 = -0.2240464
+ lk2 = 0.0
+ kt2 = -0.030266136
+ lvoff = 0.0
+ eta0 = 5e-5
+ llc = -0.039
+ lln = -1
+ pvag = 0.0
+ etab = -5e-5
+ lu0 = 0.0
+ vsat = 90000.01
+ beta0 = 11.59263
+ nch = 3.9e+17
+ wint = 3e-9
+ lwl = 0.0
+ lwn = 1.0
+ vth0 = 0.4365561
+ leta0 = 1.75e-14
+ mobmod = 1
+ nlx = 0.0
+ rdsw = 170.0
+ lint = 1e-8
+ wmax = 0.000900001
+ lvth0 = 0.0
+ pu0 = 0.0
+ wmin = 1e-5
+ prt = 0
+ lmax = 2.0001e-5
+ delta = 0.01
+ lmin = 1e-5
+ rsh = 6.8
+ tcj = 0.001040287
+ ua1 = 1.224e-9
+ ub1 = -1.1209314e-18
+ uc1 = 1.1643822e-11
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ tpb = 0.001554306
+ tox = 4.08e-9
+ ute = -1.5799998
+ wln = 1.0
+ wu0 = 0.0
+ nfactor = 1.0
+ hdif = 2e-7
+ wwl = 0.0
+ wwn = 1
+ xti = 3
+ mjsw = 0.2003879
+ tcjswg = 0.000645489
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0006999999
+ pdiblcb = 0.01
+ tcjsw = 0.000645489
+ cdsc = 0.0
+ pvoff = 0.0
+ cgdo = 3.665e-10
+ binunit = 2
+ cgso = 3.665e-10
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 7.5e-21
+ pvth0 = 0.0
+ )

.model nch_tt_2 nmos (
+ level = 49
+ wmax = 0.000900001
+ wmin = 1e-5
+ lkt2 = -4.553491e-12
+ lmax = 1e-5
+ lmin = 1.2e-6
+ la0 = -3.496093e-7
+ jsw = 1.45e-12
+ kt1 = -0.2240468
+ lk1 = 1.4908844e-8
+ kt2 = -0.03026568
+ lk2 = -1.111338e-8
+ llc = -0.039
+ lln = -1
+ lketa = -4.320781e-8
+ lu0 = 3.291809e-9
+ lua = -4.643216e-16
+ lub = 7.375677e-25
+ luc = 3.898355e-17
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ xpart = 1
+ pnfactor = 0.0
+ nlx = 0.0
+ hdif = 2e-7
+ wnfactor = 0.0
+ capmod = 3
+ lub1 = 4.527317e-28
+ luc1 = 7.827772e-20
+ nfactor = 1.0
+ pu0 = 0.0
+ mjsw = 0.2003879
+ prt = 0
+ pbswg = 0.6882682
+ lute = -5.743953e-11
+ lvoff = -1.0471328e-8
+ rsh = 6.8
+ tcj = 0.001040287
+ ua1 = 1.224e-9
+ ub1 = -1.1209769e-18
+ uc1 = 1.1635963e-11
+ mobmod = 1
+ beta0 = 11.59263
+ tpb = 0.001554306
+ tox = 4.08e-9
+ lnfactor = 0.0
+ leta0 = 1.75e-14
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0003968181
+ cdsc = 0.0
+ pdiblcb = 0.01
+ lpscbe1 = 262.58185
+ ute = -1.5799941
+ lvsat = -0.006562638
+ cgdo = 3.665e-10
+ wln = 1.0
+ lvth0 = 6.061287e-8
+ wu0 = 0.0
+ wwl = 0.0
+ wwn = 1
+ cgso = 3.665e-10
+ xti = 3
+ delta = 0.01
+ lpdiblc2 = 3.0196912e-9
+ binunit = 2
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ cjsw = 2.040547e-10
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ tnom = 25.0
+ tcjswg = 0.000645489
+ a0 = 0.4051808
+ a1 = 0.0
+ a2 = 0.99
+ b0 = 0.0
+ b1 = 0.0
+ at = 20000.0
+ cf = 0
+ cj = 0.001000266
+ ef = 0.874
+ k1 = 0.5127332
+ k2 = 0.015913647
+ k3 = 0.0
+ em = 30000000.0
+ toxm = 4.08e-9
+ js = 3.5e-7
+ ll = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ u0 = 0.04187289
+ pb = 0.6882682
+ w0 = 0.0
+ pbsw = 0.6882682
+ rd = 0
+ pclm = 0.7736172
+ rs = 0
+ ua = -5.656554e-10
+ ub = 2.2395009e-18
+ uc = 1.0484686e-10
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ tcjsw = 0.000645489
+ version = 3.24
+ pvoff = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 7.5e-21
+ pvth0 = 0.0
+ keta = 0.013601619
+ drout = 0.0
+ tpbsw = 0.001554306
+ dsub = 0.0
+ cjswg = 3.340547e-10
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ mjswg = 0.43879
+ pscbe1 = 173636400.0
+ pscbe2 = 1e-6
+ lcit = 2.6652053e-10
+ wvoff = 0.0
+ voff = -0.1395267
+ ldif = 9e-8
+ ags = 0.02
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ weta0 = 0
+ nqsmod = 0
+ eta0 = 5e-5
+ tpbswg = 0.001554306
+ pvag = 0.0
+ etab = -5e-5
+ cit = -0.00012675911
+ noimod = 2
+ wvsat = 0.0
+ vsat = 90658.91
+ wint = 3e-9
+ dlc = 3e-9
+ lpclm = 2.6277317e-7
+ wvth0 = 0.0
+ vth0 = 0.4304705
+ k3b = 0.0
+ rdsw = 170.0
+ dwb = 0.0
+ dwg = 0.0
+ lint = 1e-8
+ )

.model nch_tt_3 nmos (
+ level = 49
+ beta0 = 11.59263
+ leta0 = 3.813178e-11
+ letab = -3.811428e-11
+ lvsat = -0.0007622857
+ version = 3.24
+ lvth0 = 3.942757e-9
+ delta = 0.01
+ keta = -0.015927497
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ dsub = 0.0
+ pnfactor = 0.0
+ lags = -3.044698e-8
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ tcjswg = 0.000645489
+ wnfactor = 0.0
+ lcit = 3.0262734e-10
+ voff = -0.1621186
+ ldif = 9e-8
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ eta0 = 1.7142866e-5
+ pvag = 0.0
+ etab = -1.7142866e-5
+ vsat = 85658.6
+ tcjsw = 0.000645489
+ lnfactor = 0.0
+ wint = 3e-9
+ vth0 = 0.479324
+ rdsw = 170.0
+ pvoff = 0.0
+ lint = 1e-8
+ wmax = 0.000900001
+ wmin = 1e-5
+ cdscb = 0.0
+ cdscd = 0.0
+ lkt1 = 5.782678e-9
+ lkt2 = 1.5570838e-9
+ peta0 = 7.5e-21
+ lmax = 1.2e-6
+ lpdiblc2 = 1.525682e-9
+ lmin = 5e-7
+ pvth0 = 0.0
+ ags = 0.0462474
+ drout = 0.0
+ tpbsw = 0.001554306
+ cit = -0.00015788565
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ dlc = 3e-9
+ cjswg = 3.340547e-10
+ k3b = 0.0
+ pscbe1 = 400000100.0
+ pscbe2 = 1e-6
+ mjswg = 0.43879
+ dwb = 0.0
+ dwg = 0.0
+ hdif = 2e-7
+ lua1 = -3.0446746e-18
+ lub1 = -1.2004175e-24
+ luc1 = -6.517273e-17
+ wvoff = 0.0
+ mjsw = 0.2003879
+ nqsmod = 0
+ tpbswg = 0.001554306
+ noimod = 2
+ nfactor = 1.0
+ lute = -2.6630502e-7
+ weta0 = 0
+ la0 = 4.581426e-7
+ wvsat = 0.0
+ jsw = 1.45e-12
+ kt1 = -0.2290285
+ lk1 = -7.214246e-9
+ kt2 = -0.031611919
+ lk2 = 1.703151e-9
+ lpclm = 1.5245718e-7
+ wvth0 = 0.0
+ a0 = -0.2911571
+ a1 = 0.0
+ a2 = 0.99
+ b0 = 0.0
+ b1 = 0.0
+ llc = -0.039
+ cdsc = 0.0
+ lln = -1
+ lu0 = 1.0406079e-9
+ at = 20000.0
+ cf = 0
+ cj = 0.001000266
+ ef = 0.874
+ k1 = 0.5318048
+ k2 = 0.004864913
+ k3 = 0.0
+ em = 30000000.0
+ lua = 7.982966e-17
+ lub = -1.5630905e-25
+ luc = -9.669895e-18
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ js = 3.5e-7
+ cgdo = 3.665e-10
+ ll = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0016847569
+ u0 = 0.04381358
+ pb = 0.6882682
+ w0 = 0.0
+ rd = 0
+ nlx = 0.0
+ rs = 0
+ pdiblcb = 0.01
+ ua = -1.0347512e-9
+ ub = 3.0100842e-18
+ uc = 1.4678947e-10
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ cgso = 3.665e-10
+ pu0 = 0.0
+ prt = 0
+ cjsw = 2.040547e-10
+ binunit = 2
+ rsh = 6.8
+ tcj = 0.001040287
+ ua1 = 1.2266247e-9
+ ub1 = -8.574386e-20
+ uc1 = 6.788683e-11
+ lketa = -8.954029e-9
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ tpb = 0.001554306
+ tox = 4.08e-9
+ capmod = 3
+ xpart = 1
+ ute = -1.3504703
+ tnom = 25.0
+ wln = 1.0
+ wu0 = 0.0
+ pbswg = 0.6882682
+ wwl = 0.0
+ wwn = 1
+ xti = 3
+ toxm = 4.08e-9
+ mobmod = 1
+ lvoff = 1.5735258e-8
+ pbsw = 0.6882682
+ pclm = 0.8687172
+ )

.model nch_tt_4 nmos (
+ level = 49
+ lua1 = 8.039099e-19
+ lub1 = 3.824101e-25
+ luc1 = 2.9606131e-17
+ mjsw = 0.2003879
+ lute = 7.030476e-8
+ ags = -0.019916179
+ tcjsw = 0.000645489
+ nfactor = 1.0
+ cdsc = 0.0
+ cit = 0.000271889
+ pvoff = 0.0
+ dlc = 3e-9
+ cgdo = 3.665e-10
+ k3b = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cgso = 3.665e-10
+ peta0 = 7.5e-21
+ pdiblc1 = 1e-6
+ pdiblc2 = -0.00593541
+ pdiblcb = 0.01
+ pvth0 = 0.0
+ drout = 0.0
+ alpha0 = 0.0
+ cjsw = 2.040547e-10
+ alpha1 = 0.448150714
+ tpbsw = 0.001554306
+ la0 = 7.545271e-8
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ pscbe1 = 400000000.0
+ pscbe2 = 1e-6
+ binunit = 2
+ jsw = 1.45e-12
+ kt1 = -0.22715
+ lk1 = 4.899558e-8
+ kt2 = -0.029537767
+ lk2 = -2.3341336e-8
+ cjswg = 3.340547e-10
+ pnfactor = 0.0
+ llc = -0.039
+ lln = -1
+ mjswg = 0.43879
+ lu0 = 1.2517989e-9
+ wnfactor = 0.0
+ lua = -1.0530929e-18
+ lub = 5.559478e-27
+ luc = 4.133919e-18
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ tnom = 25.0
+ nqsmod = 0
+ tpbswg = 0.001554306
+ wvoff = 0.0
+ nlx = 0.0
+ noimod = 2
+ toxm = 4.08e-9
+ pu0 = 0.0
+ weta0 = 0
+ pbsw = 0.6882682
+ pclm = 1.1076791
+ prt = 0
+ wvsat = 0.0
+ lnfactor = 0.0
+ lpclm = 4.253467e-8
+ wvth0 = 0.0
+ rsh = 6.8
+ tcj = 0.001040287
+ ua1 = 1.2182583e-9
+ ub1 = -3.526674e-18
+ uc1 = -1.381542e-10
+ tpb = 0.001554306
+ tox = 4.08e-9
+ ute = -2.0822308
+ version = 3.24
+ wln = 1.0
+ wu0 = 0.0
+ lpdiblc2 = 5.030957e-9
+ wwl = 0.0
+ wwn = 1
+ xti = 3
+ keta = -0.04182327
+ capmod = 3
+ dsub = 0.0
+ lketa = 2.9580252e-9
+ xpart = 1
+ lags = -1.1735286e-11
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ lcit = 1.0493098e-10
+ voff = -0.1245498
+ pbswg = 0.6882682
+ mobmod = 1
+ ldif = 9e-8
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ lvoff = -1.5463618e-9
+ eta0 = -0.0002937502
+ pvag = 0.0
+ etab = 0.0013875004
+ beta0 = 11.59263
+ vsat = 84438.96
+ wint = 3e-9
+ leta0 = 1.8114255999999999e-10
+ vth0 = 0.4752311
+ letab = -6.842502e-10
+ rdsw = 170.0
+ lvsat = -0.00020125005
+ lint = 1e-8
+ lvth0 = 5.825501e-9
+ wmax = 0.000900001
+ wmin = 1e-5
+ lkt1 = 4.918561e-9
+ lkt2 = 6.029743e-10
+ delta = 0.01
+ lmax = 5e-7
+ a0 = 0.5407774
+ a1 = 0.0
+ a2 = 0.99
+ b0 = 0.0
+ b1 = 0.0
+ lmin = 1.8e-7
+ at = 20000.0
+ cf = 0
+ cj = 0.001000266
+ ef = 0.874
+ k1 = 0.4096095
+ k2 = 0.05930946
+ k3 = 0.0
+ em = 30000000.0
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ js = 3.5e-7
+ ll = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ u0 = 0.04335447
+ pb = 0.6882682
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ua = -8.589192e-10
+ ub = 2.6581962e-18
+ uc = 1.1678118e-10
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ tcjswg = 0.000645489
+ hdif = 2e-7
+ )

.model nch_tt_5 nmos (
+ level = 49
+ pu0 = 0.0
+ pscbe1 = 200000030.0
+ pscbe2 = 1e-6
+ tpbsw = 0.001554306
+ prt = 0
+ dsub = 0.0
+ cjswg = 3.340547e-10
+ rsh = 6.8
+ tcj = 0.001040287
+ ua1 = 1.224e-9
+ ub1 = -1.0684574e-18
+ a0 = 0.3702259
+ a1 = 0.0
+ a2 = 0.99
+ uc1 = 2.4230474e-11
+ b0 = 0.0
+ b1 = 0.0
+ mjswg = 0.43879
+ nqsmod = 0
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ tpbswg = 0.001554306
+ at = 20000.0
+ cf = 0
+ cj = 0.001000266
+ ef = 0.874
+ k1 = 0.5102321
+ k2 = 0.016091494
+ k3 = 0.0
+ tpb = 0.001554306
+ noimod = 2
+ em = 30000000.0
+ tox = 4.08e-9
+ js = 3.5e-7
+ wa0 = -1.4643313e-9
+ ll = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ wvoff = 8.907224e-10
+ u0 = 0.0430359
+ pb = 0.6882682
+ w0 = 0.0
+ rd = 0
+ ute = -1.5803809
+ rs = 0
+ ua = -5.885942e-10
+ ub = 2.3329335e-18
+ uc = 1.1057788e-10
+ voff = -0.1406671
+ wk1 = 3.995606e-8
+ wk2 = -1.2928737e-8
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -2e-8
+ ww = 0.0
+ ldif = 9e-8
+ xw = 0.0
+ wln = 1.0
+ wu0 = -8.320099e-9
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ puc1 = -1.4905616e-28
+ weta0 = 0
+ wua = -2.3665659e-16
+ wub = -1.936796e-25
+ wuc = -1.815927e-17
+ wwl = 0.0
+ wwn = 1
+ eta0 = 5e-5
+ xti = 3
+ wvsat = 0.0
+ pvag = 0.0
+ etab = -5e-5
+ vsat = 90000.01
+ wvth0 = 6.876114e-10
+ wint = 3e-9
+ vth0 = 0.4364873
+ rdsw = 170.0
+ wkt1 = -8.215166e-9
+ wkt2 = 1.6245854e-9
+ lint = 1e-8
+ wmax = 1e-5
+ wmin = 1.2e-6
+ lmax = 2.0001e-5
+ lmin = 1e-5
+ capmod = 3
+ xpart = 1
+ wub1 = -5.244247e-25
+ pnfactor = 0.0
+ wuc1 = -1.257911e-16
+ wnfactor = 0.0
+ hdif = 2e-7
+ mobmod = 1
+ wute = 3.808433e-9
+ pbswg = 0.6882682
+ mjsw = 0.2003879
+ lvoff = 0.0
+ beta0 = 11.59263
+ lnfactor = 0.0
+ leta0 = 1.75e-14
+ cdsc = 0.0
+ nfactor = 1.0
+ lvth0 = 0.0
+ cgdo = 3.665e-10
+ cgso = 3.665e-10
+ delta = 0.01
+ dvt0w = 0.0
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0006999999
+ dvt1w = 0.0
+ dvt2w = 0.0
+ pdiblcb = 0.01
+ cjsw = 2.040547e-10
+ tcjswg = 0.000645489
+ ags = 0.02
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ cit = -0.00010000001
+ binunit = 2
+ dlc = 3e-9
+ tnom = 25.0
+ k3b = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ toxm = 4.08e-9
+ pbsw = 0.6882682
+ pclm = 0.8000001
+ tcjsw = 0.000645489
+ pvoff = 0.0
+ jsw = 1.45e-12
+ kt1 = -0.2232244
+ kt2 = -0.030428693
+ lk2 = 0.0
+ llc = -0.039
+ lln = -1
+ lu0 = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ nch = 3.9e+17
+ peta0 = 7.5e-21
+ lwl = 0.0
+ lwn = 1.0
+ nlx = 0.0
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ version = 3.24
+ wketa = -1.0935369e-8
+ pvth0 = 0.0
+ keta = 0.010357677
+ drout = 0.0
+ )

.model nch_tt_6 nmos (
+ level = 49
+ nfactor = 1.0
+ cgso = 3.665e-10
+ capmod = 3
+ cjsw = 2.040547e-10
+ lketa = -4.518989e-8
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0003968181
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ pdiblcb = 0.01
+ lpscbe1 = 262.58185
+ xpart = 1
+ mobmod = 1
+ tnom = 25.0
+ pbswg = 0.6882682
+ binunit = 2
+ toxm = 4.08e-9
+ lvoff = -1.0806052e-8
+ a0 = 0.40626
+ a1 = 0.0
+ a2 = 0.99
+ b0 = 0.0
+ b1 = 0.0
+ pbsw = 0.6882682
+ pclm = 0.7755287
+ at = 20000.0
+ cf = 0
+ cj = 0.001000266
+ ef = 0.874
+ k1 = 0.508509
+ beta0 = 11.59263
+ k2 = 0.01731023
+ k3 = 0.0
+ em = 30000000.0
+ js = 3.5e-7
+ ll = 0.0
+ leta0 = 1.75e-14
+ mj = 0.3595262
+ lw = 0.0
+ u0 = 0.04273027
+ pb = 0.6882682
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ags = 0.02
+ ua = -5.377125e-10
+ ub = 2.2537915e-18
+ uc = 1.0657759e-10
+ lvsat = -0.006753025
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ lvth0 = 6.070609e-8
+ cit = -0.00012675911
+ ppclm = 1.9027247e-13
+ delta = 0.01
+ dlc = 3e-9
+ k3b = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ tcjswg = 0.000645489
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ pkt1 = 4.710912e-15
+ pkt2 = -4.130377e-15
+ keta = 0.014894814
+ version = 3.24
+ dsub = 0.0
+ pnfactor = 0.0
+ la0 = -3.588995e-7
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ wnfactor = 0.0
+ jsw = 1.45e-12
+ lk1 = 1.7161611e-8
+ kt1 = -0.2231775
+ lk2 = -1.2138612e-8
+ kt2 = -0.030469729
+ pketa = 1.9809019e-14
+ llc = -0.039
+ lln = -1
+ lu0 = 3.0440912e-9
+ lcit = 2.6652053e-10
+ voff = -0.1395822
+ lua = -5.067804e-16
+ lub = 7.882536e-25
+ luc = 3.984287e-17
+ nch = 3.9e+17
+ ldif = 9e-8
+ lwl = 0.0
+ lwn = 1.0
+ wpclm = -1.9103656e-8
+ kt1l = 0.0
+ pa0 = 9.284546e-14
+ prwb = 0.0
+ prwg = 0.0
+ pub1 = 4.176128e-31
+ nlx = 0.0
+ puc1 = 7.417578e-23
+ eta0 = 5e-5
+ pk1 = -2.2514154e-14
+ pk2 = 1.0246181e-14
+ pvag = 0.0
+ etab = -5e-5
+ tcjsw = 0.000645489
+ pu0 = 2.4756895e-15
+ vsat = 90678.02
+ lnfactor = 0.0
+ wint = 3e-9
+ pute = -5.708167e-14
+ prt = 0
+ pua = 4.243342e-22
+ pub = -5.065558e-31
+ puc = -8.588134e-24
+ vth0 = 0.4303924
+ rdsw = 170.0
+ pvoff = 3.345241e-15
+ wkt1 = -8.688151e-9
+ wkt2 = 2.0392819e-9
+ rsh = 6.8
+ lint = 1e-8
+ tcj = 0.001040287
+ ua1 = 1.224e-9
+ ub1 = -1.0643074e-18
+ uc1 = 2.4967807e-11
+ wmax = 1e-5
+ wmin = 1.2e-6
+ cdscb = 0.0
+ cdscd = 0.0
+ tpb = 0.001554306
+ peta0 = 7.5e-21
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ tox = 4.08e-9
+ lkt1 = -4.674615e-10
+ lkt2 = 4.087321e-10
+ wa0 = -1.0786144e-8
+ lpdiblc2 = 3.0196912e-9
+ lmax = 1e-5
+ pvsat = 1.9027204e-9
+ ute = -1.5809486
+ pscbe1 = 173636400.0
+ pscbe2 = 1e-6
+ wk1 = 4.221652e-8
+ wk2 = -1.3957471e-8
+ lmin = 1.2e-6
+ wketa = -1.292423e-8
+ pvth0 = -9.316875e-16
+ wln = 1.0
+ drout = 0.0
+ wu0 = -8.568663e-9
+ tpbsw = 0.001554306
+ wua = -2.7926046e-16
+ wub = -1.4282058e-25
+ wuc = -1.7297008e-17
+ wwl = 0.0
+ wwn = 1
+ xti = 3
+ nqsmod = 0
+ tpbswg = 0.001554306
+ cjswg = 3.340547e-10
+ noimod = 2
+ wub1 = -5.663537e-25
+ wuc1 = -1.3323848e-16
+ mjswg = 0.43879
+ hdif = 2e-7
+ wvoff = 5.548539e-10
+ lub1 = -4.133362e-26
+ luc1 = -7.343755e-18
+ wute = 9.539526e-9
+ mjsw = 0.2003879
+ weta0 = 0
+ lute = 5.654154e-9
+ wvsat = -0.00019104627
+ lpclm = 2.4373449e-7
+ wvth0 = 7.811502e-10
+ cdsc = 0.0
+ cgdo = 3.665e-10
+ )

.model nch_tt_7 nmos (
+ level = 49
+ beta0 = 11.59263
+ pvag = 0.0
+ etab = -1.7142869e-5
+ vsat = 85513.59
+ leta0 = 3.813178e-11
+ wint = 3e-9
+ pute = 4.357466e-13
+ letab = -3.811428e-11
+ vth0 = 0.4799949
+ lvsat = -0.0007622865
+ rdsw = 170.0
+ lvth0 = 3.167132e-9
+ wkt1 = -3.681822e-9
+ wkt2 = -1.3190541e-9
+ lint = 1e-8
+ wmax = 1e-5
+ la0 = 4.645035e-7
+ ppclm = 7.258032e-15
+ wmin = 1.2e-6
+ jsw = 1.45e-12
+ lk1 = -1.1179709e-8
+ kt1 = -0.2286601
+ lk2 = 3.431065e-9
+ kt2 = -0.031479932
+ delta = 0.01
+ tcjswg = 0.000645489
+ lkt1 = 5.892387e-9
+ lkt2 = 1.5805686e-9
+ llc = -0.039
+ lln = -1
+ lmax = 1.2e-6
+ lu0 = 9.604713e-10
+ lmin = 5e-7
+ lua = 6.148926e-17
+ lub = -1.2783527e-25
+ luc = -6.505068e-18
+ nch = 3.9e+17
+ dvt0w = 0.0
+ lwl = 0.0
+ lwn = 1.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ pa0 = -6.357063e-14
+ nlx = 0.0
+ pk1 = 3.963084e-14
+ pk2 = -1.7268767e-14
+ pu0 = 8.008865e-16
+ prt = 0
+ pua = 1.8329395e-22
+ pub = -2.8456703e-31
+ puc = -3.16293e-23
+ wua1 = -3.55913e-18
+ wub1 = -1.6132161e-24
+ wuc1 = -1.8047248e-16
+ hdif = 2e-7
+ rsh = 6.8
+ pketa = 9.843987e-15
+ tcj = 0.001040287
+ ua1 = 1.2269809e-9
+ ub1 = 7.567455e-20
+ lua1 = -3.457781e-18
+ uc1 = 8.594492e-11
+ lub1 = -1.3637128e-24
+ luc1 = -7.807721e-17
+ wute = -4.153124e-7
+ mjsw = 0.2003879
+ tpb = 0.001554306
+ tox = 4.08e-9
+ wa0 = 1.2405528e-7
+ wpclm = 1.3866737e-7
+ ute = -1.3089141
+ lute = -3.0990586e-7
+ wk1 = -1.1356744e-8
+ wk2 = 9.762311e-9
+ wln = 1.0
+ tcjsw = 0.000645489
+ wu0 = -7.124867e-9
+ wua = -7.146715e-17
+ wub = -3.341902e-25
+ wuc = 2.5660584e-18
+ wwl = 0.0
+ wwn = 1
+ xti = 3
+ cdsc = 0.0
+ pvoff = -3.013814e-15
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ cgdo = 3.665e-10
+ a0 = -0.3035701
+ a1 = 0.0
+ a2 = 0.99
+ b0 = 0.0
+ b1 = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 7.5e-21
+ at = 20000.0
+ cf = 0
+ cj = 0.001000266
+ pscbe1 = 400000100.0
+ pscbe2 = 1e-6
+ ef = 0.874
+ k1 = 0.5329412
+ k2 = 0.003888095
+ k3 = 0.0
+ em = 30000000.0
+ cgso = 3.665e-10
+ js = 3.5e-7
+ ll = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ u0 = 0.04452649
+ pb = 0.6882682
+ nfactor = 1.0
+ w0 = 0.0
+ rd = 0
+ wketa = -4.333682e-9
+ rs = 0
+ ua = -1.0276002e-9
+ ub = 3.0435232e-18
+ uc = 1.4653272e-10
+ pvth0 = 7.751598e-15
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ drout = 0.0
+ tpbsw = 0.001554306
+ nqsmod = 0
+ cjsw = 2.040547e-10
+ tpbswg = 0.001554306
+ noimod = 2
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ cjswg = 3.340547e-10
+ pnfactor = 0.0
+ mjswg = 0.43879
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0017737894
+ pdiblcb = 0.01
+ wnfactor = 0.0
+ tnom = 25.0
+ wvoff = 6.036798e-9
+ pags = 4.128623e-14
+ toxm = 4.08e-9
+ weta0 = 0
+ ppdiblc2 = 1.0321563e-15
+ binunit = 2
+ pbsw = 0.6882682
+ pclm = 0.8548421
+ wvsat = 0.0014492224
+ wpdiblc2 = -8.897895e-10
+ lpclm = 1.5173094e-7
+ wvth0 = -6.704436e-9
+ lnfactor = 0.0
+ capmod = 3
+ lpdiblc2 = 1.4224044e-9
+ pkt1 = -1.0964308e-15
+ pkt2 = -2.3470743e-16
+ keta = -0.01549387
+ lketa = -9.939018e-9
+ mobmod = 1
+ wags = -3.559157e-8
+ dsub = 0.0
+ version = 3.24
+ xpart = 1
+ ags = 0.04980868
+ lags = -3.457808e-8
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ cit = -0.00015788565
+ pbswg = 0.6882682
+ lcit = 3.0262734e-10
+ voff = -0.1627226
+ ldif = 9e-8
+ dlc = 3e-9
+ k3b = 0.0
+ kt1l = 0.0
+ lvoff = 1.6036822e-8
+ pua1 = 4.128591e-24
+ prwb = 0.0
+ prwg = 0.0
+ pub1 = 1.6319734e-30
+ puc1 = 1.2896722e-22
+ dwb = 0.0
+ dwg = 0.0
+ eta0 = 1.7142869e-5
+ )

.model nch_tt_8 nmos (
+ level = 49
+ pketa = -2.7027957e-15
+ tnom = 25.0
+ pdiblc1 = 1e-6
+ pdiblc2 = -0.006119013
+ pdiblcb = 0.01
+ pags = -1.0838496e-14
+ toxm = 4.08e-9
+ wpclm = 6.656068e-8
+ pcit = 1.4220811e-17
+ pbsw = 0.6882682
+ pclm = 1.1010191
+ tcjsw = 0.000645489
+ binunit = 2
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ pvoff = -9.75415e-16
+ pscbe1 = 400000000.0
+ pscbe2 = 1e-6
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = -1.3746218e-18
+ petab = 1.6959704e-18
+ pvsat = 1.5350395e-12
+ wketa = 2.2941933e-8
+ nqsmod = 0
+ pvth0 = 4.508938e-15
+ tpbswg = 0.001554306
+ drout = 0.0
+ noimod = 2
+ pkt1 = -1.7512235e-15
+ pkt2 = 7.382567e-17
+ keta = -0.04411884
+ tpbsw = 0.001554306
+ wags = 7.772305e-8
+ dsub = 0.0
+ cjswg = 3.340547e-10
+ mjswg = 0.43879
+ lags = 1.0727657e-9
+ wcit = -3.0914837e-11
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ version = 3.24
+ wvoff = 1.6054964e-9
+ lcit = 1.0350804e-10
+ voff = -0.1247105
+ ldif = 9e-8
+ weta0 = 3.0046217e-12
+ kt1l = 0.0
+ pua1 = -1.0901051e-24
+ prwb = 0.0
+ prwg = 0.0
+ pub1 = -4.238914e-31
+ puc1 = -2.7204607e-23
+ wetab = -3.686654e-12
+ wvsat = 0.0014459029
+ eta0 = -0.00029405078
+ pvag = 0.0
+ etab = 0.0013878694
+ lpclm = 3.848953e-8
+ wvth0 = 3.448236e-10
+ vsat = 84294.28
+ wint = 3e-9
+ pute = -1.178615e-13
+ vth0 = 0.4751966
+ rdsw = 170.0
+ capmod = 3
+ wkt1 = -2.2583577e-9
+ wkt2 = -1.9897783e-9
+ lint = 1e-8
+ ags = -0.027693154
+ wmax = 1e-5
+ wmin = 1.2e-6
+ lkt1 = 5.093789e-9
+ lkt2 = 5.955873e-10
+ lmax = 5e-7
+ cit = 0.00027498236
+ lmin = 1.8e-7
+ dlc = 3e-9
+ mobmod = 1
+ k3b = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ a0 = 0.5262308
+ a1 = 0.0
+ a2 = 0.99
+ lketa = 3.228467e-9
+ b0 = 0.0
+ b1 = 0.0
+ at = 20000.0
+ cf = 0
+ cj = 0.001000266
+ ef = 0.874
+ k1 = 0.4007356
+ k2 = 0.0631886
+ k3 = 0.0
+ em = 30000000.0
+ xpart = 1
+ js = 3.5e-7
+ ll = 0.0
+ pnfactor = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ u0 = 0.04384084
+ wua1 = 7.785862e-18
+ pb = 0.6882682
+ wub1 = 2.8560549e-24
+ w0 = 0.0
+ wuc1 = 1.5903152e-16
+ rd = 0
+ rs = 0
+ ua = -9.017296e-10
+ ub = 2.7527719e-18
+ uc = 1.2291169e-10
+ wnfactor = 0.0
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ hdif = 2e-7
+ lua1 = 9.129858e-19
+ lub1 = 4.248247e-25
+ la0 = 8.279508e-8
+ luc1 = 3.232822e-17
+ pbswg = 0.6882682
+ wute = 7.881835e-7
+ mjsw = 0.2003879
+ jsw = 1.45e-12
+ lk1 = 4.963488e-8
+ kt1 = -0.226924
+ lk2 = -2.3847164e-8
+ kt2 = -0.029338669
+ llc = -0.039
+ lvoff = -1.4487617e-9
+ lln = -1
+ lu0 = 1.2758692e-9
+ ppdiblc2 = -2.2121929e-16
+ lute = 8.209799e-8
+ lua = 3.588764e-18
+ lub = 5.910339e-27
+ luc = 4.360599e-18
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ wpdiblc2 = 1.8349379e-9
+ beta0 = 11.59263
+ pa0 = -7.337964e-14
+ lnfactor = 0.0
+ nlx = 0.0
+ leta0 = 1.8128084e-10
+ letab = -6.844199e-10
+ pk1 = -6.389182e-15
+ pk2 = 5.055259e-15
+ lvsat = -0.00020140363
+ cdsc = 0.0
+ pu0 = -2.4055863e-16
+ lvth0 = 5.374336e-9
+ prt = 0
+ pua = -4.639069e-23
+ pub = -3.506499e-33
+ puc = -2.2654354e-24
+ cgdo = 3.665e-10
+ tcjswg = 0.000645489
+ ppclm = 4.042711e-14
+ delta = 0.01
+ cgso = 3.665e-10
+ rsh = 6.8
+ tcj = 0.001040287
+ lpdiblc2 = 5.053093e-9
+ ua1 = 1.2174792e-9
+ ub1 = -3.81245e-18
+ uc1 = -1.540669e-10
+ tpb = 0.001554306
+ tox = 4.08e-9
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ wa0 = 1.4537927e-7
+ nfactor = 1.0
+ ute = -2.1610963
+ cjsw = 2.040547e-10
+ wk1 = 8.868675e-8
+ wk2 = -3.876818e-8
+ wln = 1.0
+ wu0 = -4.860856e-9
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ wua = 4.278473e-16
+ wub = -9.451913e-25
+ wuc = -6.126842e-17
+ wwl = 0.0
+ wwn = 1
+ xti = 3
+ )

.model nch_tt_9 nmos (
+ level = 49
+ cjswg = 3.340547e-10
+ mjswg = 0.43879
+ wub1 = -7.675553e-27
+ wuc1 = -1.4706552e-17
+ hdif = 2e-7
+ wvoff = -8.66569e-10
+ ags = 0.02
+ wute = 3.836007e-8
+ mjsw = 0.2003879
+ weta0 = 0
+ cit = -0.00010000004
+ wvsat = 0.0
+ dlc = 3e-9
+ k3b = 0.0
+ wvth0 = -4.263109e-9
+ dwb = 0.0
+ dwg = 0.0
+ capmod = 3
+ cdsc = 0.0
+ cgdo = 3.665e-10
+ cgso = 3.665e-10
+ mobmod = 1
+ jsw = 1.45e-12
+ kt1 = -0.2313184
+ lk2 = 0.0
+ kt2 = -0.029076951
+ llc = -0.039
+ lln = -1
+ lu0 = 0.0
+ cjsw = 2.040547e-10
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ nlx = 0.0
+ nfactor = 1.0
+ xpart = 1
+ pu0 = 0.0
+ prt = 0
+ tnom = 25.0
+ pbswg = 0.6882682
+ rsh = 6.8
+ tcj = 0.001040287
+ ua1 = 1.224e-9
+ pdiblc1 = 1e-6
+ toxm = 4.08e-9
+ pdiblc2 = 0.0007000003
+ ub1 = -1.5012456e-18
+ lvoff = 0.0
+ uc1 = -6.880516e-11
+ pdiblcb = 0.01
+ pbsw = 0.6882682
+ tpb = 0.001554306
+ pclm = 0.8000001
+ tox = 4.08e-9
+ beta0 = 11.59263
+ wa0 = 7.667051e-8
+ leta0 = 1.75e-14
+ ute = -1.6093186
+ wk1 = -2.074723e-8
+ wk2 = 4.920634e-9
+ tcjswg = 0.000645489
+ wln = 1.0
+ wu0 = 1.0362965e-9
+ lvth0 = 0.0
+ binunit = 2
+ wua = 1.4309126e-16
+ wub = -1.5411778e-25
+ wuc = -1.4141237e-17
+ wwl = 0.0
+ wwn = 1
+ xti = 3
+ delta = 0.01
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ keta = 0.0010152902
+ dsub = 0.0
+ pnfactor = 0.0
+ wnfactor = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ a0 = 0.3047864
+ a1 = 0.0
+ a2 = 0.99
+ b0 = 0.0
+ b1 = 0.0
+ voff = -0.1391954
+ version = 3.24
+ at = 20000.0
+ cf = 0
+ cj = 0.001000266
+ ldif = 9e-8
+ ef = 0.874
+ k1 = 0.5610723
+ k2 = 0.0011422717
+ k3 = 0.0
+ em = 30000000.0
+ kt1l = 0.0
+ js = 3.5e-7
+ prwb = 0.0
+ ll = 0.0
+ prwg = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ u0 = 0.03519972
+ pb = 0.6882682
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ua = -9.066409e-10
+ ub = 2.2997995e-18
+ uc = 1.072127e-10
+ eta0 = 5e-5
+ wl = 0.0
+ tcjsw = 0.000645489
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -2e-8
+ ww = 0.0
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ xw = 0.0
+ pvag = 0.0
+ etab = -5e-5
+ lnfactor = 0.0
+ vsat = 90000.01
+ wint = 3e-9
+ pscbe1 = 200000030.0
+ pscbe2 = 1e-6
+ vth0 = 0.4406337
+ pvoff = 0.0
+ rdsw = 170.0
+ wkt1 = 1.4490446e-9
+ wkt2 = 1.0605161e-11
+ lint = 1e-8
+ wmax = 1.2e-6
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 7.5e-21
+ wmin = 5e-7
+ nqsmod = 0
+ tpbswg = 0.001554306
+ noimod = 2
+ lmax = 2.0001e-5
+ wketa = 2.1944087e-10
+ pvth0 = 0.0
+ lmin = 1e-5
+ drout = 0.0
+ tpbsw = 0.001554306
+ )

.model nch_tt_10 nmos (
+ level = 49
+ lute = -1.2190513e-8
+ nqsmod = 0
+ tpbswg = 0.001554306
+ noimod = 2
+ cdsc = 0.0
+ cgdo = 3.665e-10
+ nfactor = 1.0
+ lketa = -2.8027248e-8
+ cgso = 3.665e-10
+ xpart = 1
+ cjsw = 2.040547e-10
+ pbswg = 0.6882682
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0003968185
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ pdiblcb = 0.01
+ lpscbe1 = 262.58185
+ lvoff = -3.602222e-9
+ capmod = 3
+ beta0 = 11.59263
+ tnom = 25.0
+ leta0 = 1.75e-14
+ binunit = 2
+ lvsat = -0.006201102
+ toxm = 4.08e-9
+ lvth0 = 6.592048e-8
+ pcit = 4.302753e-19
+ pbsw = 0.6882682
+ pclm = 0.7699873
+ ppclm = 1.243718e-13
+ mobmod = 1
+ delta = 0.01
+ ags = 0.02
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ cit = -0.00012672294
+ dlc = 3e-9
+ k3b = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ pnfactor = 0.0
+ pkt1 = 7.833639e-15
+ pkt2 = 9.747044e-16
+ keta = 0.00382927
+ wnfactor = 0.0
+ pketa = -6.831802e-16
+ version = 3.24
+ dsub = 0.0
+ wpclm = -1.2487239e-8
+ wcit = -4.317371e-14
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ la0 = -1.9725388e-7
+ tcjsw = 0.000645489
+ jsw = 1.45e-12
+ tcjswg = 0.000645489
+ lk1 = 1.0512358e-8
+ kt1 = -0.2310088
+ lk2 = -5.410051e-9
+ kt2 = -0.028688708
+ lcit = 2.6616018e-10
+ llc = -0.039
+ lln = -1
+ voff = -0.1388337
+ lu0 = 3.705752e-9
+ lnfactor = 0.0
+ ldif = 9e-8
+ lua = -1.9124487e-16
+ lub = 4.117038e-25
+ luc = 4.038815e-17
+ nch = 3.9e+17
+ pvoff = -5.256132e-15
+ lwl = 0.0
+ lwn = 1.0
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ pub1 = -1.8996434e-32
+ puc1 = 1.3569954e-23
+ pa0 = -1.0015934e-13
+ nlx = 0.0
+ eta0 = 5e-5
+ pk1 = -1.457495e-14
+ pk2 = 2.2122807e-15
+ pvag = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ etab = -5e-5
+ peta0 = 7.5e-21
+ vsat = 90622.61
+ wint = 3e-9
+ pu0 = 1.6856667e-15
+ pute = -3.577514e-14
+ pvsat = 1.2437262e-9
+ vth0 = 0.4340151
+ prt = 0
+ pua = 4.758471e-23
+ pub = -5.695533e-32
+ puc = -9.239189e-24
+ lpdiblc2 = 3.0196912e-9
+ wketa = 2.8803285e-10
+ rdsw = 170.0
+ pvth0 = -7.157672e-15
+ wkt1 = 6.625341e-10
+ wkt2 = -8.725676e-11
+ drout = 0.0
+ lint = 1e-8
+ rsh = 6.8
+ tpbsw = 0.001554306
+ wmax = 1.2e-6
+ tcj = 0.001040287
+ ua1 = 1.224e-9
+ ub1 = -1.5338095e-18
+ uc1 = -7.316409e-11
+ wmin = 5e-7
+ lkt1 = -3.0828107e-9
+ lkt2 = -3.866881e-9
+ tpb = 0.001554306
+ tox = 4.08e-9
+ cjswg = 3.340547e-10
+ lmax = 1e-5
+ wa0 = 8.672666e-8
+ lmin = 1.2e-6
+ ute = -1.6080947
+ mjswg = 0.43879
+ wk1 = -1.9283881e-8
+ wk2 = 4.698517e-9
+ wln = 1.0
+ wu0 = 8.670528e-10
+ wvoff = -3.388445e-10
+ wua = 1.3831368e-16
+ wub = -1.4839938e-25
+ wuc = -1.3213606e-17
+ wwl = 0.0
+ wwn = 1
+ xti = 3
+ a0 = 0.324591
+ a1 = 0.0
+ a2 = 0.99
+ b0 = 0.0
+ b1 = 0.0
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ wub1 = -5.768295e-27
+ wuc1 = -1.6068998e-17
+ weta0 = 0
+ at = 20000.0
+ cf = 0
+ cj = 0.001000266
+ ef = 0.874
+ k1 = 0.5600169
+ k2 = 0.0016854487
+ k3 = 0.0
+ em = 30000000.0
+ hdif = 2e-7
+ wvsat = -0.00012487893
+ js = 3.5e-7
+ pscbe1 = 173636400.0
+ pscbe2 = 1e-6
+ ll = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ u0 = 0.03482766
+ pb = 0.6882682
+ lub1 = 3.243357e-25
+ lpclm = 2.9892766e-7
+ wvth0 = -3.544466e-9
+ luc1 = 4.341489e-17
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ wute = 4.195195e-8
+ ua = -8.874397e-10
+ ub = 2.2584638e-18
+ uc = 1.0315766e-10
+ mjsw = 0.2003879
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ )

.model nch_tt_11 nmos (
+ level = 49
+ lvoff = 1.116323e-8
+ wcit = 5.431231e-13
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ ags = 0.02
+ beta0 = 11.59263
+ leta0 = 3.81318e-11
+ lcit = 3.0283653e-10
+ cit = -0.0001583405
+ letab = -3.81143e-11
+ voff = -0.1515625
+ ldif = 9e-8
+ lvsat = -0.0007659488
+ dlc = 3e-9
+ kt1l = 0.0
+ mobmod = 1
+ prwb = 0.0
+ lvth0 = 1.0109751e-8
+ prwg = 0.0
+ pub1 = -5.874811e-31
+ puc1 = -3.67348e-23
+ a0 = -0.1914371
+ a1 = 0.0
+ a2 = 0.99
+ k3b = 0.0
+ b0 = 0.0
+ b1 = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ eta0 = 1.7142847e-5
+ at = 20000.0
+ cf = 0
+ cj = 0.001000266
+ ef = 0.874
+ k1 = 0.5552615
+ ppclm = 7.308824e-14
+ k2 = 0.003544799
+ k3 = 0.0
+ em = 30000000.0
+ pvag = 0.0
+ etab = -1.7142847e-5
+ delta = 0.01
+ js = 3.5e-7
+ vsat = 85937.13
+ ll = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ u0 = 0.03581186
+ pb = 0.6882682
+ wint = 3e-9
+ pute = -2.0303331e-13
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ua = -1.3333591e-9
+ ub = 2.969086e-18
+ uc = 1.6160392e-10
+ vth0 = 0.4821278
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ rdsw = 170.0
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ wkt1 = 1.1898274e-8
+ wkt2 = 2.0987987e-9
+ lint = 1e-8
+ wmax = 1.2e-6
+ la0 = 4.013388e-7
+ wmin = 5e-7
+ lkt1 = 9.329063e-9
+ lkt2 = 2.691467e-9
+ jsw = 1.45e-12
+ lk1 = 1.6028618e-8
+ kt1 = -0.2417087
+ lk2 = -7.566896e-9
+ kt2 = -0.03434246
+ lmax = 1.2e-6
+ llc = -0.039
+ lln = -1
+ lu0 = 2.5640821e-9
+ lmin = 5e-7
+ lua = 3.260216e-16
+ lub = -4.12618e-25
+ luc = -2.7409531e-17
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ pketa = 1.4501565e-15
+ pa0 = 1.1848049e-14
+ nlx = 0.0
+ pk1 = 7.144098e-15
+ pk2 = -4.137203e-15
+ pu0 = -1.1138246e-15
+ wpclm = 3.172275e-8
+ wub1 = 4.843047e-25
+ prt = 0
+ wuc1 = 2.7297169e-17
+ pua = -1.3255767e-22
+ pub = 5.546348e-32
+ puc = -6.669366e-24
+ tcjswg = 0.000645489
+ hdif = 2e-7
+ tcjsw = 0.000645489
+ rsh = 6.8
+ lub1 = 4.951269e-25
+ luc1 = 6.070172e-17
+ tcj = 0.001040287
+ ua1 = 1.224e-9
+ ub1 = -1.6810433e-18
+ uc1 = -8.806652e-11
+ wute = 1.8614003e-7
+ mjsw = 0.2003879
+ pvoff = 2.8052535e-15
+ tpb = 0.001554306
+ tox = 4.08e-9
+ wa0 = -9.831444e-9
+ lute = 2.2508574e-7
+ ute = -1.8126432
+ wk1 = -3.80072e-8
+ wk2 = 1.0172209e-8
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 7.5e-21
+ wln = 1.0
+ wu0 = 3.280407e-9
+ wua = 2.9360883e-16
+ pvsat = 4.380818e-12
+ wub = -2.4531215e-25
+ wuc = -1.542897e-17
+ wwl = 0.0
+ wwn = 1
+ cdsc = 0.0
+ wketa = -1.5510503e-9
+ pvth0 = -5.378882e-16
+ xti = 3
+ drout = 0.0
+ cgdo = 3.665e-10
+ tpbsw = 0.001554306
+ cgso = 3.665e-10
+ cjswg = 3.340547e-10
+ nfactor = 1.0
+ mjswg = 0.43879
+ pnfactor = 0.0
+ cjsw = 2.040547e-10
+ wnfactor = 0.0
+ wvoff = -7.288315e-9
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ weta0 = 0
+ pscbe1 = 400000100.0
+ pscbe2 = 1e-6
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0011219129
+ pdiblcb = 0.01
+ wvsat = 0.0009435224
+ ppdiblc2 = 1.2928064e-16
+ tnom = 25.0
+ lpclm = 9.659676e-8
+ wvth0 = -9.251178e-9
+ wpdiblc2 = -1.1144895e-10
+ lnfactor = 0.0
+ nqsmod = 0
+ tpbswg = 0.001554306
+ toxm = 4.08e-9
+ noimod = 2
+ pcit = -2.4980728e-19
+ binunit = 2
+ pbsw = 0.6882682
+ pclm = 0.9444105
+ lpdiblc2 = 2.1785818e-9
+ lketa = -2.9090079e-9
+ xpart = 1
+ pkt1 = -5.199821e-15
+ pkt2 = -1.5611203e-15
+ keta = -0.017824383
+ pbswg = 0.6882682
+ dsub = 0.0
+ capmod = 3
+ version = 3.24
+ )

.model nch_tt_12 nmos (
+ level = 49
+ tpb = 0.001554306
+ tox = 4.08e-9
+ wa0 = 1.7605426e-7
+ pketa = -7.367843e-16
+ cjsw = 2.040547e-10
+ nfactor = 1.0
+ ute = -1.2073984
+ wk1 = -1.7855582e-8
+ wk2 = 1.6966123e-9
+ tcjswg = 0.000645489
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ wln = 1.0
+ wu0 = -4.268465e-11
+ wpclm = 1.9327061e-7
+ wua = -1.9101984e-17
+ wub = -5.11281e-26
+ wuc = -9.012729e-18
+ wwl = 0.0
+ wwn = 1
+ xti = 3
+ tcjsw = 0.000645489
+ tnom = 25.0
+ pdiblc1 = 1e-6
+ pdiblc2 = -0.00401322
+ pags = 1.8981756e-15
+ pdiblcb = 0.01
+ pvoff = -2.2207474e-15
+ toxm = 4.08e-9
+ pcit = -1.4232223e-17
+ pbsw = 0.6882682
+ pclm = 0.9948969
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = -1.1364491000000001e-17
+ petab = 1.3954016e-17
+ binunit = 2
+ pvsat = 1.606088e-11
+ wketa = 3.203169e-9
+ pvth0 = 2.716016e-15
+ drout = 0.0
+ tpbsw = 0.001554306
+ a0 = 0.5005398
+ a1 = 0.0
+ a2 = 0.99
+ b0 = 0.0
+ b1 = 0.0
+ at = 20000.0
+ cf = 0
+ cj = 0.001000266
+ ef = 0.874
+ k1 = 0.489967
+ k2 = 0.029298484
+ k3 = 0.0
+ em = 30000000.0
+ js = 3.5e-7
+ cjswg = 3.340547e-10
+ ll = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ u0 = 0.03980552
+ pb = 0.6882682
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ua = -5.274002e-10
+ ub = 2.0039751e-18
+ uc = 7.914647e-11
+ mjswg = 0.43879
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ pkt1 = 2.3961372e-15
+ pkt2 = 8.832021e-16
+ keta = -0.027587207
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ wvoff = 3.637774e-9
+ wags = -4.12647e-9
+ dsub = 0.0
+ pscbe1 = 400000000.0
+ pscbe2 = 1e-6
+ weta0 = 2.4721704e-11
+ lags = -9.594464e-9
+ wetab = -3.0334849e-11
+ wcit = 3.093965e-11
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ wvsat = 0.000918131
+ version = 3.24
+ nqsmod = 0
+ lpclm = 7.337301e-8
+ wvth0 = -1.6324883e-8
+ tpbswg = 0.001554306
+ noimod = 2
+ lcit = 1.2733804e-10
+ voff = -0.1264125
+ ldif = 9e-8
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ pub1 = 1.6165291e-31
+ puc1 = 2.0250814e-23
+ eta0 = -0.00031223928
+ pvag = 0.0
+ etab = 0.0014101875
+ vsat = 84736.3
+ wint = 3e-9
+ pute = 4.383575e-14
+ vth0 = 0.4891579
+ rdsw = 170.0
+ wkt1 = -4.614678e-9
+ wkt2 = -3.214946e-9
+ lint = 1e-8
+ wmax = 1.2e-6
+ ags = 0.04085753
+ lketa = 1.5818911e-9
+ wmin = 5e-7
+ lkt1 = 1.6202869e-9
+ lkt2 = -8.228257e-11
+ lmax = 5e-7
+ xpart = 1
+ cit = 0.00022317801
+ lmin = 1.8e-7
+ pnfactor = 0.0
+ dlc = 3e-9
+ wnfactor = 0.0
+ k3b = 0.0
+ capmod = 3
+ dwb = 0.0
+ dwg = 0.0
+ pbswg = 0.6882682
+ lvoff = -4.057695e-10
+ wub1 = -1.1442477e-24
+ wuc1 = -9.658459e-17
+ ppdiblc2 = 3.905237e-16
+ hdif = 2e-7
+ beta0 = 11.59263
+ wpdiblc2 = -6.793707e-10
+ lub1 = -6.558089e-26
+ leta0 = 1.8964756e-10
+ luc1 = -7.416688e-18
+ wute = -3.505318e-7
+ mobmod = 1
+ la0 = 8.302936e-8
+ letab = -6.946862e-10
+ lnfactor = 0.0
+ mjsw = 0.2003879
+ lvsat = -0.00021356932
+ jsw = 1.45e-12
+ lk1 = 4.606408e-8
+ kt1 = -0.2249505
+ lk2 = -1.9413593e-8
+ kt2 = -0.028312566
+ lvth0 = 6.875945e-9
+ llc = -0.039
+ lln = -1
+ lute = -5.332685e-8
+ lu0 = 7.269945e-10
+ lua = -4.471944e-17
+ lub = 3.1333025e-26
+ luc = 1.0520902e-17
+ ppclm = -1.2237712e-15
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ delta = 0.01
+ pa0 = -7.365936e-14
+ nlx = 0.0
+ lpdiblc2 = 4.540744e-9
+ cdsc = 0.0
+ pk1 = -2.1256446e-15
+ pk2 = -2.3842633e-16
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ pu0 = 4.147977e-16
+ cgdo = 3.665e-10
+ prt = 0
+ pua = 1.1289303e-23
+ pub = -3.386118e-32
+ puc = -9.620837e-24
+ cgso = 3.665e-10
+ rsh = 6.8
+ tcj = 0.001040287
+ ua1 = 1.224e-9
+ ub1 = -4.621132e-19
+ uc1 = 6.001696e-11
+ )

.model nch_tt_13 nmos (
+ level = 49
+ drout = 0.0
+ wkt1 = 5.128653e-9
+ wkt2 = 3.532295e-9
+ tpbsw = 0.001554306
+ lint = 1e-8
+ wmax = 5e-7
+ wmin = 2.2e-7
+ cjswg = 3.340547e-10
+ lmax = 2.0001e-5
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ mjswg = 0.43879
+ lmin = 1e-5
+ pscbe1 = 200000030.0
+ pscbe2 = 1e-6
+ wvoff = -1.7276782e-9
+ weta0 = 0
+ nqsmod = 0
+ wub1 = -4.432931e-26
+ wuc1 = -1.7086574e-17
+ tpbswg = 0.001554306
+ wvsat = 0.0
+ noimod = 2
+ hdif = 2e-7
+ wvth0 = -1.5455745e-8
+ ags = 0.02
+ wute = 2.5547985e-8
+ mjsw = 0.2003879
+ cit = -9.999998e-5
+ dlc = 3e-9
+ k3b = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ cdsc = 0.0
+ cgdo = 3.665e-10
+ cgso = 3.665e-10
+ xpart = 1
+ jsw = 1.45e-12
+ capmod = 3
+ kt1 = -0.238767
+ lk2 = 0.0
+ kt2 = -0.03620588
+ llc = -0.039
+ cjsw = 2.040547e-10
+ lln = -1
+ a0 = 0.352982
+ a1 = 0.0
+ a2 = 0.99
+ lu0 = 0.0
+ b0 = 0.0
+ b1 = 0.0
+ pbswg = 0.6882682
+ nch = 3.9e+17
+ at = 20000.0
+ cf = 0
+ cj = 0.001000266
+ lwl = 0.0
+ lwn = 1.0
+ ef = 0.874
+ k1 = 0.5220979
+ k2 = 0.016542569
+ k3 = 0.0
+ em = 30000000.0
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ nfactor = 1.0
+ js = 3.5e-7
+ ll = 0.0
+ nlx = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ lvoff = 0.0
+ u0 = 0.03533742
+ pb = 0.6882682
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ua = -5.860608e-10
+ ub = 1.7266676e-18
+ uc = 7.252202e-11
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ mobmod = 1
+ beta0 = 11.59263
+ pu0 = 0.0
+ tnom = 25.0
+ leta0 = 1.75e-14
+ prt = 0
+ toxm = 4.08e-9
+ rsh = 6.8
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0006999999
+ lvth0 = 0.0
+ tcj = 0.001040287
+ ua1 = 1.224e-9
+ ub1 = -1.4270478e-18
+ uc1 = -6.39873e-11
+ pdiblcb = 0.01
+ pbsw = 0.6882682
+ pclm = 0.7999999
+ tpb = 0.001554306
+ tox = 4.08e-9
+ delta = 0.01
+ wa0 = 5.286186e-8
+ ute = -1.5833832
+ wk1 = -1.4938487e-9
+ wk2 = -2.6871128e-9
+ dvt0w = 0.0
+ dvt1w = 0.0
+ wln = 1.0
+ dvt2w = 0.0
+ wu0 = 9.682726e-10
+ binunit = 2
+ wua = -1.5275344e-17
+ wub = 1.2900942e-25
+ wuc = 2.9959555e-18
+ wwl = 0.0
+ wwn = 1
+ xti = 3
+ pnfactor = 0.0
+ keta = 0.002064252
+ tcjswg = 0.000645489
+ wnfactor = 0.0
+ dsub = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ tcjsw = 0.000645489
+ lnfactor = 0.0
+ voff = -0.1374522
+ version = 3.24
+ pvoff = 0.0
+ ldif = 9e-8
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ eta0 = 5e-5
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 7.5e-21
+ pvag = 0.0
+ etab = -5e-5
+ vsat = 89999.99
+ wint = 3e-9
+ vth0 = 0.4632908
+ wketa = -2.9874625e-10
+ pvth0 = 0.0
+ rdsw = 170.0
+ )

.model nch_tt_14 nmos (
+ level = 49
+ la0 = -2.4964379e-7
+ pcit = 1.5653096e-18
+ pbsw = 0.6882682
+ pclm = 0.7606163
+ jsw = 1.45e-12
+ lk1 = -6.331243e-8
+ kt1 = -0.2407974
+ lk2 = 2.0798732e-8
+ kt2 = -0.03589625
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0003968183
+ pdiblcb = 0.01
+ lpscbe1 = 262.58182
+ llc = -0.039
+ lln = -1
+ lu0 = 9.894555e-9
+ lpdiblc2 = 3.0196909e-9
+ lua = -1.2876533e-16
+ lub = 7.836163e-25
+ luc = 7.064626e-17
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ pa0 = -7.427873e-14
+ nlx = 0.0
+ pk1 = 2.1894499e-14
+ pk2 = -1.0734859e-14
+ lketa = -3.0377027e-8
+ binunit = 2
+ pu0 = -1.3716021e-15
+ capmod = 3
+ prt = 0
+ pua = 1.6719826e-23
+ pub = -2.4068014e-31
+ xpart = 1
+ puc = -2.4186704e-23
+ pkt1 = -3.679308e-15
+ pkt2 = 5.879336e-16
+ rsh = 6.8
+ keta = 0.005114151
+ tcj = 0.001040287
+ ua1 = 1.224e-9
+ ub1 = -1.4513121e-18
+ uc1 = -6.991786e-11
+ pbswg = 0.6882682
+ tpb = 0.001554306
+ tox = 4.08e-9
+ dsub = 0.0
+ wa0 = 6.031956e-8
+ lvoff = -1.9727372e-8
+ mobmod = 1
+ ute = -1.5785241
+ wk1 = -3.692092e-9
+ wk2 = -1.6093152e-9
+ wcit = -1.5715551e-13
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ wln = 1.0
+ beta0 = 11.59263
+ wu0 = 1.1059835e-9
+ wua = -1.6954039e-17
+ wub = 1.5317406e-25
+ wuc = 5.42434e-18
+ leta0 = 1.75e-14
+ wwl = 0.0
+ wwn = 1
+ lcit = 2.6386249e-10
+ xti = 3
+ voff = -0.1354716
+ lvsat = -0.005267757
+ ldif = 9e-8
+ lvth0 = 5.627824e-8
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ pub1 = 2.1839324e-32
+ puc1 = 5.837128e-24
+ version = 3.24
+ ppclm = 7.826515e-14
+ eta0 = 5e-5
+ delta = 0.01
+ pvag = 0.0
+ etab = -5e-5
+ vsat = 90528.88
+ wint = 3e-9
+ pute = -1.7889165e-14
+ vth0 = 0.4576404
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ rdsw = 170.0
+ wkt1 = 5.498062e-9
+ wkt2 = 3.473265e-9
+ lint = 1e-8
+ wmax = 5e-7
+ wmin = 2.2e-7
+ lkt1 = 2.0222748e-8
+ lkt2 = -3.0839447e-9
+ lmax = 1e-5
+ tcjswg = 0.000645489
+ lmin = 1.2e-6
+ pketa = 4.776125e-16
+ wpclm = -7.857923e-9
+ wub1 = -4.652201e-26
+ wuc1 = -1.7672629e-17
+ tcjsw = 0.000645489
+ hdif = 2e-7
+ lub1 = 2.4167225e-25
+ a0 = 0.3780467
+ a1 = 0.0
+ a2 = 0.99
+ luc1 = 5.906839e-17
+ b0 = 0.0
+ b1 = 0.0
+ wute = 2.7344081e-8
+ mjsw = 0.2003879
+ at = 20000.0
+ pvoff = 2.7096929e-15
+ cf = 0
+ cj = 0.001000266
+ ef = 0.874
+ k1 = 0.5284545
+ k2 = 0.014454342
+ k3 = 0.0
+ em = 30000000.0
+ js = 3.5e-7
+ ll = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ u0 = 0.034344
+ pb = 0.6882682
+ w0 = 0.0
+ rd = 0
+ lute = -4.839696e-8
+ rs = 0
+ ua = -5.731325e-10
+ ub = 1.6479914e-18
+ uc = 6.542903e-11
+ cdscb = 0.0
+ cdscd = 0.0
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -2e-8
+ ww = 0.0
+ peta0 = 7.5e-21
+ xw = 0.0
+ pvsat = 7.826533e-10
+ wketa = -3.466991e-10
+ pvth0 = -2.3944025e-15
+ cdsc = 0.0
+ drout = 0.0
+ tpbsw = 0.001554306
+ cgdo = 3.665e-10
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ cgso = 3.665e-10
+ cjswg = 3.340547e-10
+ pscbe1 = 173636400.0
+ pscbe2 = 1e-6
+ mjswg = 0.43879
+ ags = 0.02
+ pnfactor = 0.0
+ wnfactor = 0.0
+ wvoff = -1.9997353e-9
+ cjsw = 2.040547e-10
+ cit = -0.00012649217
+ nqsmod = 0
+ dlc = 3e-9
+ tpbswg = 0.001554306
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ noimod = 2
+ k3b = 0.0
+ weta0 = 0
+ dwb = 0.0
+ dwg = 0.0
+ wvsat = -7.857954e-5
+ nfactor = 1.0
+ lpclm = 3.92261e-7
+ wvth0 = -1.5215344e-8
+ tnom = 25.0
+ lnfactor = 0.0
+ toxm = 4.08e-9
+ )

.model nch_tt_15 nmos (
+ level = 49
+ wub1 = -1.0574451e-25
+ wuc1 = -4.040928e-17
+ ppdiblc2 = 4.703685e-16
+ beta0 = 11.59263
+ hdif = 2e-7
+ wpdiblc2 = -4.054901e-10
+ leta0 = 3.813178e-11
+ lub1 = -8.773805e-25
+ luc1 = -7.886598e-17
+ letab = -3.811428e-11
+ lnfactor = 0.0
+ wute = 1.9757099e-8
+ lvsat = -0.0007893788
+ mjsw = 0.2003879
+ lvth0 = 8.859259e-9
+ lute = -1.6751561e-7
+ ppclm = 4.863229e-14
+ delta = 0.01
+ lpdiblc2 = 1.4881204e-9
+ dvt0w = 0.0
+ cdsc = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ cgdo = 3.665e-10
+ tcjswg = 0.000645489
+ cgso = 3.665e-10
+ pketa = 3.1429577e-15
+ cjsw = 2.040547e-10
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ wpclm = 1.7687656e-8
+ tcjsw = 0.000645489
+ tnom = 25.0
+ nfactor = 1.0
+ pvoff = -1.3837542e-15
+ toxm = 4.08e-9
+ ags = 0.02
+ pcit = -9.088336e-19
+ pbsw = 0.6882682
+ pclm = 0.9728217
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 7.5e-21
+ pvsat = 1.5955267e-11
+ cit = -0.00016124053
+ wketa = -2.6444102e-9
+ pvth0 = 7.985465e-17
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0017171376
+ dlc = 3e-9
+ drout = 0.0
+ pdiblcb = 0.01
+ k3b = 0.0
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ tpbsw = 0.001554306
+ dwb = 0.0
+ dwg = 0.0
+ pscbe1 = 400000100.0
+ pscbe2 = 1e-6
+ cjswg = 3.340547e-10
+ mjswg = 0.43879
+ binunit = 2
+ pkt1 = -1.1651986e-14
+ pkt2 = -1.4582807e-15
+ keta = -0.015611105
+ nqsmod = 0
+ wvoff = 1.529098e-9
+ tpbswg = 0.001554306
+ la0 = 2.7901473e-7
+ noimod = 2
+ jsw = 1.45e-12
+ dsub = 0.0
+ lk1 = 6.936774e-8
+ kt1 = -0.2426658
+ lk2 = -3.1528607e-8
+ kt2 = -0.04069558
+ llc = -0.039
+ lln = -1
+ weta0 = 0
+ lu0 = -1.7446106e-9
+ lua = 6.135559e-17
+ lub = -2.9489129e-25
+ luc = -2.7169401e-17
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ wvsat = 0.0005823669
+ wcit = 1.975718e-12
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ pa0 = 7.227613e-14
+ nlx = 0.0
+ lpclm = 1.4610272e-7
+ wvth0 = -1.7348324e-8
+ pk1 = -1.920543e-14
+ pk2 = 7.699883e-15
+ lcit = 3.0417063e-10
+ voff = -0.1694116
+ pu0 = 1.0146696e-15
+ ldif = 9e-8
+ prt = 0
+ pua = -1.8126578e-24
+ pub = -2.6935e-33
+ puc = -6.78799e-24
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ pub1 = 9.053745e-32
+ puc1 = 3.221165e-23
+ eta0 = 1.7142866e-5
+ rsh = 6.8
+ pvag = 0.0
+ etab = -1.7142866e-5
+ tcj = 0.001040287
+ ua1 = 1.224e-9
+ ub1 = -4.866116e-19
+ uc1 = 4.899104e-11
+ vsat = 86668.21
+ version = 3.24
+ a0 = -0.07769345
+ wint = 3e-9
+ a1 = 0.0
+ a2 = 0.99
+ pute = -9.088265e-15
+ b0 = 0.0
+ b1 = 0.0
+ tpb = 0.001554306
+ vth0 = 0.4985188
+ tox = 4.08e-9
+ at = 20000.0
+ cf = 0
+ cj = 0.001000266
+ ef = 0.874
+ k1 = 0.4140751
+ k2 = 0.05956412
+ k3 = 0.0
+ rdsw = 170.0
+ wa0 = -6.602082e-8
+ em = 30000000.0
+ js = 3.5e-7
+ wkt1 = 1.2371058e-8
+ wkt2 = 5.237243e-9
+ ute = -1.4758356
+ ll = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ lint = 1e-8
+ u0 = 0.04437776
+ pb = 0.6882682
+ wk1 = 3.173889e-8
+ wk2 = -1.7501334e-8
+ w0 = 0.0
+ rd = 0
+ wmax = 5e-7
+ lketa = -6.33573e-9
+ capmod = 3
+ rs = 0
+ ua = -7.370299e-10
+ ub = 2.5777392e-18
+ uc = 1.4975288e-10
+ wln = 1.0
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -2e-8
+ ww = 0.0
+ wmin = 2.2e-7
+ wu0 = -9.511471e-10
+ xw = 0.0
+ lkt1 = 2.2390124e-8
+ wua = -9.777621e-19
+ lkt2 = 2.4832894e-9
+ wub = -5.19868e-26
+ wuc = -9.57455e-18
+ xpart = 1
+ wwl = 0.0
+ wwn = 1
+ lmax = 1.2e-6
+ xti = 3
+ lmin = 5e-7
+ pnfactor = 0.0
+ wnfactor = 0.0
+ pbswg = 0.6882682
+ mobmod = 1
+ lvoff = 1.9643004e-8
+ )

.model nch_tt_16 nmos (
+ level = 49
+ at = 20000.0
+ cf = 0
+ cj = 0.001000266
+ ef = 0.874
+ k1 = 0.4942783
+ k2 = 0.023518253
+ k3 = 0.0
+ em = 30000000.0
+ pketa = -1.9609824e-16
+ pkt1 = 3.435378e-15
+ pkt2 = -8.505888e-17
+ wnfactor = 0.0
+ keta = -0.030443965
+ js = 3.5e-7
+ ll = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ ags = 0.0548038
+ u0 = 0.0371035
+ pb = 0.6882682
+ w0 = 0.0
+ binunit = 2
+ rd = 0
+ rs = 0
+ ua = -6.614348e-10
+ ub = 2.1301375e-18
+ uc = 1.2526492e-10
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ wags = -1.1015922e-8
+ xl = -2e-8
+ ww = 0.0
+ dsub = 0.0
+ xw = 0.0
+ wpclm = 1.2379924e-7
+ cit = 0.00029138371
+ lags = -1.6009743e-8
+ dlc = 3e-9
+ wcit = -2.7539906e-12
+ ppdiblc2 = -1.1422951e-16
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ tcjsw = 0.000645489
+ k3b = 0.0
+ wpdiblc2 = 8.65375e-10
+ dwb = 0.0
+ dwg = 0.0
+ lnfactor = 0.0
+ lcit = 9.596344e-11
+ pvoff = -4.969337e-16
+ voff = -0.1182414
+ ldif = 9e-8
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ pub1 = -3.181536e-32
+ puc1 = -1.1609298e-23
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 7.5e-21
+ eta0 = -0.00026219533
+ pvag = 0.0
+ etab = 0.0013487812
+ pvsat = 1.2452966e-11
+ la0 = 1.1871046e-7
+ vsat = 85400.58
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ wint = 3e-9
+ pute = -6.731688e-15
+ wketa = 4.614407e-9
+ lpdiblc2 = 5.562512e-9
+ pvth0 = -1.0421574e-15
+ jsw = 1.45e-12
+ vth0 = 0.486292
+ lk1 = 3.247429e-8
+ kt1 = -0.1929406
+ lk2 = -1.4947512e-8
+ kt2 = -0.03937921
+ drout = 0.0
+ rdsw = 170.0
+ llc = -0.039
+ lln = -1
+ tpbsw = 0.001554306
+ pscbe1 = 400000000.0
+ pscbe2 = 1e-6
+ lu0 = 1.6015452e-9
+ version = 3.24
+ wkt1 = -2.0427562e-8
+ wkt2 = 2.2519782e-9
+ lint = 1e-8
+ lua = 2.6581833e-17
+ lub = -8.899446e-26
+ luc = -1.5904941e-17
+ nch = 3.9e+17
+ wmax = 5e-7
+ lwl = 0.0
+ lwn = 1.0
+ wmin = 2.2e-7
+ pa0 = -9.128582e-14
+ nlx = 0.0
+ cjswg = 3.340547e-10
+ lkt1 = -4.834396e-10
+ lkt2 = 1.8777602e-9
+ mjswg = 0.43879
+ pk1 = 4.587708e-15
+ pk2 = -2.4446703e-15
+ lmax = 5e-7
+ nqsmod = 0
+ tpbswg = 0.001554306
+ lmin = 1.8e-7
+ noimod = 2
+ pu0 = -1.7230291e-17
+ prt = 0
+ pua = -2.3933522e-23
+ pub = 2.5580594e-32
+ puc = 3.433529e-24
+ wvoff = -3.98773e-10
+ rsh = 6.8
+ tcj = 0.001040287
+ ua1 = 1.224e-9
+ ub1 = -3.1027764e-18
+ uc1 = -2.4653823e-10
+ weta0 = 0
+ tpb = 0.001554306
+ wub1 = 1.602399e-25
+ wuc1 = 5.485366e-17
+ tox = 4.08e-9
+ wvsat = 0.0005899806
+ wa0 = 2.8954867e-7
+ hdif = 2e-7
+ lpclm = 7.125815e-8
+ wvth0 = -1.4909164e-8
+ ute = -1.9466008
+ wk1 = -1.9985334e-8
+ wk2 = 4.552045e-9
+ lub1 = 3.260553e-25
+ luc1 = 5.707747e-17
+ wute = 1.4634106e-8
+ wln = 1.0
+ mjsw = 0.2003879
+ wu0 = 1.2921135e-9
+ wua = 4.711108e-17
+ wub = -1.1345223e-25
+ wuc = -3.179524e-17
+ wwl = 0.0
+ wwn = 1
+ xti = 3
+ lute = 4.90364e-8
+ cdsc = 0.0
+ capmod = 3
+ cgdo = 3.665e-10
+ lketa = 4.87385e-10
+ cgso = 3.665e-10
+ xpart = 1
+ mobmod = 1
+ cjsw = 2.040547e-10
+ pbswg = 0.6882682
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ lvoff = -3.895271e-9
+ beta0 = 11.59263
+ leta0 = 1.6662733999999999e-10
+ tnom = 25.0
+ letab = -6.664392e-10
+ lvsat = -0.00020626588
+ pags = 5.067323e-15
+ lvth0 = 1.4483583e-8
+ toxm = 4.08e-9
+ nfactor = 1.0
+ pcit = 1.266836e-18
+ ppclm = -1.7902992e-16
+ pbsw = 0.6882682
+ pclm = 1.1355271
+ delta = 0.01
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ tcjswg = 0.000645489
+ pdiblc1 = 1e-6
+ pdiblc2 = -0.007140237
+ pdiblcb = 0.01
+ a0 = 0.270794
+ a1 = 0.0
+ a2 = 0.99
+ b0 = 0.0
+ b1 = 0.0
+ pnfactor = 0.0
+ )

.model nch_fs_1 nmos (
+ level = 49
+ cjsw = 1.93852e-10
+ drout = 0.0
+ tpbsw = 0.001554306
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ cjswg = 3.17352e-10
+ pnfactor = 0.0
+ mjswg = 0.43879
+ wnfactor = 0.0
+ tnom = 25.0
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ wvoff = 6.32688e-10
+ pscbe1 = 200000030.0
+ pscbe2 = 1e-6
+ toxm = 4.08e-9
+ version = 3.24
+ pbsw = 0.6882682
+ pclm = 0.8000001
+ weta0 = 0
+ wvsat = 0.0
+ nqsmod = 0
+ lnfactor = -4.5192e-8
+ tpbswg = 0.001554306
+ wvth0 = -5.9653440000000004e-9
+ noimod = 2
+ ags = 0.02
+ keta = 0.009263485
+ cit = -0.00010000001
+ a0 = 0.3700794
+ a1 = 0.0
+ a2 = 0.99
+ b0 = 0.0
+ b1 = 0.0
+ dlc = 3e-9
+ dsub = 0.0
+ k3b = 0.0
+ at = 20000.0
+ cf = 0
+ cj = 0.0009502527
+ ef = 0.874
+ k1 = 0.5142301
+ k2 = 0.007567123999999999
+ k3 = 0.0
+ em = 30000000.0
+ dwb = 0.0
+ dwg = 0.0
+ js = 3.5e-7
+ ll = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ u0 = 0.04401107
+ pb = 0.6882682
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ dvt0 = 0.0
+ ua = -6.12274e-10
+ dvt1 = 0.0
+ ub = 2.3135539e-18
+ xpart = 1
+ dvt2 = 0.0
+ uc = 1.0876087e-10
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ voff = -0.13786648
+ capmod = 3
+ ldif = 9e-8
+ pbswg = 0.6882682
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ jsw = 1.45e-12
+ kt1 = -0.2240464
+ lk2 = -3.6153600000000002e-9
+ kt2 = -0.030266136
+ lvoff = 9.038400000000001e-10
+ eta0 = 5e-5
+ llc = -0.039
+ lln = -1
+ pvag = 0.0
+ etab = -5e-5
+ lu0 = 4.5192000000000003e-10
+ vsat = 93615.37
+ beta0 = 11.59263
+ nch = 3.9e+17
+ wint = 3e-9
+ lwl = 0.0
+ lwn = 1.0
+ vth0 = 0.41802738
+ leta0 = 3.163440009680917e-10
+ mobmod = 1
+ nlx = 0.0
+ rdsw = 170.0
+ lint = 1e-8
+ wmax = 0.000900001
+ lvth0 = -2.621136e-9
+ pu0 = 0.0
+ wmin = 1e-5
+ prt = 0
+ lmax = 2.0001e-5
+ delta = 0.01
+ lmin = 1e-5
+ rsh = 6.8
+ tcj = 0.001040287
+ ua1 = 1.224e-9
+ ub1 = -1.1209314e-18
+ uc1 = 1.1643822e-11
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ tpb = 0.001554306
+ tox = 4.08e-9
+ ute = -1.5799998
+ wln = 1.0
+ wu0 = 0.0
+ nfactor = 1.0
+ hdif = 2e-7
+ wwl = 0.0
+ wwn = 1
+ xti = 3
+ mjsw = 0.2003879
+ tcjswg = 0.000645489
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0006999999
+ pdiblcb = 0.01
+ tcjsw = 0.000645489
+ cdsc = 0.0
+ pvoff = 9.038400000000001e-16
+ cgdo = 3.665e-10
+ binunit = 2
+ cgso = 3.665e-10
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 1.3557600041489644e-16
+ pvth0 = -2.71152e-15
+ )

.model nch_fs_2 nmos (
+ level = 49
+ wmax = 0.000900001
+ wmin = 1e-5
+ lkt2 = -4.553491e-12
+ lmax = 1e-5
+ lmin = 1.2e-6
+ la0 = -3.496093e-7
+ jsw = 1.45e-12
+ kt1 = -0.2240468
+ lk1 = 1.4908844e-8
+ kt2 = -0.03026568
+ lk2 = -1.472874e-8
+ llc = -0.039
+ lln = -1
+ lketa = -4.320781e-8
+ lu0 = 3.743729e-9
+ lua = -4.643216e-16
+ lub = 7.375677e-25
+ luc = 3.898355e-17
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ xpart = 1
+ pnfactor = 0.0
+ nlx = 0.0
+ hdif = 2e-7
+ wnfactor = 0.0
+ capmod = 3
+ lub1 = 4.527317e-28
+ luc1 = 7.827772e-20
+ nfactor = 1.0
+ pu0 = 0.0
+ mjsw = 0.2003879
+ prt = 0
+ pbswg = 0.6882682
+ lute = -5.743953e-11
+ lvoff = -9.567488e-9
+ rsh = 6.8
+ tcj = 0.001040287
+ ua1 = 1.224e-9
+ ub1 = -1.1209769e-18
+ uc1 = 1.1635963e-11
+ mobmod = 1
+ beta0 = 11.59263
+ tpb = 0.001554306
+ tox = 4.08e-9
+ lnfactor = -4.5192e-8
+ leta0 = 3.163440009680917e-10
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0003968181
+ cdsc = 0.0
+ pdiblcb = 0.01
+ lpscbe1 = 262.58185
+ ute = -1.5799941
+ lvsat = -0.006562638
+ cgdo = 3.665e-10
+ wln = 1.0
+ lvth0 = 5.799173400000001e-8
+ wu0 = 0.0
+ wwl = 0.0
+ wwn = 1
+ cgso = 3.665e-10
+ xti = 3
+ delta = 0.01
+ lpdiblc2 = 3.0196912e-9
+ binunit = 2
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ cjsw = 1.93852e-10
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ tnom = 25.0
+ tcjswg = 0.000645489
+ a0 = 0.4051808
+ a1 = 0.0
+ a2 = 0.99
+ b0 = 0.0
+ b1 = 0.0
+ at = 20000.0
+ cf = 0
+ cj = 0.0009502527
+ ef = 0.874
+ k1 = 0.5127332
+ k2 = 0.008682927
+ k3 = 0.0
+ em = 30000000.0
+ toxm = 4.08e-9
+ js = 3.5e-7
+ ll = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ u0 = 0.04368057
+ pb = 0.6882682
+ w0 = 0.0
+ pbsw = 0.6882682
+ rd = 0
+ pclm = 0.7736172
+ rs = 0
+ ua = -5.656554e-10
+ ub = 2.2395009e-18
+ uc = 1.0484686e-10
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ tcjsw = 0.000645489
+ version = 3.24
+ pvoff = 9.038400000000001e-16
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 1.3557600041489644e-16
+ pvth0 = -2.71152e-15
+ keta = 0.013601619
+ drout = 0.0
+ tpbsw = 0.001554306
+ dsub = 0.0
+ cjswg = 3.17352e-10
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ mjswg = 0.43879
+ pscbe1 = 173636400.0
+ pscbe2 = 1e-6
+ lcit = 2.6652053e-10
+ wvoff = 6.32688e-10
+ voff = -0.13681518
+ ldif = 9e-8
+ ags = 0.02
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ weta0 = 0
+ nqsmod = 0
+ eta0 = 5e-5
+ tpbswg = 0.001554306
+ pvag = 0.0
+ etab = -5e-5
+ cit = -0.00012675911
+ noimod = 2
+ wvsat = 0.0
+ vsat = 94274.27
+ wint = 3e-9
+ dlc = 3e-9
+ lpclm = 2.6277317e-7
+ wvth0 = -5.9653440000000004e-9
+ vth0 = 0.41194178
+ k3b = 0.0
+ rdsw = 170.0
+ dwb = 0.0
+ dwg = 0.0
+ lint = 1e-8
+ )

.model nch_fs_3 nmos (
+ level = 49
+ beta0 = 11.59263
+ leta0 = 3.544582809680917e-10
+ letab = -3.811428e-11
+ lvsat = -0.0007622857
+ version = 3.24
+ lvth0 = 1.3216209999999997e-9
+ delta = 0.01
+ keta = -0.015927497
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ dsub = 0.0
+ pnfactor = 0.0
+ lags = -3.044698e-8
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ tcjswg = 0.000645489
+ wnfactor = 0.0
+ lcit = 3.0262734e-10
+ voff = -0.15940708
+ ldif = 9e-8
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ eta0 = 1.7142866e-5
+ pvag = 0.0
+ etab = -1.7142866e-5
+ vsat = 89273.96
+ tcjsw = 0.000645489
+ lnfactor = -4.5192e-8
+ wint = 3e-9
+ vth0 = 0.46079528
+ rdsw = 170.0
+ pvoff = 9.038400000000001e-16
+ lint = 1e-8
+ wmax = 0.000900001
+ wmin = 1e-5
+ cdscb = 0.0
+ cdscd = 0.0
+ lkt1 = 5.782678e-9
+ lkt2 = 1.5570838e-9
+ peta0 = 1.3557600041489644e-16
+ lmax = 1.2e-6
+ lpdiblc2 = 1.525682e-9
+ lmin = 5e-7
+ pvth0 = -2.71152e-15
+ ags = 0.0462474
+ drout = 0.0
+ tpbsw = 0.001554306
+ cit = -0.00015788565
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ dlc = 3e-9
+ cjswg = 3.17352e-10
+ k3b = 0.0
+ pscbe1 = 400000100.0
+ pscbe2 = 1e-6
+ mjswg = 0.43879
+ dwb = 0.0
+ dwg = 0.0
+ hdif = 2e-7
+ lua1 = -3.0446746e-18
+ lub1 = -1.2004175e-24
+ luc1 = -6.517273e-17
+ wvoff = 6.32688e-10
+ mjsw = 0.2003879
+ nqsmod = 0
+ tpbswg = 0.001554306
+ noimod = 2
+ nfactor = 1.0
+ lute = -2.6630502e-7
+ weta0 = 0
+ la0 = 4.581426e-7
+ wvsat = 0.0
+ jsw = 1.45e-12
+ kt1 = -0.2290285
+ lk1 = -7.214246e-9
+ kt2 = -0.031611919
+ lk2 = -1.9122090000000005e-9
+ lpclm = 1.5245718e-7
+ wvth0 = -5.9653440000000004e-9
+ a0 = -0.2911571
+ a1 = 0.0
+ a2 = 0.99
+ b0 = 0.0
+ b1 = 0.0
+ llc = -0.039
+ cdsc = 0.0
+ lln = -1
+ lu0 = 1.4925279e-9
+ at = 20000.0
+ cf = 0
+ cj = 0.0009502527
+ ef = 0.874
+ k1 = 0.5318048
+ k2 = -0.002365807
+ k3 = 0.0
+ em = 30000000.0
+ lua = 7.982966e-17
+ lub = -1.5630905e-25
+ luc = -9.669895e-18
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ js = 3.5e-7
+ cgdo = 3.665e-10
+ ll = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0016847569
+ u0 = 0.04562126
+ pb = 0.6882682
+ w0 = 0.0
+ rd = 0
+ nlx = 0.0
+ rs = 0
+ pdiblcb = 0.01
+ ua = -1.0347512e-9
+ ub = 3.0100842e-18
+ uc = 1.4678947e-10
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ cgso = 3.665e-10
+ pu0 = 0.0
+ prt = 0
+ cjsw = 1.93852e-10
+ binunit = 2
+ rsh = 6.8
+ tcj = 0.001040287
+ ua1 = 1.2266247e-9
+ ub1 = -8.574386e-20
+ uc1 = 6.788683e-11
+ lketa = -8.954029e-9
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ tpb = 0.001554306
+ tox = 4.08e-9
+ capmod = 3
+ xpart = 1
+ ute = -1.3504703
+ tnom = 25.0
+ wln = 1.0
+ wu0 = 0.0
+ pbswg = 0.6882682
+ wwl = 0.0
+ wwn = 1
+ xti = 3
+ toxm = 4.08e-9
+ mobmod = 1
+ lvoff = 1.6639098000000002e-8
+ pbsw = 0.6882682
+ pclm = 0.8687172
+ )

.model nch_fs_4 nmos (
+ level = 49
+ lua1 = 8.039099e-19
+ lub1 = 3.824101e-25
+ luc1 = 2.9606131e-17
+ mjsw = 0.2003879
+ lute = 7.030476e-8
+ ags = -0.019916179
+ tcjsw = 0.000645489
+ nfactor = 1.0
+ cdsc = 0.0
+ cit = 0.000271889
+ pvoff = 9.038400000000001e-16
+ dlc = 3e-9
+ cgdo = 3.665e-10
+ k3b = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cgso = 3.665e-10
+ peta0 = 1.3557600041489644e-16
+ pdiblc1 = 1e-6
+ pdiblc2 = -0.00593541
+ pdiblcb = 0.01
+ pvth0 = -2.71152e-15
+ drout = 0.0
+ alpha0 = 0.0
+ cjsw = 1.93852e-10
+ alpha1 = 0.448150714
+ tpbsw = 0.001554306
+ la0 = 7.545271e-8
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ pscbe1 = 400000000.0
+ pscbe2 = 1e-6
+ binunit = 2
+ jsw = 1.45e-12
+ kt1 = -0.22715
+ lk1 = 4.899558e-8
+ kt2 = -0.029537767
+ lk2 = -2.6956696000000003e-8
+ cjswg = 3.17352e-10
+ pnfactor = 0.0
+ llc = -0.039
+ lln = -1
+ mjswg = 0.43879
+ lu0 = 1.7037189e-9
+ wnfactor = 0.0
+ lua = -1.0530929e-18
+ lub = 5.559478e-27
+ luc = 4.133919e-18
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ tnom = 25.0
+ nqsmod = 0
+ tpbswg = 0.001554306
+ wvoff = 6.32688e-10
+ nlx = 0.0
+ noimod = 2
+ toxm = 4.08e-9
+ pu0 = 0.0
+ weta0 = 0
+ pbsw = 0.6882682
+ pclm = 1.1076791
+ prt = 0
+ wvsat = 0.0
+ lnfactor = -4.5192e-8
+ lpclm = 4.253467e-8
+ wvth0 = -5.9653440000000004e-9
+ rsh = 6.8
+ tcj = 0.001040287
+ ua1 = 1.2182583e-9
+ ub1 = -3.526674e-18
+ uc1 = -1.381542e-10
+ tpb = 0.001554306
+ tox = 4.08e-9
+ ute = -2.0822308
+ version = 3.24
+ wln = 1.0
+ wu0 = 0.0
+ lpdiblc2 = 5.030957e-9
+ wwl = 0.0
+ wwn = 1
+ xti = 3
+ keta = -0.04182327
+ capmod = 3
+ dsub = 0.0
+ lketa = 2.9580252e-9
+ xpart = 1
+ lags = -1.1735286e-11
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ lcit = 1.0493098e-10
+ voff = -0.12183828000000001
+ pbswg = 0.6882682
+ mobmod = 1
+ ldif = 9e-8
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ lvoff = -6.425217999999999e-10
+ eta0 = -0.0002937502
+ pvag = 0.0
+ etab = 0.0013875004
+ beta0 = 11.59263
+ vsat = 88054.32
+ wint = 3e-9
+ leta0 = 4.974690609680917e-10
+ vth0 = 0.45670238
+ letab = -6.842502e-10
+ rdsw = 170.0
+ lvsat = -0.00020125005
+ lint = 1e-8
+ lvth0 = 3.2043650000000002e-9
+ wmax = 0.000900001
+ wmin = 1e-5
+ lkt1 = 4.918561e-9
+ lkt2 = 6.029743e-10
+ delta = 0.01
+ lmax = 5e-7
+ a0 = 0.5407774
+ a1 = 0.0
+ a2 = 0.99
+ b0 = 0.0
+ b1 = 0.0
+ lmin = 1.8e-7
+ at = 20000.0
+ cf = 0
+ cj = 0.0009502527
+ ef = 0.874
+ k1 = 0.4096095
+ k2 = 0.05207874
+ k3 = 0.0
+ em = 30000000.0
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ js = 3.5e-7
+ ll = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ u0 = 0.04516215
+ pb = 0.6882682
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ua = -8.589192e-10
+ ub = 2.6581962e-18
+ uc = 1.1678118e-10
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ tcjswg = 0.000645489
+ hdif = 2e-7
+ )

.model nch_fs_5 nmos (
+ level = 49
+ pu0 = 0.0
+ pscbe1 = 200000030.0
+ pscbe2 = 1e-6
+ tpbsw = 0.001554306
+ prt = 0
+ dsub = 0.0
+ cjswg = 3.17352e-10
+ rsh = 6.8
+ tcj = 0.001040287
+ ua1 = 1.224e-9
+ ub1 = -1.0684574e-18
+ a0 = 0.3702259
+ a1 = 0.0
+ a2 = 0.99
+ uc1 = 2.4230474e-11
+ b0 = 0.0
+ b1 = 0.0
+ mjswg = 0.43879
+ nqsmod = 0
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ tpbswg = 0.001554306
+ at = 20000.0
+ cf = 0
+ cj = 0.0009502527
+ ef = 0.874
+ k1 = 0.5102321
+ k2 = 0.008860774000000002
+ k3 = 0.0
+ tpb = 0.001554306
+ noimod = 2
+ em = 30000000.0
+ tox = 4.08e-9
+ js = 3.5e-7
+ wa0 = -1.4643313e-9
+ ll = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ wvoff = 1.5234104e-9
+ u0 = 0.04484358
+ pb = 0.6882682
+ w0 = 0.0
+ rd = 0
+ ute = -1.5803809
+ rs = 0
+ ua = -5.885942e-10
+ ub = 2.3329335e-18
+ uc = 1.1057788e-10
+ voff = -0.13795558
+ wk1 = 3.995606e-8
+ wk2 = -1.2928737e-8
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -2e-8
+ ww = 0.0
+ ldif = 9e-8
+ xw = 0.0
+ wln = 1.0
+ wu0 = -8.320099e-9
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ puc1 = -1.4905616e-28
+ weta0 = 0
+ wua = -2.3665659e-16
+ wub = -1.936796e-25
+ wuc = -1.815927e-17
+ wwl = 0.0
+ wwn = 1
+ eta0 = 5e-5
+ xti = 3
+ wvsat = 0.0
+ pvag = 0.0
+ etab = -5e-5
+ vsat = 93615.37
+ wvth0 = -5.2777326e-9
+ wint = 3e-9
+ vth0 = 0.41795858
+ rdsw = 170.0
+ wkt1 = -8.215166e-9
+ wkt2 = 1.6245854e-9
+ lint = 1e-8
+ wmax = 1e-5
+ wmin = 1.2e-6
+ lmax = 2.0001e-5
+ lmin = 1e-5
+ capmod = 3
+ xpart = 1
+ wub1 = -5.244247e-25
+ pnfactor = 0.0
+ wuc1 = -1.257911e-16
+ wnfactor = 0.0
+ hdif = 2e-7
+ mobmod = 1
+ wute = 3.808433e-9
+ pbswg = 0.6882682
+ mjsw = 0.2003879
+ lvoff = 9.038400000000001e-10
+ beta0 = 11.59263
+ lnfactor = -4.5192e-8
+ leta0 = 3.163440009680917e-10
+ cdsc = 0.0
+ nfactor = 1.0
+ lvth0 = -2.621136e-9
+ cgdo = 3.665e-10
+ cgso = 3.665e-10
+ delta = 0.01
+ dvt0w = 0.0
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0006999999
+ dvt1w = 0.0
+ dvt2w = 0.0
+ pdiblcb = 0.01
+ cjsw = 1.93852e-10
+ tcjswg = 0.000645489
+ ags = 0.02
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ cit = -0.00010000001
+ binunit = 2
+ dlc = 3e-9
+ tnom = 25.0
+ k3b = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ toxm = 4.08e-9
+ pbsw = 0.6882682
+ pclm = 0.8000001
+ tcjsw = 0.000645489
+ pvoff = 9.038400000000001e-16
+ jsw = 1.45e-12
+ kt1 = -0.2232244
+ kt2 = -0.030428693
+ lk2 = -3.6153600000000002e-9
+ llc = -0.039
+ lln = -1
+ lu0 = 4.5192000000000003e-10
+ cdscb = 0.0
+ cdscd = 0.0
+ nch = 3.9e+17
+ peta0 = 1.3557600041489644e-16
+ lwl = 0.0
+ lwn = 1.0
+ nlx = 0.0
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ version = 3.24
+ wketa = -1.0935369e-8
+ pvth0 = -2.71152e-15
+ keta = 0.010357677
+ drout = 0.0
+ )

.model nch_fs_6 nmos (
+ level = 49
+ nfactor = 1.0
+ cgso = 3.665e-10
+ capmod = 3
+ cjsw = 1.93852e-10
+ lketa = -4.518989e-8
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0003968181
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ pdiblcb = 0.01
+ lpscbe1 = 262.58185
+ xpart = 1
+ mobmod = 1
+ tnom = 25.0
+ pbswg = 0.6882682
+ binunit = 2
+ toxm = 4.08e-9
+ lvoff = -9.902212e-9
+ a0 = 0.40626
+ a1 = 0.0
+ a2 = 0.99
+ b0 = 0.0
+ b1 = 0.0
+ pbsw = 0.6882682
+ pclm = 0.7755287
+ at = 20000.0
+ cf = 0
+ cj = 0.0009502527
+ ef = 0.874
+ k1 = 0.508509
+ beta0 = 11.59263
+ k2 = 0.01007951
+ k3 = 0.0
+ em = 30000000.0
+ js = 3.5e-7
+ ll = 0.0
+ leta0 = 3.163440009680917e-10
+ mj = 0.3595262
+ lw = 0.0
+ u0 = 0.04453795
+ pb = 0.6882682
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ags = 0.02
+ ua = -5.377125e-10
+ ub = 2.2537915e-18
+ uc = 1.0657759e-10
+ lvsat = -0.006753025
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ lvth0 = 5.8084954e-8
+ cit = -0.00012675911
+ ppclm = 1.9027247e-13
+ delta = 0.01
+ dlc = 3e-9
+ k3b = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ tcjswg = 0.000645489
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ pkt1 = 4.710912e-15
+ pkt2 = -4.130377e-15
+ keta = 0.014894814
+ version = 3.24
+ dsub = 0.0
+ pnfactor = 0.0
+ la0 = -3.588995e-7
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ wnfactor = 0.0
+ jsw = 1.45e-12
+ lk1 = 1.7161611e-8
+ kt1 = -0.2231775
+ lk2 = -1.5753972e-8
+ kt2 = -0.030469729
+ pketa = 1.9809019e-14
+ llc = -0.039
+ lln = -1
+ lu0 = 3.4960111999999998e-9
+ lcit = 2.6652053e-10
+ voff = -0.13687068
+ lua = -5.067804e-16
+ lub = 7.882536e-25
+ luc = 3.984287e-17
+ nch = 3.9e+17
+ ldif = 9e-8
+ lwl = 0.0
+ lwn = 1.0
+ wpclm = -1.9103656e-8
+ kt1l = 0.0
+ pa0 = 9.284546e-14
+ prwb = 0.0
+ prwg = 0.0
+ pub1 = 4.176128e-31
+ nlx = 0.0
+ puc1 = 7.417578e-23
+ eta0 = 5e-5
+ pk1 = -2.2514154e-14
+ pk2 = 1.0246181e-14
+ pvag = 0.0
+ etab = -5e-5
+ tcjsw = 0.000645489
+ pu0 = 2.4756895e-15
+ vsat = 94293.38
+ lnfactor = -4.5192e-8
+ wint = 3e-9
+ pute = -5.708167e-14
+ prt = 0
+ pua = 4.243342e-22
+ pub = -5.065558e-31
+ puc = -8.588134e-24
+ vth0 = 0.41186368
+ rdsw = 170.0
+ pvoff = 4.249081000000001e-15
+ wkt1 = -8.688151e-9
+ wkt2 = 2.0392819e-9
+ rsh = 6.8
+ lint = 1e-8
+ tcj = 0.001040287
+ ua1 = 1.224e-9
+ ub1 = -1.0643074e-18
+ uc1 = 2.4967807e-11
+ wmax = 1e-5
+ wmin = 1.2e-6
+ cdscb = 0.0
+ cdscd = 0.0
+ tpb = 0.001554306
+ peta0 = 1.3557600041489644e-16
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ tox = 4.08e-9
+ lkt1 = -4.674615e-10
+ lkt2 = 4.087321e-10
+ wa0 = -1.0786144e-8
+ lpdiblc2 = 3.0196912e-9
+ lmax = 1e-5
+ pvsat = 1.9027204e-9
+ ute = -1.5809486
+ pscbe1 = 173636400.0
+ pscbe2 = 1e-6
+ wk1 = 4.221652e-8
+ wk2 = -1.3957471e-8
+ lmin = 1.2e-6
+ wketa = -1.292423e-8
+ pvth0 = -3.6432075e-15
+ wln = 1.0
+ drout = 0.0
+ wu0 = -8.568663e-9
+ tpbsw = 0.001554306
+ wua = -2.7926046e-16
+ wub = -1.4282058e-25
+ wuc = -1.7297008e-17
+ wwl = 0.0
+ wwn = 1
+ xti = 3
+ nqsmod = 0
+ tpbswg = 0.001554306
+ cjswg = 3.17352e-10
+ noimod = 2
+ wub1 = -5.663537e-25
+ wuc1 = -1.3323848e-16
+ mjswg = 0.43879
+ hdif = 2e-7
+ wvoff = 1.1875419e-9
+ lub1 = -4.133362e-26
+ luc1 = -7.343755e-18
+ wute = 9.539526e-9
+ mjsw = 0.2003879
+ weta0 = 0
+ lute = 5.654154e-9
+ wvsat = -0.00019104627
+ lpclm = 2.4373449e-7
+ wvth0 = -5.184193800000001e-9
+ cdsc = 0.0
+ cgdo = 3.665e-10
+ )

.model nch_fs_7 nmos (
+ level = 49
+ beta0 = 11.59263
+ pvag = 0.0
+ etab = -1.7142869e-5
+ vsat = 89128.95
+ leta0 = 3.544582809680917e-10
+ wint = 3e-9
+ pute = 4.357466e-13
+ letab = -3.811428e-11
+ vth0 = 0.46146618
+ lvsat = -0.0007622865
+ rdsw = 170.0
+ lvth0 = 5.459959999999999e-10
+ wkt1 = -3.681822e-9
+ wkt2 = -1.3190541e-9
+ lint = 1e-8
+ wmax = 1e-5
+ la0 = 4.645035e-7
+ ppclm = 7.258032e-15
+ wmin = 1.2e-6
+ jsw = 1.45e-12
+ lk1 = -1.1179709e-8
+ kt1 = -0.2286601
+ lk2 = -1.8429500000000034e-10
+ kt2 = -0.031479932
+ delta = 0.01
+ tcjswg = 0.000645489
+ lkt1 = 5.892387e-9
+ lkt2 = 1.5805686e-9
+ llc = -0.039
+ lln = -1
+ lmax = 1.2e-6
+ lu0 = 1.4123913000000001e-9
+ lmin = 5e-7
+ lua = 6.148926e-17
+ lub = -1.2783527e-25
+ luc = -6.505068e-18
+ nch = 3.9e+17
+ dvt0w = 0.0
+ lwl = 0.0
+ lwn = 1.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ pa0 = -6.357063e-14
+ nlx = 0.0
+ pk1 = 3.963084e-14
+ pk2 = -1.7268767e-14
+ pu0 = 8.008865e-16
+ prt = 0
+ pua = 1.8329395e-22
+ pub = -2.8456703e-31
+ puc = -3.16293e-23
+ wua1 = -3.55913e-18
+ wub1 = -1.6132161e-24
+ wuc1 = -1.8047248e-16
+ hdif = 2e-7
+ rsh = 6.8
+ pketa = 9.843987e-15
+ tcj = 0.001040287
+ ua1 = 1.2269809e-9
+ ub1 = 7.567455e-20
+ lua1 = -3.457781e-18
+ uc1 = 8.594492e-11
+ lub1 = -1.3637128e-24
+ luc1 = -7.807721e-17
+ wute = -4.153124e-7
+ mjsw = 0.2003879
+ tpb = 0.001554306
+ tox = 4.08e-9
+ wa0 = 1.2405528e-7
+ wpclm = 1.3866737e-7
+ ute = -1.3089141
+ lute = -3.0990586e-7
+ wk1 = -1.1356744e-8
+ wk2 = 9.762311e-9
+ wln = 1.0
+ tcjsw = 0.000645489
+ wu0 = -7.124867e-9
+ wua = -7.146715e-17
+ wub = -3.341902e-25
+ wuc = 2.5660584e-18
+ wwl = 0.0
+ wwn = 1
+ xti = 3
+ cdsc = 0.0
+ pvoff = -2.109974e-15
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ cgdo = 3.665e-10
+ a0 = -0.3035701
+ a1 = 0.0
+ a2 = 0.99
+ b0 = 0.0
+ b1 = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 1.3557600041489644e-16
+ at = 20000.0
+ cf = 0
+ cj = 0.0009502527
+ pscbe1 = 400000100.0
+ pscbe2 = 1e-6
+ ef = 0.874
+ k1 = 0.5329412
+ k2 = -0.0033426250000000005
+ k3 = 0.0
+ em = 30000000.0
+ cgso = 3.665e-10
+ js = 3.5e-7
+ ll = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ u0 = 0.04633417
+ pb = 0.6882682
+ nfactor = 1.0
+ w0 = 0.0
+ rd = 0
+ wketa = -4.333682e-9
+ rs = 0
+ ua = -1.0276002e-9
+ ub = 3.0435232e-18
+ uc = 1.4653272e-10
+ pvth0 = 5.040078e-15
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ drout = 0.0
+ tpbsw = 0.001554306
+ nqsmod = 0
+ cjsw = 1.93852e-10
+ tpbswg = 0.001554306
+ noimod = 2
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ cjswg = 3.17352e-10
+ pnfactor = 0.0
+ mjswg = 0.43879
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0017737894
+ pdiblcb = 0.01
+ wnfactor = 0.0
+ tnom = 25.0
+ wvoff = 6.6694859999999994e-9
+ pags = 4.128623e-14
+ toxm = 4.08e-9
+ weta0 = 0
+ ppdiblc2 = 1.0321563e-15
+ binunit = 2
+ pbsw = 0.6882682
+ pclm = 0.8548421
+ wvsat = 0.0014492224
+ wpdiblc2 = -8.897895e-10
+ lpclm = 1.5173094e-7
+ wvth0 = -1.266978e-8
+ lnfactor = -4.5192e-8
+ capmod = 3
+ lpdiblc2 = 1.4224044e-9
+ pkt1 = -1.0964308e-15
+ pkt2 = -2.3470743e-16
+ keta = -0.01549387
+ lketa = -9.939018e-9
+ mobmod = 1
+ wags = -3.559157e-8
+ dsub = 0.0
+ version = 3.24
+ xpart = 1
+ ags = 0.04980868
+ lags = -3.457808e-8
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ cit = -0.00015788565
+ pbswg = 0.6882682
+ lcit = 3.0262734e-10
+ voff = -0.16001108
+ ldif = 9e-8
+ dlc = 3e-9
+ k3b = 0.0
+ kt1l = 0.0
+ lvoff = 1.6940662e-8
+ pua1 = 4.128591e-24
+ prwb = 0.0
+ prwg = 0.0
+ pub1 = 1.6319734e-30
+ puc1 = 1.2896722e-22
+ dwb = 0.0
+ dwg = 0.0
+ eta0 = 1.7142869e-5
+ )

.model nch_fs_8 nmos (
+ level = 49
+ pketa = -2.7027957e-15
+ tnom = 25.0
+ pdiblc1 = 1e-6
+ pdiblc2 = -0.006119013
+ pdiblcb = 0.01
+ pags = -1.0838496e-14
+ toxm = 4.08e-9
+ wpclm = 6.656068e-8
+ pcit = 1.4220811e-17
+ pbsw = 0.6882682
+ pclm = 1.1010191
+ tcjsw = 0.000645489
+ binunit = 2
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ pvoff = -7.157499999999998e-17
+ pscbe1 = 400000000.0
+ pscbe2 = 1e-6
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 1.3419387861489644e-16
+ petab = 1.6959704e-18
+ pvsat = 1.5350395e-12
+ wketa = 2.2941933e-8
+ nqsmod = 0
+ pvth0 = 1.797418e-15
+ tpbswg = 0.001554306
+ drout = 0.0
+ noimod = 2
+ pkt1 = -1.7512235e-15
+ pkt2 = 7.382567e-17
+ keta = -0.04411884
+ tpbsw = 0.001554306
+ wags = 7.772305e-8
+ dsub = 0.0
+ cjswg = 3.17352e-10
+ mjswg = 0.43879
+ lags = 1.0727657e-9
+ wcit = -3.0914837e-11
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ version = 3.24
+ wvoff = 2.2381844e-9
+ lcit = 1.0350804e-10
+ voff = -0.12199898
+ ldif = 9e-8
+ weta0 = 3.0046217e-12
+ kt1l = 0.0
+ pua1 = -1.0901051e-24
+ prwb = 0.0
+ prwg = 0.0
+ pub1 = -4.238914e-31
+ puc1 = -2.7204607e-23
+ wetab = -3.686654e-12
+ wvsat = 0.0014459029
+ eta0 = -0.00029405078
+ pvag = 0.0
+ etab = 0.0013878694
+ lpclm = 3.848953e-8
+ wvth0 = -5.6205204000000005e-9
+ vsat = 87909.64
+ wint = 3e-9
+ pute = -1.178615e-13
+ vth0 = 0.45666788
+ rdsw = 170.0
+ capmod = 3
+ wkt1 = -2.2583577e-9
+ wkt2 = -1.9897783e-9
+ lint = 1e-8
+ ags = -0.027693154
+ wmax = 1e-5
+ wmin = 1.2e-6
+ lkt1 = 5.093789e-9
+ lkt2 = 5.955873e-10
+ lmax = 5e-7
+ cit = 0.00027498236
+ lmin = 1.8e-7
+ dlc = 3e-9
+ mobmod = 1
+ k3b = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ a0 = 0.5262308
+ a1 = 0.0
+ a2 = 0.99
+ lketa = 3.228467e-9
+ b0 = 0.0
+ b1 = 0.0
+ at = 20000.0
+ cf = 0
+ cj = 0.0009502527
+ ef = 0.874
+ k1 = 0.4007356
+ k2 = 0.055957879999999995
+ k3 = 0.0
+ em = 30000000.0
+ xpart = 1
+ js = 3.5e-7
+ ll = 0.0
+ pnfactor = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ u0 = 0.04564852
+ wua1 = 7.785862e-18
+ pb = 0.6882682
+ wub1 = 2.8560549e-24
+ w0 = 0.0
+ wuc1 = 1.5903152e-16
+ rd = 0
+ rs = 0
+ ua = -9.017296e-10
+ ub = 2.7527719e-18
+ uc = 1.2291169e-10
+ wnfactor = 0.0
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ hdif = 2e-7
+ lua1 = 9.129858e-19
+ lub1 = 4.248247e-25
+ la0 = 8.279508e-8
+ luc1 = 3.232822e-17
+ pbswg = 0.6882682
+ wute = 7.881835e-7
+ mjsw = 0.2003879
+ jsw = 1.45e-12
+ lk1 = 4.963488e-8
+ kt1 = -0.226924
+ lk2 = -2.7462524e-8
+ kt2 = -0.029338669
+ llc = -0.039
+ lvoff = -5.449216999999999e-10
+ lln = -1
+ lu0 = 1.7277892e-9
+ ppdiblc2 = -2.2121929e-16
+ lute = 8.209799e-8
+ lua = 3.588764e-18
+ lub = 5.910339e-27
+ luc = 4.360599e-18
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ wpdiblc2 = 1.8349379e-9
+ beta0 = 11.59263
+ pa0 = -7.337964e-14
+ lnfactor = -4.5192e-8
+ nlx = 0.0
+ leta0 = 4.976073409680917e-10
+ letab = -6.844199e-10
+ pk1 = -6.389182e-15
+ pk2 = 5.055259e-15
+ lvsat = -0.00020140363
+ cdsc = 0.0
+ pu0 = -2.4055863e-16
+ lvth0 = 2.7532000000000004e-9
+ prt = 0
+ pua = -4.639069e-23
+ pub = -3.506499e-33
+ puc = -2.2654354e-24
+ cgdo = 3.665e-10
+ tcjswg = 0.000645489
+ ppclm = 4.042711e-14
+ delta = 0.01
+ cgso = 3.665e-10
+ rsh = 6.8
+ tcj = 0.001040287
+ lpdiblc2 = 5.053093e-9
+ ua1 = 1.2174792e-9
+ ub1 = -3.81245e-18
+ uc1 = -1.540669e-10
+ tpb = 0.001554306
+ tox = 4.08e-9
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ wa0 = 1.4537927e-7
+ nfactor = 1.0
+ ute = -2.1610963
+ cjsw = 1.93852e-10
+ wk1 = 8.868675e-8
+ wk2 = -3.876818e-8
+ wln = 1.0
+ wu0 = -4.860856e-9
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ wua = 4.278473e-16
+ wub = -9.451913e-25
+ wuc = -6.126842e-17
+ wwl = 0.0
+ wwn = 1
+ xti = 3
+ )

.model nch_fs_9 nmos (
+ level = 49
+ cjswg = 3.17352e-10
+ mjswg = 0.43879
+ wub1 = -7.675553e-27
+ wuc1 = -1.4706552e-17
+ hdif = 2e-7
+ wvoff = -2.3388100000000003e-10
+ ags = 0.02
+ wute = 3.836007e-8
+ mjsw = 0.2003879
+ weta0 = 0
+ cit = -0.00010000004
+ wvsat = 0.0
+ dlc = 3e-9
+ k3b = 0.0
+ wvth0 = -1.0228453e-8
+ dwb = 0.0
+ dwg = 0.0
+ capmod = 3
+ cdsc = 0.0
+ cgdo = 3.665e-10
+ cgso = 3.665e-10
+ mobmod = 1
+ jsw = 1.45e-12
+ kt1 = -0.2313184
+ lk2 = -3.6153600000000002e-9
+ kt2 = -0.029076951
+ llc = -0.039
+ lln = -1
+ lu0 = 4.5192000000000003e-10
+ cjsw = 1.93852e-10
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ nlx = 0.0
+ nfactor = 1.0
+ xpart = 1
+ pu0 = 0.0
+ prt = 0
+ tnom = 25.0
+ pbswg = 0.6882682
+ rsh = 6.8
+ tcj = 0.001040287
+ ua1 = 1.224e-9
+ pdiblc1 = 1e-6
+ toxm = 4.08e-9
+ pdiblc2 = 0.0007000003
+ ub1 = -1.5012456e-18
+ lvoff = 9.038400000000001e-10
+ uc1 = -6.880516e-11
+ pdiblcb = 0.01
+ pbsw = 0.6882682
+ tpb = 0.001554306
+ pclm = 0.8000001
+ tox = 4.08e-9
+ beta0 = 11.59263
+ wa0 = 7.667051e-8
+ leta0 = 3.163440009680917e-10
+ ute = -1.6093186
+ wk1 = -2.074723e-8
+ wk2 = 4.920634e-9
+ tcjswg = 0.000645489
+ wln = 1.0
+ wu0 = 1.0362965e-9
+ lvth0 = -2.621136e-9
+ binunit = 2
+ wua = 1.4309126e-16
+ wub = -1.5411778e-25
+ wuc = -1.4141237e-17
+ wwl = 0.0
+ wwn = 1
+ xti = 3
+ delta = 0.01
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ keta = 0.0010152902
+ dsub = 0.0
+ pnfactor = 0.0
+ wnfactor = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ a0 = 0.3047864
+ a1 = 0.0
+ a2 = 0.99
+ b0 = 0.0
+ b1 = 0.0
+ voff = -0.13648388
+ version = 3.24
+ at = 20000.0
+ cf = 0
+ cj = 0.0009502527
+ ldif = 9e-8
+ ef = 0.874
+ k1 = 0.5610723
+ k2 = -0.0060884483
+ k3 = 0.0
+ em = 30000000.0
+ kt1l = 0.0
+ js = 3.5e-7
+ prwb = 0.0
+ ll = 0.0
+ prwg = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ u0 = 0.037007399999999996
+ pb = 0.6882682
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ua = -9.066409e-10
+ ub = 2.2997995e-18
+ uc = 1.072127e-10
+ eta0 = 5e-5
+ wl = 0.0
+ tcjsw = 0.000645489
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -2e-8
+ ww = 0.0
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ xw = 0.0
+ pvag = 0.0
+ etab = -5e-5
+ lnfactor = -4.5192e-8
+ vsat = 93615.37
+ wint = 3e-9
+ pscbe1 = 200000030.0
+ pscbe2 = 1e-6
+ vth0 = 0.42210498
+ pvoff = 9.038400000000001e-16
+ rdsw = 170.0
+ wkt1 = 1.4490446e-9
+ wkt2 = 1.0605161e-11
+ lint = 1e-8
+ wmax = 1.2e-6
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 1.3557600041489644e-16
+ wmin = 5e-7
+ nqsmod = 0
+ tpbswg = 0.001554306
+ noimod = 2
+ lmax = 2.0001e-5
+ wketa = 2.1944087e-10
+ pvth0 = -2.71152e-15
+ lmin = 1e-5
+ drout = 0.0
+ tpbsw = 0.001554306
+ )

.model nch_fs_10 nmos (
+ level = 49
+ lute = -1.2190513e-8
+ nqsmod = 0
+ tpbswg = 0.001554306
+ noimod = 2
+ cdsc = 0.0
+ cgdo = 3.665e-10
+ nfactor = 1.0
+ lketa = -2.8027248e-8
+ cgso = 3.665e-10
+ xpart = 1
+ cjsw = 1.93852e-10
+ pbswg = 0.6882682
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0003968185
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ pdiblcb = 0.01
+ lpscbe1 = 262.58185
+ lvoff = -2.6983819999999998e-9
+ capmod = 3
+ beta0 = 11.59263
+ tnom = 25.0
+ leta0 = 3.163440009680917e-10
+ binunit = 2
+ lvsat = -0.006201102
+ toxm = 4.08e-9
+ lvth0 = 6.329934400000001e-8
+ pcit = 4.302753e-19
+ pbsw = 0.6882682
+ pclm = 0.7699873
+ ppclm = 1.243718e-13
+ mobmod = 1
+ delta = 0.01
+ ags = 0.02
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ cit = -0.00012672294
+ dlc = 3e-9
+ k3b = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ pnfactor = 0.0
+ pkt1 = 7.833639e-15
+ pkt2 = 9.747044e-16
+ keta = 0.00382927
+ wnfactor = 0.0
+ pketa = -6.831802e-16
+ version = 3.24
+ dsub = 0.0
+ wpclm = -1.2487239e-8
+ wcit = -4.317371e-14
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ la0 = -1.9725388e-7
+ tcjsw = 0.000645489
+ jsw = 1.45e-12
+ tcjswg = 0.000645489
+ lk1 = 1.0512358e-8
+ kt1 = -0.2310088
+ lk2 = -9.025411e-9
+ kt2 = -0.028688708
+ lcit = 2.6616018e-10
+ llc = -0.039
+ lln = -1
+ voff = -0.13612218
+ lu0 = 4.157672e-9
+ lnfactor = -4.5192e-8
+ ldif = 9e-8
+ lua = -1.9124487e-16
+ lub = 4.117038e-25
+ luc = 4.038815e-17
+ nch = 3.9e+17
+ pvoff = -4.352292e-15
+ lwl = 0.0
+ lwn = 1.0
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ pub1 = -1.8996434e-32
+ puc1 = 1.3569954e-23
+ pa0 = -1.0015934e-13
+ nlx = 0.0
+ eta0 = 5e-5
+ pk1 = -1.457495e-14
+ pk2 = 2.2122807e-15
+ pvag = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ etab = -5e-5
+ peta0 = 1.3557600041489644e-16
+ vsat = 94237.97
+ wint = 3e-9
+ pu0 = 1.6856667e-15
+ pute = -3.577514e-14
+ pvsat = 1.2437262e-9
+ vth0 = 0.41548638
+ prt = 0
+ pua = 4.758471e-23
+ pub = -5.695533e-32
+ puc = -9.239189e-24
+ lpdiblc2 = 3.0196912e-9
+ wketa = 2.8803285e-10
+ rdsw = 170.0
+ pvth0 = -9.869192e-15
+ wkt1 = 6.625341e-10
+ wkt2 = -8.725676e-11
+ drout = 0.0
+ lint = 1e-8
+ rsh = 6.8
+ tpbsw = 0.001554306
+ wmax = 1.2e-6
+ tcj = 0.001040287
+ ua1 = 1.224e-9
+ ub1 = -1.5338095e-18
+ uc1 = -7.316409e-11
+ wmin = 5e-7
+ lkt1 = -3.0828107e-9
+ lkt2 = -3.866881e-9
+ tpb = 0.001554306
+ tox = 4.08e-9
+ cjswg = 3.17352e-10
+ lmax = 1e-5
+ wa0 = 8.672666e-8
+ lmin = 1.2e-6
+ ute = -1.6080947
+ mjswg = 0.43879
+ wk1 = -1.9283881e-8
+ wk2 = 4.698517e-9
+ wln = 1.0
+ wu0 = 8.670528e-10
+ wvoff = 2.938435e-10
+ wua = 1.3831368e-16
+ wub = -1.4839938e-25
+ wuc = -1.3213606e-17
+ wwl = 0.0
+ wwn = 1
+ xti = 3
+ a0 = 0.324591
+ a1 = 0.0
+ a2 = 0.99
+ b0 = 0.0
+ b1 = 0.0
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ wub1 = -5.768295e-27
+ wuc1 = -1.6068998e-17
+ weta0 = 0
+ at = 20000.0
+ cf = 0
+ cj = 0.0009502527
+ ef = 0.874
+ k1 = 0.5600169
+ k2 = -0.005545271300000001
+ k3 = 0.0
+ em = 30000000.0
+ hdif = 2e-7
+ wvsat = -0.00012487893
+ js = 3.5e-7
+ pscbe1 = 173636400.0
+ pscbe2 = 1e-6
+ ll = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ u0 = 0.03663534
+ pb = 0.6882682
+ lub1 = 3.243357e-25
+ lpclm = 2.9892766e-7
+ wvth0 = -9.50981e-9
+ luc1 = 4.341489e-17
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ wute = 4.195195e-8
+ ua = -8.874397e-10
+ ub = 2.2584638e-18
+ uc = 1.0315766e-10
+ mjsw = 0.2003879
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ )

.model nch_fs_11 nmos (
+ level = 49
+ lvoff = 1.2067069999999999e-8
+ wcit = 5.431231e-13
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ ags = 0.02
+ beta0 = 11.59263
+ leta0 = 3.544583009680917e-10
+ lcit = 3.0283653e-10
+ cit = -0.0001583405
+ letab = -3.81143e-11
+ voff = -0.14885098
+ ldif = 9e-8
+ lvsat = -0.0007659488
+ dlc = 3e-9
+ kt1l = 0.0
+ mobmod = 1
+ prwb = 0.0
+ lvth0 = 7.488615e-9
+ prwg = 0.0
+ pub1 = -5.874811e-31
+ puc1 = -3.67348e-23
+ a0 = -0.1914371
+ a1 = 0.0
+ a2 = 0.99
+ k3b = 0.0
+ b0 = 0.0
+ b1 = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ eta0 = 1.7142847e-5
+ at = 20000.0
+ cf = 0
+ cj = 0.0009502527
+ ef = 0.874
+ k1 = 0.5552615
+ ppclm = 7.308824e-14
+ k2 = -0.0036859210000000004
+ k3 = 0.0
+ em = 30000000.0
+ pvag = 0.0
+ etab = -1.7142847e-5
+ delta = 0.01
+ js = 3.5e-7
+ vsat = 89552.49
+ ll = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ u0 = 0.03761954
+ pb = 0.6882682
+ wint = 3e-9
+ pute = -2.0303331e-13
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ua = -1.3333591e-9
+ ub = 2.969086e-18
+ uc = 1.6160392e-10
+ vth0 = 0.46359908
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ rdsw = 170.0
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ wkt1 = 1.1898274e-8
+ wkt2 = 2.0987987e-9
+ lint = 1e-8
+ wmax = 1.2e-6
+ la0 = 4.013388e-7
+ wmin = 5e-7
+ lkt1 = 9.329063e-9
+ lkt2 = 2.691467e-9
+ jsw = 1.45e-12
+ lk1 = 1.6028618e-8
+ kt1 = -0.2417087
+ lk2 = -1.1182256000000001e-8
+ kt2 = -0.03434246
+ lmax = 1.2e-6
+ llc = -0.039
+ lln = -1
+ lu0 = 3.0160021e-9
+ lmin = 5e-7
+ lua = 3.260216e-16
+ lub = -4.12618e-25
+ luc = -2.7409531e-17
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ pketa = 1.4501565e-15
+ pa0 = 1.1848049e-14
+ nlx = 0.0
+ pk1 = 7.144098e-15
+ pk2 = -4.137203e-15
+ pu0 = -1.1138246e-15
+ wpclm = 3.172275e-8
+ wub1 = 4.843047e-25
+ prt = 0
+ wuc1 = 2.7297169e-17
+ pua = -1.3255767e-22
+ pub = 5.546348e-32
+ puc = -6.669366e-24
+ tcjswg = 0.000645489
+ hdif = 2e-7
+ tcjsw = 0.000645489
+ rsh = 6.8
+ lub1 = 4.951269e-25
+ luc1 = 6.070172e-17
+ tcj = 0.001040287
+ ua1 = 1.224e-9
+ ub1 = -1.6810433e-18
+ uc1 = -8.806652e-11
+ wute = 1.8614003e-7
+ mjsw = 0.2003879
+ pvoff = 3.7090935e-15
+ tpb = 0.001554306
+ tox = 4.08e-9
+ wa0 = -9.831444e-9
+ lute = 2.2508574e-7
+ ute = -1.8126432
+ wk1 = -3.80072e-8
+ wk2 = 1.0172209e-8
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 1.3557600041489644e-16
+ wln = 1.0
+ wu0 = 3.280407e-9
+ wua = 2.9360883e-16
+ pvsat = 4.380818e-12
+ wub = -2.4531215e-25
+ wuc = -1.542897e-17
+ wwl = 0.0
+ wwn = 1
+ cdsc = 0.0
+ wketa = -1.5510503e-9
+ pvth0 = -3.2494082e-15
+ xti = 3
+ drout = 0.0
+ cgdo = 3.665e-10
+ tpbsw = 0.001554306
+ cgso = 3.665e-10
+ cjswg = 3.17352e-10
+ nfactor = 1.0
+ mjswg = 0.43879
+ pnfactor = 0.0
+ cjsw = 1.93852e-10
+ wnfactor = 0.0
+ wvoff = -6.655627e-9
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ weta0 = 0
+ pscbe1 = 400000100.0
+ pscbe2 = 1e-6
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0011219129
+ pdiblcb = 0.01
+ wvsat = 0.0009435224
+ ppdiblc2 = 1.2928064e-16
+ tnom = 25.0
+ lpclm = 9.659676e-8
+ wvth0 = -1.5216522e-8
+ wpdiblc2 = -1.1144895e-10
+ lnfactor = -4.5192e-8
+ nqsmod = 0
+ tpbswg = 0.001554306
+ toxm = 4.08e-9
+ noimod = 2
+ pcit = -2.4980728e-19
+ binunit = 2
+ pbsw = 0.6882682
+ pclm = 0.9444105
+ lpdiblc2 = 2.1785818e-9
+ lketa = -2.9090079e-9
+ xpart = 1
+ pkt1 = -5.199821e-15
+ pkt2 = -1.5611203e-15
+ keta = -0.017824383
+ pbswg = 0.6882682
+ dsub = 0.0
+ capmod = 3
+ version = 3.24
+ )

.model nch_fs_12 nmos (
+ level = 49
+ tpb = 0.001554306
+ tox = 4.08e-9
+ wa0 = 1.7605426e-7
+ pketa = -7.367843e-16
+ cjsw = 1.93852e-10
+ nfactor = 1.0
+ ute = -1.2073984
+ wk1 = -1.7855582e-8
+ wk2 = 1.6966123e-9
+ tcjswg = 0.000645489
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ wln = 1.0
+ wu0 = -4.268465e-11
+ wpclm = 1.9327061e-7
+ wua = -1.9101984e-17
+ wub = -5.11281e-26
+ wuc = -9.012729e-18
+ wwl = 0.0
+ wwn = 1
+ xti = 3
+ tcjsw = 0.000645489
+ tnom = 25.0
+ pdiblc1 = 1e-6
+ pdiblc2 = -0.00401322
+ pags = 1.8981756e-15
+ pdiblcb = 0.01
+ pvoff = -1.3169074e-15
+ toxm = 4.08e-9
+ pcit = -1.4232223e-17
+ pbsw = 0.6882682
+ pclm = 0.9948969
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 1.2420400941489644e-16
+ petab = 1.3954016e-17
+ binunit = 2
+ pvsat = 1.606088e-11
+ wketa = 3.203169e-9
+ pvth0 = 4.495999999999906e-18
+ drout = 0.0
+ tpbsw = 0.001554306
+ a0 = 0.5005398
+ a1 = 0.0
+ a2 = 0.99
+ b0 = 0.0
+ b1 = 0.0
+ at = 20000.0
+ cf = 0
+ cj = 0.0009502527
+ ef = 0.874
+ k1 = 0.489967
+ k2 = 0.022067764
+ k3 = 0.0
+ em = 30000000.0
+ js = 3.5e-7
+ cjswg = 3.17352e-10
+ ll = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ u0 = 0.041613199999999996
+ pb = 0.6882682
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ua = -5.274002e-10
+ ub = 2.0039751e-18
+ uc = 7.914647e-11
+ mjswg = 0.43879
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ pkt1 = 2.3961372e-15
+ pkt2 = 8.832021e-16
+ keta = -0.027587207
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ wvoff = 4.2704619999999996e-9
+ wags = -4.12647e-9
+ dsub = 0.0
+ pscbe1 = 400000000.0
+ pscbe2 = 1e-6
+ weta0 = 2.4721704e-11
+ lags = -9.594464e-9
+ wetab = -3.0334849e-11
+ wcit = 3.093965e-11
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ wvsat = 0.000918131
+ version = 3.24
+ nqsmod = 0
+ lpclm = 7.337301e-8
+ wvth0 = -2.2290227000000003e-8
+ tpbswg = 0.001554306
+ noimod = 2
+ lcit = 1.2733804e-10
+ voff = -0.12370098000000002
+ ldif = 9e-8
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ pub1 = 1.6165291e-31
+ puc1 = 2.0250814e-23
+ eta0 = -0.00031223928
+ pvag = 0.0
+ etab = 0.0014101875
+ vsat = 88351.66
+ wint = 3e-9
+ pute = 4.383575e-14
+ vth0 = 0.47062918
+ rdsw = 170.0
+ wkt1 = -4.614678e-9
+ wkt2 = -3.214946e-9
+ lint = 1e-8
+ wmax = 1.2e-6
+ ags = 0.04085753
+ lketa = 1.5818911e-9
+ wmin = 5e-7
+ lkt1 = 1.6202869e-9
+ lkt2 = -8.228257e-11
+ lmax = 5e-7
+ xpart = 1
+ cit = 0.00022317801
+ lmin = 1.8e-7
+ pnfactor = 0.0
+ dlc = 3e-9
+ wnfactor = 0.0
+ k3b = 0.0
+ capmod = 3
+ dwb = 0.0
+ dwg = 0.0
+ pbswg = 0.6882682
+ lvoff = 4.980705000000001e-10
+ wub1 = -1.1442477e-24
+ wuc1 = -9.658459e-17
+ ppdiblc2 = 3.905237e-16
+ hdif = 2e-7
+ beta0 = 11.59263
+ wpdiblc2 = -6.793707e-10
+ lub1 = -6.558089e-26
+ leta0 = 5.059740609680917e-10
+ luc1 = -7.416688e-18
+ wute = -3.505318e-7
+ mobmod = 1
+ la0 = 8.302936e-8
+ letab = -6.946862e-10
+ lnfactor = -4.5192e-8
+ mjsw = 0.2003879
+ lvsat = -0.00021356932
+ jsw = 1.45e-12
+ lk1 = 4.606408e-8
+ kt1 = -0.2249505
+ lk2 = -2.3028953000000002e-8
+ kt2 = -0.028312566
+ lvth0 = 4.254808999999999e-9
+ llc = -0.039
+ lln = -1
+ lute = -5.332685e-8
+ lu0 = 1.1789145e-9
+ lua = -4.471944e-17
+ lub = 3.1333025e-26
+ luc = 1.0520902e-17
+ ppclm = -1.2237712e-15
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ delta = 0.01
+ pa0 = -7.365936e-14
+ nlx = 0.0
+ lpdiblc2 = 4.540744e-9
+ cdsc = 0.0
+ pk1 = -2.1256446e-15
+ pk2 = -2.3842633e-16
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ pu0 = 4.147977e-16
+ cgdo = 3.665e-10
+ prt = 0
+ pua = 1.1289303e-23
+ pub = -3.386118e-32
+ puc = -9.620837e-24
+ cgso = 3.665e-10
+ rsh = 6.8
+ tcj = 0.001040287
+ ua1 = 1.224e-9
+ ub1 = -4.621132e-19
+ uc1 = 6.001696e-11
+ )

.model nch_fs_13 nmos (
+ level = 49
+ drout = 0.0
+ wkt1 = 5.128653e-9
+ wkt2 = 3.532295e-9
+ tpbsw = 0.001554306
+ lint = 1e-8
+ wmax = 5e-7
+ wmin = 2.2e-7
+ cjswg = 3.17352e-10
+ lmax = 2.0001e-5
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ mjswg = 0.43879
+ lmin = 1e-5
+ pscbe1 = 200000030.0
+ pscbe2 = 1e-6
+ wvoff = -1.0949902e-9
+ weta0 = 0
+ nqsmod = 0
+ wub1 = -4.432931e-26
+ wuc1 = -1.7086574e-17
+ tpbswg = 0.001554306
+ wvsat = 0.0
+ noimod = 2
+ hdif = 2e-7
+ wvth0 = -2.1421089000000002e-8
+ ags = 0.02
+ wute = 2.5547985e-8
+ mjsw = 0.2003879
+ cit = -9.999998e-5
+ dlc = 3e-9
+ k3b = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ cdsc = 0.0
+ cgdo = 3.665e-10
+ cgso = 3.665e-10
+ xpart = 1
+ jsw = 1.45e-12
+ capmod = 3
+ kt1 = -0.238767
+ lk2 = -3.6153600000000002e-9
+ kt2 = -0.03620588
+ llc = -0.039
+ cjsw = 1.93852e-10
+ lln = -1
+ a0 = 0.352982
+ a1 = 0.0
+ a2 = 0.99
+ lu0 = 4.5192000000000003e-10
+ b0 = 0.0
+ b1 = 0.0
+ pbswg = 0.6882682
+ nch = 3.9e+17
+ at = 20000.0
+ cf = 0
+ cj = 0.0009502527
+ lwl = 0.0
+ lwn = 1.0
+ ef = 0.874
+ k1 = 0.5220979
+ k2 = 0.009311849
+ k3 = 0.0
+ em = 30000000.0
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ nfactor = 1.0
+ js = 3.5e-7
+ ll = 0.0
+ nlx = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ lvoff = 9.038400000000001e-10
+ u0 = 0.0371451
+ pb = 0.6882682
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ua = -5.860608e-10
+ ub = 1.7266676e-18
+ uc = 7.252202e-11
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ mobmod = 1
+ beta0 = 11.59263
+ pu0 = 0.0
+ tnom = 25.0
+ leta0 = 3.163440009680917e-10
+ prt = 0
+ toxm = 4.08e-9
+ rsh = 6.8
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0006999999
+ lvth0 = -2.621136e-9
+ tcj = 0.001040287
+ ua1 = 1.224e-9
+ ub1 = -1.4270478e-18
+ uc1 = -6.39873e-11
+ pdiblcb = 0.01
+ pbsw = 0.6882682
+ pclm = 0.7999999
+ tpb = 0.001554306
+ tox = 4.08e-9
+ delta = 0.01
+ wa0 = 5.286186e-8
+ ute = -1.5833832
+ wk1 = -1.4938487e-9
+ wk2 = -2.6871128e-9
+ dvt0w = 0.0
+ dvt1w = 0.0
+ wln = 1.0
+ dvt2w = 0.0
+ wu0 = 9.682726e-10
+ binunit = 2
+ wua = -1.5275344e-17
+ wub = 1.2900942e-25
+ wuc = 2.9959555e-18
+ wwl = 0.0
+ wwn = 1
+ xti = 3
+ pnfactor = 0.0
+ keta = 0.002064252
+ tcjswg = 0.000645489
+ wnfactor = 0.0
+ dsub = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ tcjsw = 0.000645489
+ lnfactor = -4.5192e-8
+ voff = -0.13474068
+ version = 3.24
+ pvoff = 9.038400000000001e-16
+ ldif = 9e-8
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ eta0 = 5e-5
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 1.3557600041489644e-16
+ pvag = 0.0
+ etab = -5e-5
+ vsat = 93615.35
+ wint = 3e-9
+ vth0 = 0.44476208
+ wketa = -2.9874625e-10
+ pvth0 = -2.71152e-15
+ rdsw = 170.0
+ )

.model nch_fs_14 nmos (
+ level = 49
+ la0 = -2.4964379e-7
+ pcit = 1.5653096e-18
+ pbsw = 0.6882682
+ pclm = 0.7606163
+ jsw = 1.45e-12
+ lk1 = -6.331243e-8
+ kt1 = -0.2407974
+ lk2 = 1.7183372000000002e-8
+ kt2 = -0.03589625
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0003968183
+ pdiblcb = 0.01
+ lpscbe1 = 262.58182
+ llc = -0.039
+ lln = -1
+ lu0 = 1.0346475000000001e-8
+ lpdiblc2 = 3.0196909e-9
+ lua = -1.2876533e-16
+ lub = 7.836163e-25
+ luc = 7.064626e-17
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ pa0 = -7.427873e-14
+ nlx = 0.0
+ pk1 = 2.1894499e-14
+ pk2 = -1.0734859e-14
+ lketa = -3.0377027e-8
+ binunit = 2
+ pu0 = -1.3716021e-15
+ capmod = 3
+ prt = 0
+ pua = 1.6719826e-23
+ pub = -2.4068014e-31
+ xpart = 1
+ puc = -2.4186704e-23
+ pkt1 = -3.679308e-15
+ pkt2 = 5.879336e-16
+ rsh = 6.8
+ keta = 0.005114151
+ tcj = 0.001040287
+ ua1 = 1.224e-9
+ ub1 = -1.4513121e-18
+ uc1 = -6.991786e-11
+ pbswg = 0.6882682
+ tpb = 0.001554306
+ tox = 4.08e-9
+ dsub = 0.0
+ wa0 = 6.031956e-8
+ lvoff = -1.8823532e-8
+ mobmod = 1
+ ute = -1.5785241
+ wk1 = -3.692092e-9
+ wk2 = -1.6093152e-9
+ wcit = -1.5715551e-13
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ wln = 1.0
+ beta0 = 11.59263
+ wu0 = 1.1059835e-9
+ wua = -1.6954039e-17
+ wub = 1.5317406e-25
+ wuc = 5.42434e-18
+ leta0 = 3.163440009680917e-10
+ wwl = 0.0
+ wwn = 1
+ lcit = 2.6386249e-10
+ xti = 3
+ voff = -0.13276008
+ lvsat = -0.005267757
+ ldif = 9e-8
+ lvth0 = 5.3657104e-8
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ pub1 = 2.1839324e-32
+ puc1 = 5.837128e-24
+ version = 3.24
+ ppclm = 7.826515e-14
+ eta0 = 5e-5
+ delta = 0.01
+ pvag = 0.0
+ etab = -5e-5
+ vsat = 94144.24
+ wint = 3e-9
+ pute = -1.7889165e-14
+ vth0 = 0.43911168
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ rdsw = 170.0
+ wkt1 = 5.498062e-9
+ wkt2 = 3.473265e-9
+ lint = 1e-8
+ wmax = 5e-7
+ wmin = 2.2e-7
+ lkt1 = 2.0222748e-8
+ lkt2 = -3.0839447e-9
+ lmax = 1e-5
+ tcjswg = 0.000645489
+ lmin = 1.2e-6
+ pketa = 4.776125e-16
+ wpclm = -7.857923e-9
+ wub1 = -4.652201e-26
+ wuc1 = -1.7672629e-17
+ tcjsw = 0.000645489
+ hdif = 2e-7
+ lub1 = 2.4167225e-25
+ a0 = 0.3780467
+ a1 = 0.0
+ a2 = 0.99
+ luc1 = 5.906839e-17
+ b0 = 0.0
+ b1 = 0.0
+ wute = 2.7344081e-8
+ mjsw = 0.2003879
+ at = 20000.0
+ pvoff = 3.6135329e-15
+ cf = 0
+ cj = 0.0009502527
+ ef = 0.874
+ k1 = 0.5284545
+ k2 = 0.007223622
+ k3 = 0.0
+ em = 30000000.0
+ js = 3.5e-7
+ ll = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ u0 = 0.03615168
+ pb = 0.6882682
+ w0 = 0.0
+ rd = 0
+ lute = -4.839696e-8
+ rs = 0
+ ua = -5.731325e-10
+ ub = 1.6479914e-18
+ uc = 6.542903e-11
+ cdscb = 0.0
+ cdscd = 0.0
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -2e-8
+ ww = 0.0
+ peta0 = 1.3557600041489644e-16
+ xw = 0.0
+ pvsat = 7.826533e-10
+ wketa = -3.466991e-10
+ pvth0 = -5.1059225e-15
+ cdsc = 0.0
+ drout = 0.0
+ tpbsw = 0.001554306
+ cgdo = 3.665e-10
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ cgso = 3.665e-10
+ cjswg = 3.17352e-10
+ pscbe1 = 173636400.0
+ pscbe2 = 1e-6
+ mjswg = 0.43879
+ ags = 0.02
+ pnfactor = 0.0
+ wnfactor = 0.0
+ wvoff = -1.3670473000000001e-9
+ cjsw = 1.93852e-10
+ cit = -0.00012649217
+ nqsmod = 0
+ dlc = 3e-9
+ tpbswg = 0.001554306
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ noimod = 2
+ k3b = 0.0
+ weta0 = 0
+ dwb = 0.0
+ dwg = 0.0
+ wvsat = -7.857954e-5
+ nfactor = 1.0
+ lpclm = 3.92261e-7
+ wvth0 = -2.1180688000000003e-8
+ tnom = 25.0
+ lnfactor = -4.5192e-8
+ toxm = 4.08e-9
+ )

.model nch_fs_15 nmos (
+ level = 49
+ wub1 = -1.0574451e-25
+ wuc1 = -4.040928e-17
+ ppdiblc2 = 4.703685e-16
+ beta0 = 11.59263
+ hdif = 2e-7
+ wpdiblc2 = -4.054901e-10
+ leta0 = 3.544582809680917e-10
+ lub1 = -8.773805e-25
+ luc1 = -7.886598e-17
+ letab = -3.811428e-11
+ lnfactor = -4.5192e-8
+ wute = 1.9757099e-8
+ lvsat = -0.0007893788
+ mjsw = 0.2003879
+ lvth0 = 6.2381230000000005e-9
+ lute = -1.6751561e-7
+ ppclm = 4.863229e-14
+ delta = 0.01
+ lpdiblc2 = 1.4881204e-9
+ dvt0w = 0.0
+ cdsc = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ cgdo = 3.665e-10
+ tcjswg = 0.000645489
+ cgso = 3.665e-10
+ pketa = 3.1429577e-15
+ cjsw = 1.93852e-10
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ wpclm = 1.7687656e-8
+ tcjsw = 0.000645489
+ tnom = 25.0
+ nfactor = 1.0
+ pvoff = -4.799142e-16
+ toxm = 4.08e-9
+ ags = 0.02
+ pcit = -9.088336e-19
+ pbsw = 0.6882682
+ pclm = 0.9728217
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 1.3557600041489644e-16
+ pvsat = 1.5955267e-11
+ cit = -0.00016124053
+ wketa = -2.6444102e-9
+ pvth0 = -2.63166535e-15
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0017171376
+ dlc = 3e-9
+ drout = 0.0
+ pdiblcb = 0.01
+ k3b = 0.0
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ tpbsw = 0.001554306
+ dwb = 0.0
+ dwg = 0.0
+ pscbe1 = 400000100.0
+ pscbe2 = 1e-6
+ cjswg = 3.17352e-10
+ mjswg = 0.43879
+ binunit = 2
+ pkt1 = -1.1651986e-14
+ pkt2 = -1.4582807e-15
+ keta = -0.015611105
+ nqsmod = 0
+ wvoff = 2.1617860000000002e-9
+ tpbswg = 0.001554306
+ la0 = 2.7901473e-7
+ noimod = 2
+ jsw = 1.45e-12
+ dsub = 0.0
+ lk1 = 6.936774e-8
+ kt1 = -0.2426658
+ lk2 = -3.5143967e-8
+ kt2 = -0.04069558
+ llc = -0.039
+ lln = -1
+ weta0 = 0
+ lu0 = -1.2926906e-9
+ lua = 6.135559e-17
+ lub = -2.9489129e-25
+ luc = -2.7169401e-17
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ wvsat = 0.0005823669
+ wcit = 1.975718e-12
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ pa0 = 7.227613e-14
+ nlx = 0.0
+ lpclm = 1.4610272e-7
+ wvth0 = -2.3313668000000003e-8
+ pk1 = -1.920543e-14
+ pk2 = 7.699883e-15
+ lcit = 3.0417063e-10
+ voff = -0.16670008
+ pu0 = 1.0146696e-15
+ ldif = 9e-8
+ prt = 0
+ pua = -1.8126578e-24
+ pub = -2.6935e-33
+ puc = -6.78799e-24
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ pub1 = 9.053745e-32
+ puc1 = 3.221165e-23
+ eta0 = 1.7142866e-5
+ rsh = 6.8
+ pvag = 0.0
+ etab = -1.7142866e-5
+ tcj = 0.001040287
+ ua1 = 1.224e-9
+ ub1 = -4.866116e-19
+ uc1 = 4.899104e-11
+ vsat = 90283.57
+ version = 3.24
+ a0 = -0.07769345
+ wint = 3e-9
+ a1 = 0.0
+ a2 = 0.99
+ pute = -9.088265e-15
+ b0 = 0.0
+ b1 = 0.0
+ tpb = 0.001554306
+ vth0 = 0.47999008
+ tox = 4.08e-9
+ at = 20000.0
+ cf = 0
+ cj = 0.0009502527
+ ef = 0.874
+ k1 = 0.4140751
+ k2 = 0.052333399999999995
+ k3 = 0.0
+ rdsw = 170.0
+ wa0 = -6.602082e-8
+ em = 30000000.0
+ js = 3.5e-7
+ wkt1 = 1.2371058e-8
+ wkt2 = 5.237243e-9
+ ute = -1.4758356
+ ll = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ lint = 1e-8
+ u0 = 0.04618544
+ pb = 0.6882682
+ wk1 = 3.173889e-8
+ wk2 = -1.7501334e-8
+ w0 = 0.0
+ rd = 0
+ wmax = 5e-7
+ lketa = -6.33573e-9
+ capmod = 3
+ rs = 0
+ ua = -7.370299e-10
+ ub = 2.5777392e-18
+ uc = 1.4975288e-10
+ wln = 1.0
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -2e-8
+ ww = 0.0
+ wmin = 2.2e-7
+ wu0 = -9.511471e-10
+ xw = 0.0
+ lkt1 = 2.2390124e-8
+ wua = -9.777621e-19
+ lkt2 = 2.4832894e-9
+ wub = -5.19868e-26
+ wuc = -9.57455e-18
+ xpart = 1
+ wwl = 0.0
+ wwn = 1
+ lmax = 1.2e-6
+ xti = 3
+ lmin = 5e-7
+ pnfactor = 0.0
+ wnfactor = 0.0
+ pbswg = 0.6882682
+ mobmod = 1
+ lvoff = 2.0546844000000002e-8
+ )

.model nch_fs_16 nmos (
+ level = 49
+ at = 20000.0
+ cf = 0
+ cj = 0.0009502527
+ ef = 0.874
+ k1 = 0.4942783
+ k2 = 0.016287533
+ k3 = 0.0
+ em = 30000000.0
+ pketa = -1.9609824e-16
+ pkt1 = 3.435378e-15
+ pkt2 = -8.505888e-17
+ wnfactor = 0.0
+ keta = -0.030443965
+ js = 3.5e-7
+ ll = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ ags = 0.0548038
+ u0 = 0.03891118
+ pb = 0.6882682
+ w0 = 0.0
+ binunit = 2
+ rd = 0
+ rs = 0
+ ua = -6.614348e-10
+ ub = 2.1301375e-18
+ uc = 1.2526492e-10
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ wags = -1.1015922e-8
+ xl = -2e-8
+ ww = 0.0
+ dsub = 0.0
+ xw = 0.0
+ wpclm = 1.2379924e-7
+ cit = 0.00029138371
+ lags = -1.6009743e-8
+ dlc = 3e-9
+ wcit = -2.7539906e-12
+ ppdiblc2 = -1.1422951e-16
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ tcjsw = 0.000645489
+ k3b = 0.0
+ wpdiblc2 = 8.65375e-10
+ dwb = 0.0
+ dwg = 0.0
+ lnfactor = -4.5192e-8
+ lcit = 9.596344e-11
+ pvoff = 4.069063000000001e-16
+ voff = -0.11552988
+ ldif = 9e-8
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ pub1 = -3.181536e-32
+ puc1 = -1.1609298e-23
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 1.3557600041489644e-16
+ eta0 = -0.00026219533
+ pvag = 0.0
+ etab = 0.0013487812
+ pvsat = 1.2452966e-11
+ la0 = 1.1871046e-7
+ vsat = 89015.94
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ wint = 3e-9
+ pute = -6.731688e-15
+ wketa = 4.614407e-9
+ lpdiblc2 = 5.562512e-9
+ pvth0 = -3.7536774e-15
+ jsw = 1.45e-12
+ vth0 = 0.46776328
+ lk1 = 3.247429e-8
+ kt1 = -0.1929406
+ lk2 = -1.8562871999999998e-8
+ kt2 = -0.03937921
+ drout = 0.0
+ rdsw = 170.0
+ llc = -0.039
+ lln = -1
+ tpbsw = 0.001554306
+ pscbe1 = 400000000.0
+ pscbe2 = 1e-6
+ lu0 = 2.0534652e-9
+ version = 3.24
+ wkt1 = -2.0427562e-8
+ wkt2 = 2.2519782e-9
+ lint = 1e-8
+ lua = 2.6581833e-17
+ lub = -8.899446e-26
+ luc = -1.5904941e-17
+ nch = 3.9e+17
+ wmax = 5e-7
+ lwl = 0.0
+ lwn = 1.0
+ wmin = 2.2e-7
+ pa0 = -9.128582e-14
+ nlx = 0.0
+ cjswg = 3.17352e-10
+ lkt1 = -4.834396e-10
+ lkt2 = 1.8777602e-9
+ mjswg = 0.43879
+ pk1 = 4.587708e-15
+ pk2 = -2.4446703e-15
+ lmax = 5e-7
+ nqsmod = 0
+ tpbswg = 0.001554306
+ lmin = 1.8e-7
+ noimod = 2
+ pu0 = -1.7230291e-17
+ prt = 0
+ pua = -2.3933522e-23
+ pub = 2.5580594e-32
+ puc = 3.433529e-24
+ wvoff = 2.33915e-10
+ rsh = 6.8
+ tcj = 0.001040287
+ ua1 = 1.224e-9
+ ub1 = -3.1027764e-18
+ uc1 = -2.4653823e-10
+ weta0 = 0
+ tpb = 0.001554306
+ wub1 = 1.602399e-25
+ wuc1 = 5.485366e-17
+ tox = 4.08e-9
+ wvsat = 0.0005899806
+ wa0 = 2.8954867e-7
+ hdif = 2e-7
+ lpclm = 7.125815e-8
+ wvth0 = -2.0874508000000002e-8
+ ute = -1.9466008
+ wk1 = -1.9985334e-8
+ wk2 = 4.552045e-9
+ lub1 = 3.260553e-25
+ luc1 = 5.707747e-17
+ wute = 1.4634106e-8
+ wln = 1.0
+ mjsw = 0.2003879
+ wu0 = 1.2921135e-9
+ wua = 4.711108e-17
+ wub = -1.1345223e-25
+ wuc = -3.179524e-17
+ wwl = 0.0
+ wwn = 1
+ xti = 3
+ lute = 4.90364e-8
+ cdsc = 0.0
+ capmod = 3
+ cgdo = 3.665e-10
+ lketa = 4.87385e-10
+ cgso = 3.665e-10
+ xpart = 1
+ mobmod = 1
+ cjsw = 1.93852e-10
+ pbswg = 0.6882682
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ lvoff = -2.9914309999999998e-9
+ beta0 = 11.59263
+ leta0 = 4.829538409680917e-10
+ tnom = 25.0
+ letab = -6.664392e-10
+ lvsat = -0.00020626588
+ pags = 5.067323e-15
+ lvth0 = 1.1862447e-8
+ toxm = 4.08e-9
+ nfactor = 1.0
+ pcit = 1.266836e-18
+ ppclm = -1.7902992e-16
+ pbsw = 0.6882682
+ pclm = 1.1355271
+ delta = 0.01
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ tcjswg = 0.000645489
+ pdiblc1 = 1e-6
+ pdiblc2 = -0.007140237
+ pdiblcb = 0.01
+ a0 = 0.270794
+ a1 = 0.0
+ a2 = 0.99
+ b0 = 0.0
+ b1 = 0.0
+ pnfactor = 0.0
+ )

.model nch_sf_1 nmos (
+ level = 49
+ cjsw = 2.142574e-10
+ drout = 0.0
+ tpbsw = 0.001554306
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ cjswg = 3.507574e-10
+ pnfactor = 0.0
+ mjswg = 0.43879
+ wnfactor = 0.0
+ tnom = 25.0
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ wvoff = -6.32688e-10
+ pscbe1 = 200000030.0
+ pscbe2 = 1e-6
+ toxm = 4.08e-9
+ version = 3.24
+ pbsw = 0.6882682
+ pclm = 0.8000001
+ weta0 = 0
+ wvsat = 0.0
+ nqsmod = 0
+ lnfactor = 4.5192e-8
+ tpbswg = 0.001554306
+ wvth0 = 5.9653440000000004e-9
+ noimod = 2
+ ags = 0.02
+ keta = 0.009263485
+ cit = -0.00010000001
+ a0 = 0.3700794
+ a1 = 0.0
+ a2 = 0.99
+ b0 = 0.0
+ b1 = 0.0
+ dlc = 3e-9
+ dsub = 0.0
+ k3b = 0.0
+ at = 20000.0
+ cf = 0
+ cj = 0.001050279
+ ef = 0.874
+ k1 = 0.5142301
+ k2 = 0.022028564
+ k3 = 0.0
+ em = 30000000.0
+ dwb = 0.0
+ dwg = 0.0
+ js = 3.5e-7
+ ll = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ u0 = 0.04039571
+ pb = 0.6882682
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ dvt0 = 0.0
+ ua = -6.12274e-10
+ dvt1 = 0.0
+ ub = 2.3135539e-18
+ xpart = 1
+ dvt2 = 0.0
+ uc = 1.0876087e-10
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ voff = -0.14328952
+ capmod = 3
+ ldif = 9e-8
+ pbswg = 0.6882682
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ jsw = 1.45e-12
+ kt1 = -0.2240464
+ lk2 = 3.6153600000000002e-9
+ kt2 = -0.030266136
+ lvoff = -9.038400000000001e-10
+ eta0 = 5e-5
+ llc = -0.039
+ lln = -1
+ pvag = 0.0
+ etab = -5e-5
+ lu0 = -4.5192000000000003e-10
+ vsat = 86384.65
+ beta0 = 11.59263
+ nch = 3.9e+17
+ wint = 3e-9
+ lwl = 0.0
+ lwn = 1.0
+ vth0 = 0.45508482
+ leta0 = 9.680916984722288e-19
+ mobmod = 1
+ nlx = 0.0
+ rdsw = 170.0
+ lint = 1e-8
+ wmax = 0.000900001
+ lvth0 = 2.621136e-9
+ pu0 = 0.0
+ wmin = 1e-5
+ prt = 0
+ lmax = 2.0001e-5
+ delta = 0.01
+ lmin = 1e-5
+ rsh = 6.8
+ tcj = 0.001040287
+ ua1 = 1.224e-9
+ ub1 = -1.1209314e-18
+ uc1 = 1.1643822e-11
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ tpb = 0.001554306
+ tox = 4.08e-9
+ ute = -1.5799998
+ wln = 1.0
+ wu0 = 0.0
+ nfactor = 1.0
+ hdif = 2e-7
+ wwl = 0.0
+ wwn = 1
+ xti = 3
+ mjsw = 0.2003879
+ tcjswg = 0.000645489
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0006999999
+ pdiblcb = 0.01
+ tcjsw = 0.000645489
+ cdsc = 0.0
+ pvoff = -9.038400000000001e-16
+ cgdo = 3.665e-10
+ binunit = 2
+ cgso = 3.665e-10
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 4.148964422023837e-25
+ pvth0 = 2.71152e-15
+ )

.model nch_sf_2 nmos (
+ level = 49
+ wmax = 0.000900001
+ wmin = 1e-5
+ lkt2 = -4.553491e-12
+ lmax = 1e-5
+ lmin = 1.2e-6
+ la0 = -3.496093e-7
+ jsw = 1.45e-12
+ kt1 = -0.2240468
+ lk1 = 1.4908844e-8
+ kt2 = -0.03026568
+ lk2 = -7.49802e-9
+ llc = -0.039
+ lln = -1
+ lketa = -4.320781e-8
+ lu0 = 2.8398890000000003e-9
+ lua = -4.643216e-16
+ lub = 7.375677e-25
+ luc = 3.898355e-17
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ xpart = 1
+ pnfactor = 0.0
+ nlx = 0.0
+ hdif = 2e-7
+ wnfactor = 0.0
+ capmod = 3
+ lub1 = 4.527317e-28
+ luc1 = 7.827772e-20
+ nfactor = 1.0
+ pu0 = 0.0
+ mjsw = 0.2003879
+ prt = 0
+ pbswg = 0.6882682
+ lute = -5.743953e-11
+ lvoff = -1.1375168e-8
+ rsh = 6.8
+ tcj = 0.001040287
+ ua1 = 1.224e-9
+ ub1 = -1.1209769e-18
+ uc1 = 1.1635963e-11
+ mobmod = 1
+ beta0 = 11.59263
+ tpb = 0.001554306
+ tox = 4.08e-9
+ lnfactor = 4.5192e-8
+ leta0 = 9.680916984722288e-19
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0003968181
+ cdsc = 0.0
+ pdiblcb = 0.01
+ lpscbe1 = 262.58185
+ ute = -1.5799941
+ lvsat = -0.006562638
+ cgdo = 3.665e-10
+ wln = 1.0
+ lvth0 = 6.3234006e-8
+ wu0 = 0.0
+ wwl = 0.0
+ wwn = 1
+ cgso = 3.665e-10
+ xti = 3
+ delta = 0.01
+ lpdiblc2 = 3.0196912e-9
+ binunit = 2
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ cjsw = 2.142574e-10
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ tnom = 25.0
+ tcjswg = 0.000645489
+ a0 = 0.4051808
+ a1 = 0.0
+ a2 = 0.99
+ b0 = 0.0
+ b1 = 0.0
+ at = 20000.0
+ cf = 0
+ cj = 0.001050279
+ ef = 0.874
+ k1 = 0.5127332
+ k2 = 0.023144367
+ k3 = 0.0
+ em = 30000000.0
+ toxm = 4.08e-9
+ js = 3.5e-7
+ ll = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ u0 = 0.040065210000000004
+ pb = 0.6882682
+ w0 = 0.0
+ pbsw = 0.6882682
+ rd = 0
+ pclm = 0.7736172
+ rs = 0
+ ua = -5.656554e-10
+ ub = 2.2395009e-18
+ uc = 1.0484686e-10
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ tcjsw = 0.000645489
+ version = 3.24
+ pvoff = -9.038400000000001e-16
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 4.148964422023837e-25
+ pvth0 = 2.71152e-15
+ keta = 0.013601619
+ drout = 0.0
+ tpbsw = 0.001554306
+ dsub = 0.0
+ cjswg = 3.507574e-10
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ mjswg = 0.43879
+ pscbe1 = 173636400.0
+ pscbe2 = 1e-6
+ lcit = 2.6652053e-10
+ wvoff = -6.32688e-10
+ voff = -0.14223822
+ ldif = 9e-8
+ ags = 0.02
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ weta0 = 0
+ nqsmod = 0
+ eta0 = 5e-5
+ tpbswg = 0.001554306
+ pvag = 0.0
+ etab = -5e-5
+ cit = -0.00012675911
+ noimod = 2
+ wvsat = 0.0
+ vsat = 87043.55
+ wint = 3e-9
+ dlc = 3e-9
+ lpclm = 2.6277317e-7
+ wvth0 = 5.9653440000000004e-9
+ vth0 = 0.44899922
+ k3b = 0.0
+ rdsw = 170.0
+ dwb = 0.0
+ dwg = 0.0
+ lint = 1e-8
+ )

.model nch_sf_3 nmos (
+ level = 49
+ beta0 = 11.59263
+ leta0 = 3.8114280968091696e-11
+ letab = -3.811428e-11
+ lvsat = -0.0007622857
+ version = 3.24
+ lvth0 = 6.563892999999999e-9
+ delta = 0.01
+ keta = -0.015927497
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ dsub = 0.0
+ pnfactor = 0.0
+ lags = -3.044698e-8
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ tcjswg = 0.000645489
+ wnfactor = 0.0
+ lcit = 3.0262734e-10
+ voff = -0.16483012
+ ldif = 9e-8
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ eta0 = 1.7142866e-5
+ pvag = 0.0
+ etab = -1.7142866e-5
+ vsat = 82043.24
+ tcjsw = 0.000645489
+ lnfactor = 4.5192e-8
+ wint = 3e-9
+ vth0 = 0.49785271999999997
+ rdsw = 170.0
+ pvoff = -9.038400000000001e-16
+ lint = 1e-8
+ wmax = 0.000900001
+ wmin = 1e-5
+ cdscb = 0.0
+ cdscd = 0.0
+ lkt1 = 5.782678e-9
+ lkt2 = 1.5570838e-9
+ peta0 = 4.148964422023837e-25
+ lmax = 1.2e-6
+ lpdiblc2 = 1.525682e-9
+ lmin = 5e-7
+ pvth0 = 2.71152e-15
+ ags = 0.0462474
+ drout = 0.0
+ tpbsw = 0.001554306
+ cit = -0.00015788565
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ dlc = 3e-9
+ cjswg = 3.507574e-10
+ k3b = 0.0
+ pscbe1 = 400000100.0
+ pscbe2 = 1e-6
+ mjswg = 0.43879
+ dwb = 0.0
+ dwg = 0.0
+ hdif = 2e-7
+ lua1 = -3.0446746e-18
+ lub1 = -1.2004175e-24
+ luc1 = -6.517273e-17
+ wvoff = -6.32688e-10
+ mjsw = 0.2003879
+ nqsmod = 0
+ tpbswg = 0.001554306
+ noimod = 2
+ nfactor = 1.0
+ lute = -2.6630502e-7
+ weta0 = 0
+ la0 = 4.581426e-7
+ wvsat = 0.0
+ jsw = 1.45e-12
+ kt1 = -0.2290285
+ lk1 = -7.214246e-9
+ kt2 = -0.031611919
+ lk2 = 5.318511e-9
+ lpclm = 1.5245718e-7
+ wvth0 = 5.9653440000000004e-9
+ a0 = -0.2911571
+ a1 = 0.0
+ a2 = 0.99
+ b0 = 0.0
+ b1 = 0.0
+ llc = -0.039
+ cdsc = 0.0
+ lln = -1
+ lu0 = 5.886878999999999e-10
+ at = 20000.0
+ cf = 0
+ cj = 0.001050279
+ ef = 0.874
+ k1 = 0.5318048
+ k2 = 0.012095633000000001
+ k3 = 0.0
+ em = 30000000.0
+ lua = 7.982966e-17
+ lub = -1.5630905e-25
+ luc = -9.669895e-18
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ js = 3.5e-7
+ cgdo = 3.665e-10
+ ll = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0016847569
+ u0 = 0.0420059
+ pb = 0.6882682
+ w0 = 0.0
+ rd = 0
+ nlx = 0.0
+ rs = 0
+ pdiblcb = 0.01
+ ua = -1.0347512e-9
+ ub = 3.0100842e-18
+ uc = 1.4678947e-10
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ cgso = 3.665e-10
+ pu0 = 0.0
+ prt = 0
+ cjsw = 2.142574e-10
+ binunit = 2
+ rsh = 6.8
+ tcj = 0.001040287
+ ua1 = 1.2266247e-9
+ ub1 = -8.574386e-20
+ uc1 = 6.788683e-11
+ lketa = -8.954029e-9
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ tpb = 0.001554306
+ tox = 4.08e-9
+ capmod = 3
+ xpart = 1
+ ute = -1.3504703
+ tnom = 25.0
+ wln = 1.0
+ wu0 = 0.0
+ pbswg = 0.6882682
+ wwl = 0.0
+ wwn = 1
+ xti = 3
+ toxm = 4.08e-9
+ mobmod = 1
+ lvoff = 1.4831418000000001e-8
+ pbsw = 0.6882682
+ pclm = 0.8687172
+ )

.model nch_sf_4 nmos (
+ level = 49
+ lua1 = 8.039099e-19
+ lub1 = 3.824101e-25
+ luc1 = 2.9606131e-17
+ mjsw = 0.2003879
+ lute = 7.030476e-8
+ ags = -0.019916179
+ tcjsw = 0.000645489
+ nfactor = 1.0
+ cdsc = 0.0
+ cit = 0.000271889
+ pvoff = -9.038400000000001e-16
+ dlc = 3e-9
+ cgdo = 3.665e-10
+ k3b = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cgso = 3.665e-10
+ peta0 = 4.148964422023837e-25
+ pdiblc1 = 1e-6
+ pdiblc2 = -0.00593541
+ pdiblcb = 0.01
+ pvth0 = 2.71152e-15
+ drout = 0.0
+ alpha0 = 0.0
+ cjsw = 2.142574e-10
+ alpha1 = 0.448150714
+ tpbsw = 0.001554306
+ la0 = 7.545271e-8
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ pscbe1 = 400000000.0
+ pscbe2 = 1e-6
+ binunit = 2
+ jsw = 1.45e-12
+ kt1 = -0.22715
+ lk1 = 4.899558e-8
+ kt2 = -0.029537767
+ lk2 = -1.9725976e-8
+ cjswg = 3.507574e-10
+ pnfactor = 0.0
+ llc = -0.039
+ lln = -1
+ mjswg = 0.43879
+ lu0 = 7.998789e-10
+ wnfactor = 0.0
+ lua = -1.0530929e-18
+ lub = 5.559478e-27
+ luc = 4.133919e-18
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ tnom = 25.0
+ nqsmod = 0
+ tpbswg = 0.001554306
+ wvoff = -6.32688e-10
+ nlx = 0.0
+ noimod = 2
+ toxm = 4.08e-9
+ pu0 = 0.0
+ weta0 = 0
+ pbsw = 0.6882682
+ pclm = 1.1076791
+ prt = 0
+ wvsat = 0.0
+ lnfactor = 4.5192e-8
+ lpclm = 4.253467e-8
+ wvth0 = 5.9653440000000004e-9
+ rsh = 6.8
+ tcj = 0.001040287
+ ua1 = 1.2182583e-9
+ ub1 = -3.526674e-18
+ uc1 = -1.381542e-10
+ tpb = 0.001554306
+ tox = 4.08e-9
+ ute = -2.0822308
+ version = 3.24
+ wln = 1.0
+ wu0 = 0.0
+ lpdiblc2 = 5.030957e-9
+ wwl = 0.0
+ wwn = 1
+ xti = 3
+ keta = -0.04182327
+ capmod = 3
+ dsub = 0.0
+ lketa = 2.9580252e-9
+ xpart = 1
+ lags = -1.1735286e-11
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ lcit = 1.0493098e-10
+ voff = -0.12726132
+ pbswg = 0.6882682
+ mobmod = 1
+ ldif = 9e-8
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ lvoff = -2.4502018000000002e-9
+ eta0 = -0.0002937502
+ pvag = 0.0
+ etab = 0.0013875004
+ beta0 = 11.59263
+ vsat = 80823.6
+ wint = 3e-9
+ leta0 = 1.811250609680917e-10
+ vth0 = 0.49375982
+ letab = -6.842502e-10
+ rdsw = 170.0
+ lvsat = -0.00020125005
+ lint = 1e-8
+ lvth0 = 8.446637e-9
+ wmax = 0.000900001
+ wmin = 1e-5
+ lkt1 = 4.918561e-9
+ lkt2 = 6.029743e-10
+ delta = 0.01
+ lmax = 5e-7
+ a0 = 0.5407774
+ a1 = 0.0
+ a2 = 0.99
+ b0 = 0.0
+ b1 = 0.0
+ lmin = 1.8e-7
+ at = 20000.0
+ cf = 0
+ cj = 0.001050279
+ ef = 0.874
+ k1 = 0.4096095
+ k2 = 0.06654018
+ k3 = 0.0
+ em = 30000000.0
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ js = 3.5e-7
+ ll = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ u0 = 0.04154679
+ pb = 0.6882682
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ua = -8.589192e-10
+ ub = 2.6581962e-18
+ uc = 1.1678118e-10
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ tcjswg = 0.000645489
+ hdif = 2e-7
+ )

.model nch_sf_5 nmos (
+ level = 49
+ pu0 = 0.0
+ pscbe1 = 200000030.0
+ pscbe2 = 1e-6
+ tpbsw = 0.001554306
+ prt = 0
+ dsub = 0.0
+ cjswg = 3.507574e-10
+ rsh = 6.8
+ tcj = 0.001040287
+ ua1 = 1.224e-9
+ ub1 = -1.0684574e-18
+ a0 = 0.3702259
+ a1 = 0.0
+ a2 = 0.99
+ uc1 = 2.4230474e-11
+ b0 = 0.0
+ b1 = 0.0
+ mjswg = 0.43879
+ nqsmod = 0
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ tpbswg = 0.001554306
+ at = 20000.0
+ cf = 0
+ cj = 0.001050279
+ ef = 0.874
+ k1 = 0.5102321
+ k2 = 0.023322214
+ k3 = 0.0
+ tpb = 0.001554306
+ noimod = 2
+ em = 30000000.0
+ tox = 4.08e-9
+ js = 3.5e-7
+ wa0 = -1.4643313e-9
+ ll = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ wvoff = 2.5803440000000005e-10
+ u0 = 0.04122822
+ pb = 0.6882682
+ w0 = 0.0
+ rd = 0
+ ute = -1.5803809
+ rs = 0
+ ua = -5.885942e-10
+ ub = 2.3329335e-18
+ uc = 1.1057788e-10
+ voff = -0.14337861999999998
+ wk1 = 3.995606e-8
+ wk2 = -1.2928737e-8
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -2e-8
+ ww = 0.0
+ ldif = 9e-8
+ xw = 0.0
+ wln = 1.0
+ wu0 = -8.320099e-9
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ puc1 = -1.4905616e-28
+ weta0 = 0
+ wua = -2.3665659e-16
+ wub = -1.936796e-25
+ wuc = -1.815927e-17
+ wwl = 0.0
+ wwn = 1
+ eta0 = 5e-5
+ xti = 3
+ wvsat = 0.0
+ pvag = 0.0
+ etab = -5e-5
+ vsat = 86384.65
+ wvth0 = 6.652955400000001e-9
+ wint = 3e-9
+ vth0 = 0.45501602
+ rdsw = 170.0
+ wkt1 = -8.215166e-9
+ wkt2 = 1.6245854e-9
+ lint = 1e-8
+ wmax = 1e-5
+ wmin = 1.2e-6
+ lmax = 2.0001e-5
+ lmin = 1e-5
+ capmod = 3
+ xpart = 1
+ wub1 = -5.244247e-25
+ pnfactor = 0.0
+ wuc1 = -1.257911e-16
+ wnfactor = 0.0
+ hdif = 2e-7
+ mobmod = 1
+ wute = 3.808433e-9
+ pbswg = 0.6882682
+ mjsw = 0.2003879
+ lvoff = -9.038400000000001e-10
+ beta0 = 11.59263
+ lnfactor = 4.5192e-8
+ leta0 = 9.680916984722288e-19
+ cdsc = 0.0
+ nfactor = 1.0
+ lvth0 = 2.621136e-9
+ cgdo = 3.665e-10
+ cgso = 3.665e-10
+ delta = 0.01
+ dvt0w = 0.0
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0006999999
+ dvt1w = 0.0
+ dvt2w = 0.0
+ pdiblcb = 0.01
+ cjsw = 2.142574e-10
+ tcjswg = 0.000645489
+ ags = 0.02
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ cit = -0.00010000001
+ binunit = 2
+ dlc = 3e-9
+ tnom = 25.0
+ k3b = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ toxm = 4.08e-9
+ pbsw = 0.6882682
+ pclm = 0.8000001
+ tcjsw = 0.000645489
+ pvoff = -9.038400000000001e-16
+ jsw = 1.45e-12
+ kt1 = -0.2232244
+ kt2 = -0.030428693
+ lk2 = 3.6153600000000002e-9
+ llc = -0.039
+ lln = -1
+ lu0 = -4.5192000000000003e-10
+ cdscb = 0.0
+ cdscd = 0.0
+ nch = 3.9e+17
+ peta0 = 4.148964422023837e-25
+ lwl = 0.0
+ lwn = 1.0
+ nlx = 0.0
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ version = 3.24
+ wketa = -1.0935369e-8
+ pvth0 = 2.71152e-15
+ keta = 0.010357677
+ drout = 0.0
+ )

.model nch_sf_6 nmos (
+ level = 49
+ nfactor = 1.0
+ cgso = 3.665e-10
+ capmod = 3
+ cjsw = 2.142574e-10
+ lketa = -4.518989e-8
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0003968181
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ pdiblcb = 0.01
+ lpscbe1 = 262.58185
+ xpart = 1
+ mobmod = 1
+ tnom = 25.0
+ pbswg = 0.6882682
+ binunit = 2
+ toxm = 4.08e-9
+ lvoff = -1.1709891999999999e-8
+ a0 = 0.40626
+ a1 = 0.0
+ a2 = 0.99
+ b0 = 0.0
+ b1 = 0.0
+ pbsw = 0.6882682
+ pclm = 0.7755287
+ at = 20000.0
+ cf = 0
+ cj = 0.001050279
+ ef = 0.874
+ k1 = 0.508509
+ beta0 = 11.59263
+ k2 = 0.02454095
+ k3 = 0.0
+ em = 30000000.0
+ js = 3.5e-7
+ ll = 0.0
+ leta0 = 9.680916984722288e-19
+ mj = 0.3595262
+ lw = 0.0
+ u0 = 0.04092259
+ pb = 0.6882682
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ags = 0.02
+ ua = -5.377125e-10
+ ub = 2.2537915e-18
+ uc = 1.0657759e-10
+ lvsat = -0.006753025
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ lvth0 = 6.3327226e-8
+ cit = -0.00012675911
+ ppclm = 1.9027247e-13
+ delta = 0.01
+ dlc = 3e-9
+ k3b = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ tcjswg = 0.000645489
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ pkt1 = 4.710912e-15
+ pkt2 = -4.130377e-15
+ keta = 0.014894814
+ version = 3.24
+ dsub = 0.0
+ pnfactor = 0.0
+ la0 = -3.588995e-7
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ wnfactor = 0.0
+ jsw = 1.45e-12
+ lk1 = 1.7161611e-8
+ kt1 = -0.2231775
+ lk2 = -8.523252e-9
+ kt2 = -0.030469729
+ pketa = 1.9809019e-14
+ llc = -0.039
+ lln = -1
+ lu0 = 2.5921712e-9
+ lcit = 2.6652053e-10
+ voff = -0.14229371999999998
+ lua = -5.067804e-16
+ lub = 7.882536e-25
+ luc = 3.984287e-17
+ nch = 3.9e+17
+ ldif = 9e-8
+ lwl = 0.0
+ lwn = 1.0
+ wpclm = -1.9103656e-8
+ kt1l = 0.0
+ pa0 = 9.284546e-14
+ prwb = 0.0
+ prwg = 0.0
+ pub1 = 4.176128e-31
+ nlx = 0.0
+ puc1 = 7.417578e-23
+ eta0 = 5e-5
+ pk1 = -2.2514154e-14
+ pk2 = 1.0246181e-14
+ pvag = 0.0
+ etab = -5e-5
+ tcjsw = 0.000645489
+ pu0 = 2.4756895e-15
+ vsat = 87062.66
+ lnfactor = 4.5192e-8
+ wint = 3e-9
+ pute = -5.708167e-14
+ prt = 0
+ pua = 4.243342e-22
+ pub = -5.065558e-31
+ puc = -8.588134e-24
+ vth0 = 0.44892112
+ rdsw = 170.0
+ pvoff = 2.441401e-15
+ wkt1 = -8.688151e-9
+ wkt2 = 2.0392819e-9
+ rsh = 6.8
+ lint = 1e-8
+ tcj = 0.001040287
+ ua1 = 1.224e-9
+ ub1 = -1.0643074e-18
+ uc1 = 2.4967807e-11
+ wmax = 1e-5
+ wmin = 1.2e-6
+ cdscb = 0.0
+ cdscd = 0.0
+ tpb = 0.001554306
+ peta0 = 4.148964422023837e-25
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ tox = 4.08e-9
+ lkt1 = -4.674615e-10
+ lkt2 = 4.087321e-10
+ wa0 = -1.0786144e-8
+ lpdiblc2 = 3.0196912e-9
+ lmax = 1e-5
+ pvsat = 1.9027204e-9
+ ute = -1.5809486
+ pscbe1 = 173636400.0
+ pscbe2 = 1e-6
+ wk1 = 4.221652e-8
+ wk2 = -1.3957471e-8
+ lmin = 1.2e-6
+ wketa = -1.292423e-8
+ pvth0 = 1.7798325e-15
+ wln = 1.0
+ drout = 0.0
+ wu0 = -8.568663e-9
+ tpbsw = 0.001554306
+ wua = -2.7926046e-16
+ wub = -1.4282058e-25
+ wuc = -1.7297008e-17
+ wwl = 0.0
+ wwn = 1
+ xti = 3
+ nqsmod = 0
+ tpbswg = 0.001554306
+ cjswg = 3.507574e-10
+ noimod = 2
+ wub1 = -5.663537e-25
+ wuc1 = -1.3323848e-16
+ mjswg = 0.43879
+ hdif = 2e-7
+ wvoff = -7.783409999999999e-11
+ lub1 = -4.133362e-26
+ luc1 = -7.343755e-18
+ wute = 9.539526e-9
+ mjsw = 0.2003879
+ weta0 = 0
+ lute = 5.654154e-9
+ wvsat = -0.00019104627
+ lpclm = 2.4373449e-7
+ wvth0 = 6.7464942e-9
+ cdsc = 0.0
+ cgdo = 3.665e-10
+ )

.model nch_sf_7 nmos (
+ level = 49
+ beta0 = 11.59263
+ pvag = 0.0
+ etab = -1.7142869e-5
+ vsat = 81898.23
+ leta0 = 3.8114280968091696e-11
+ wint = 3e-9
+ pute = 4.357466e-13
+ letab = -3.811428e-11
+ vth0 = 0.49852362
+ lvsat = -0.0007622865
+ rdsw = 170.0
+ lvth0 = 5.788268e-9
+ wkt1 = -3.681822e-9
+ wkt2 = -1.3190541e-9
+ lint = 1e-8
+ wmax = 1e-5
+ la0 = 4.645035e-7
+ ppclm = 7.258032e-15
+ wmin = 1.2e-6
+ jsw = 1.45e-12
+ lk1 = -1.1179709e-8
+ kt1 = -0.2286601
+ lk2 = 7.0464250000000005e-9
+ kt2 = -0.031479932
+ delta = 0.01
+ tcjswg = 0.000645489
+ lkt1 = 5.892387e-9
+ lkt2 = 1.5805686e-9
+ llc = -0.039
+ lln = -1
+ lmax = 1.2e-6
+ lu0 = 5.085513000000001e-10
+ lmin = 5e-7
+ lua = 6.148926e-17
+ lub = -1.2783527e-25
+ luc = -6.505068e-18
+ nch = 3.9e+17
+ dvt0w = 0.0
+ lwl = 0.0
+ lwn = 1.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ pa0 = -6.357063e-14
+ nlx = 0.0
+ pk1 = 3.963084e-14
+ pk2 = -1.7268767e-14
+ pu0 = 8.008865e-16
+ prt = 0
+ pua = 1.8329395e-22
+ pub = -2.8456703e-31
+ puc = -3.16293e-23
+ wua1 = -3.55913e-18
+ wub1 = -1.6132161e-24
+ wuc1 = -1.8047248e-16
+ hdif = 2e-7
+ rsh = 6.8
+ pketa = 9.843987e-15
+ tcj = 0.001040287
+ ua1 = 1.2269809e-9
+ ub1 = 7.567455e-20
+ lua1 = -3.457781e-18
+ uc1 = 8.594492e-11
+ lub1 = -1.3637128e-24
+ luc1 = -7.807721e-17
+ wute = -4.153124e-7
+ mjsw = 0.2003879
+ tpb = 0.001554306
+ tox = 4.08e-9
+ wa0 = 1.2405528e-7
+ wpclm = 1.3866737e-7
+ ute = -1.3089141
+ lute = -3.0990586e-7
+ wk1 = -1.1356744e-8
+ wk2 = 9.762311e-9
+ wln = 1.0
+ tcjsw = 0.000645489
+ wu0 = -7.124867e-9
+ wua = -7.146715e-17
+ wub = -3.341902e-25
+ wuc = 2.5660584e-18
+ wwl = 0.0
+ wwn = 1
+ xti = 3
+ cdsc = 0.0
+ pvoff = -3.917654e-15
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ cgdo = 3.665e-10
+ a0 = -0.3035701
+ a1 = 0.0
+ a2 = 0.99
+ b0 = 0.0
+ b1 = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 4.148964422023837e-25
+ at = 20000.0
+ cf = 0
+ cj = 0.001050279
+ pscbe1 = 400000100.0
+ pscbe2 = 1e-6
+ ef = 0.874
+ k1 = 0.5329412
+ k2 = 0.011118815
+ k3 = 0.0
+ em = 30000000.0
+ cgso = 3.665e-10
+ js = 3.5e-7
+ ll = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ u0 = 0.04271881
+ pb = 0.6882682
+ nfactor = 1.0
+ w0 = 0.0
+ rd = 0
+ wketa = -4.333682e-9
+ rs = 0
+ ua = -1.0276002e-9
+ ub = 3.0435232e-18
+ uc = 1.4653272e-10
+ pvth0 = 1.0463117999999999e-14
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ drout = 0.0
+ tpbsw = 0.001554306
+ nqsmod = 0
+ cjsw = 2.142574e-10
+ tpbswg = 0.001554306
+ noimod = 2
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ cjswg = 3.507574e-10
+ pnfactor = 0.0
+ mjswg = 0.43879
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0017737894
+ pdiblcb = 0.01
+ wnfactor = 0.0
+ tnom = 25.0
+ wvoff = 5.40411e-9
+ pags = 4.128623e-14
+ toxm = 4.08e-9
+ weta0 = 0
+ ppdiblc2 = 1.0321563e-15
+ binunit = 2
+ pbsw = 0.6882682
+ pclm = 0.8548421
+ wvsat = 0.0014492224
+ wpdiblc2 = -8.897895e-10
+ lpclm = 1.5173094e-7
+ wvth0 = -7.390919999999996e-10
+ lnfactor = 4.5192e-8
+ capmod = 3
+ lpdiblc2 = 1.4224044e-9
+ pkt1 = -1.0964308e-15
+ pkt2 = -2.3470743e-16
+ keta = -0.01549387
+ lketa = -9.939018e-9
+ mobmod = 1
+ wags = -3.559157e-8
+ dsub = 0.0
+ version = 3.24
+ xpart = 1
+ ags = 0.04980868
+ lags = -3.457808e-8
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ cit = -0.00015788565
+ pbswg = 0.6882682
+ lcit = 3.0262734e-10
+ voff = -0.16543412
+ ldif = 9e-8
+ dlc = 3e-9
+ k3b = 0.0
+ kt1l = 0.0
+ lvoff = 1.5132981999999998e-8
+ pua1 = 4.128591e-24
+ prwb = 0.0
+ prwg = 0.0
+ pub1 = 1.6319734e-30
+ puc1 = 1.2896722e-22
+ dwb = 0.0
+ dwg = 0.0
+ eta0 = 1.7142869e-5
+ )

.model nch_sf_8 nmos (
+ level = 49
+ pketa = -2.7027957e-15
+ tnom = 25.0
+ pdiblc1 = 1e-6
+ pdiblc2 = -0.006119013
+ pdiblcb = 0.01
+ pags = -1.0838496e-14
+ toxm = 4.08e-9
+ wpclm = 6.656068e-8
+ pcit = 1.4220811e-17
+ pbsw = 0.6882682
+ pclm = 1.1010191
+ tcjsw = 0.000645489
+ binunit = 2
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ pvoff = -1.8792550000000002e-15
+ pscbe1 = 400000000.0
+ pscbe2 = 1e-6
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = -1.3821213851035578e-18
+ petab = 1.6959704e-18
+ pvsat = 1.5350395e-12
+ wketa = 2.2941933e-8
+ nqsmod = 0
+ pvth0 = 7.220458e-15
+ tpbswg = 0.001554306
+ drout = 0.0
+ noimod = 2
+ pkt1 = -1.7512235e-15
+ pkt2 = 7.382567e-17
+ keta = -0.04411884
+ tpbsw = 0.001554306
+ wags = 7.772305e-8
+ dsub = 0.0
+ cjswg = 3.507574e-10
+ mjswg = 0.43879
+ lags = 1.0727657e-9
+ wcit = -3.0914837e-11
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ version = 3.24
+ wvoff = 9.728084e-10
+ lcit = 1.0350804e-10
+ voff = -0.12742202
+ ldif = 9e-8
+ weta0 = 3.0046217e-12
+ kt1l = 0.0
+ pua1 = -1.0901051e-24
+ prwb = 0.0
+ prwg = 0.0
+ pub1 = -4.238914e-31
+ puc1 = -2.7204607e-23
+ wetab = -3.686654e-12
+ wvsat = 0.0014459029
+ eta0 = -0.00029405078
+ pvag = 0.0
+ etab = 0.0013878694
+ lpclm = 3.848953e-8
+ wvth0 = 6.3101676e-9
+ vsat = 80678.92
+ wint = 3e-9
+ pute = -1.178615e-13
+ vth0 = 0.49372532
+ rdsw = 170.0
+ capmod = 3
+ wkt1 = -2.2583577e-9
+ wkt2 = -1.9897783e-9
+ lint = 1e-8
+ ags = -0.027693154
+ wmax = 1e-5
+ wmin = 1.2e-6
+ lkt1 = 5.093789e-9
+ lkt2 = 5.955873e-10
+ lmax = 5e-7
+ cit = 0.00027498236
+ lmin = 1.8e-7
+ dlc = 3e-9
+ mobmod = 1
+ k3b = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ a0 = 0.5262308
+ a1 = 0.0
+ a2 = 0.99
+ lketa = 3.228467e-9
+ b0 = 0.0
+ b1 = 0.0
+ at = 20000.0
+ cf = 0
+ cj = 0.001050279
+ ef = 0.874
+ k1 = 0.4007356
+ k2 = 0.07041932
+ k3 = 0.0
+ em = 30000000.0
+ xpart = 1
+ js = 3.5e-7
+ ll = 0.0
+ pnfactor = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ u0 = 0.04203316
+ wua1 = 7.785862e-18
+ pb = 0.6882682
+ wub1 = 2.8560549e-24
+ w0 = 0.0
+ wuc1 = 1.5903152e-16
+ rd = 0
+ rs = 0
+ ua = -9.017296e-10
+ ub = 2.7527719e-18
+ uc = 1.2291169e-10
+ wnfactor = 0.0
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ hdif = 2e-7
+ lua1 = 9.129858e-19
+ lub1 = 4.248247e-25
+ la0 = 8.279508e-8
+ luc1 = 3.232822e-17
+ pbswg = 0.6882682
+ wute = 7.881835e-7
+ mjsw = 0.2003879
+ jsw = 1.45e-12
+ lk1 = 4.963488e-8
+ kt1 = -0.226924
+ lk2 = -2.0231804000000002e-8
+ kt2 = -0.029338669
+ llc = -0.039
+ lvoff = -2.3526017e-9
+ lln = -1
+ lu0 = 8.239492e-10
+ ppdiblc2 = -2.2121929e-16
+ lute = 8.209799e-8
+ lua = 3.588764e-18
+ lub = 5.910339e-27
+ luc = 4.360599e-18
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ wpdiblc2 = 1.8349379e-9
+ beta0 = 11.59263
+ pa0 = -7.337964e-14
+ lnfactor = 4.5192e-8
+ nlx = 0.0
+ leta0 = 1.812633409680917e-10
+ letab = -6.844199e-10
+ pk1 = -6.389182e-15
+ pk2 = 5.055259e-15
+ lvsat = -0.00020140363
+ cdsc = 0.0
+ pu0 = -2.4055863e-16
+ lvth0 = 7.995472e-9
+ prt = 0
+ pua = -4.639069e-23
+ pub = -3.506499e-33
+ puc = -2.2654354e-24
+ cgdo = 3.665e-10
+ tcjswg = 0.000645489
+ ppclm = 4.042711e-14
+ delta = 0.01
+ cgso = 3.665e-10
+ rsh = 6.8
+ tcj = 0.001040287
+ lpdiblc2 = 5.053093e-9
+ ua1 = 1.2174792e-9
+ ub1 = -3.81245e-18
+ uc1 = -1.540669e-10
+ tpb = 0.001554306
+ tox = 4.08e-9
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ wa0 = 1.4537927e-7
+ nfactor = 1.0
+ ute = -2.1610963
+ cjsw = 2.142574e-10
+ wk1 = 8.868675e-8
+ wk2 = -3.876818e-8
+ wln = 1.0
+ wu0 = -4.860856e-9
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ wua = 4.278473e-16
+ wub = -9.451913e-25
+ wuc = -6.126842e-17
+ wwl = 0.0
+ wwn = 1
+ xti = 3
+ )

.model nch_sf_9 nmos (
+ level = 49
+ cjswg = 3.507574e-10
+ mjswg = 0.43879
+ wub1 = -7.675553e-27
+ wuc1 = -1.4706552e-17
+ hdif = 2e-7
+ wvoff = -1.499257e-9
+ ags = 0.02
+ wute = 3.836007e-8
+ mjsw = 0.2003879
+ weta0 = 0
+ cit = -0.00010000004
+ wvsat = 0.0
+ dlc = 3e-9
+ k3b = 0.0
+ wvth0 = 1.7022350000000006e-9
+ dwb = 0.0
+ dwg = 0.0
+ capmod = 3
+ cdsc = 0.0
+ cgdo = 3.665e-10
+ cgso = 3.665e-10
+ mobmod = 1
+ jsw = 1.45e-12
+ kt1 = -0.2313184
+ lk2 = 3.6153600000000002e-9
+ kt2 = -0.029076951
+ llc = -0.039
+ lln = -1
+ lu0 = -4.5192000000000003e-10
+ cjsw = 2.142574e-10
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ nlx = 0.0
+ nfactor = 1.0
+ xpart = 1
+ pu0 = 0.0
+ prt = 0
+ tnom = 25.0
+ pbswg = 0.6882682
+ rsh = 6.8
+ tcj = 0.001040287
+ ua1 = 1.224e-9
+ pdiblc1 = 1e-6
+ toxm = 4.08e-9
+ pdiblc2 = 0.0007000003
+ ub1 = -1.5012456e-18
+ lvoff = -9.038400000000001e-10
+ uc1 = -6.880516e-11
+ pdiblcb = 0.01
+ pbsw = 0.6882682
+ tpb = 0.001554306
+ pclm = 0.8000001
+ tox = 4.08e-9
+ beta0 = 11.59263
+ wa0 = 7.667051e-8
+ leta0 = 9.680916984722288e-19
+ ute = -1.6093186
+ wk1 = -2.074723e-8
+ wk2 = 4.920634e-9
+ tcjswg = 0.000645489
+ wln = 1.0
+ wu0 = 1.0362965e-9
+ lvth0 = 2.621136e-9
+ binunit = 2
+ wua = 1.4309126e-16
+ wub = -1.5411778e-25
+ wuc = -1.4141237e-17
+ wwl = 0.0
+ wwn = 1
+ xti = 3
+ delta = 0.01
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ keta = 0.0010152902
+ dsub = 0.0
+ pnfactor = 0.0
+ wnfactor = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ a0 = 0.3047864
+ a1 = 0.0
+ a2 = 0.99
+ b0 = 0.0
+ b1 = 0.0
+ voff = -0.14190692
+ version = 3.24
+ at = 20000.0
+ cf = 0
+ cj = 0.001050279
+ ldif = 9e-8
+ ef = 0.874
+ k1 = 0.5610723
+ k2 = 0.0083729917
+ k3 = 0.0
+ em = 30000000.0
+ kt1l = 0.0
+ js = 3.5e-7
+ prwb = 0.0
+ ll = 0.0
+ prwg = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ u0 = 0.03339204
+ pb = 0.6882682
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ua = -9.066409e-10
+ ub = 2.2997995e-18
+ uc = 1.072127e-10
+ eta0 = 5e-5
+ wl = 0.0
+ tcjsw = 0.000645489
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -2e-8
+ ww = 0.0
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ xw = 0.0
+ pvag = 0.0
+ etab = -5e-5
+ lnfactor = 4.5192e-8
+ vsat = 86384.65
+ wint = 3e-9
+ pscbe1 = 200000030.0
+ pscbe2 = 1e-6
+ vth0 = 0.45916242
+ pvoff = -9.038400000000001e-16
+ rdsw = 170.0
+ wkt1 = 1.4490446e-9
+ wkt2 = 1.0605161e-11
+ lint = 1e-8
+ wmax = 1.2e-6
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 4.148964422023837e-25
+ wmin = 5e-7
+ nqsmod = 0
+ tpbswg = 0.001554306
+ noimod = 2
+ lmax = 2.0001e-5
+ wketa = 2.1944087e-10
+ pvth0 = 2.71152e-15
+ lmin = 1e-5
+ drout = 0.0
+ tpbsw = 0.001554306
+ )

.model nch_sf_10 nmos (
+ level = 49
+ lute = -1.2190513e-8
+ nqsmod = 0
+ tpbswg = 0.001554306
+ noimod = 2
+ cdsc = 0.0
+ cgdo = 3.665e-10
+ nfactor = 1.0
+ lketa = -2.8027248e-8
+ cgso = 3.665e-10
+ xpart = 1
+ cjsw = 2.142574e-10
+ pbswg = 0.6882682
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0003968185
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ pdiblcb = 0.01
+ lpscbe1 = 262.58185
+ lvoff = -4.506062e-9
+ capmod = 3
+ beta0 = 11.59263
+ tnom = 25.0
+ leta0 = 9.680916984722288e-19
+ binunit = 2
+ lvsat = -0.006201102
+ toxm = 4.08e-9
+ lvth0 = 6.8541616e-8
+ pcit = 4.302753e-19
+ pbsw = 0.6882682
+ pclm = 0.7699873
+ ppclm = 1.243718e-13
+ mobmod = 1
+ delta = 0.01
+ ags = 0.02
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ cit = -0.00012672294
+ dlc = 3e-9
+ k3b = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ pnfactor = 0.0
+ pkt1 = 7.833639e-15
+ pkt2 = 9.747044e-16
+ keta = 0.00382927
+ wnfactor = 0.0
+ pketa = -6.831802e-16
+ version = 3.24
+ dsub = 0.0
+ wpclm = -1.2487239e-8
+ wcit = -4.317371e-14
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ la0 = -1.9725388e-7
+ tcjsw = 0.000645489
+ jsw = 1.45e-12
+ tcjswg = 0.000645489
+ lk1 = 1.0512358e-8
+ kt1 = -0.2310088
+ lk2 = -1.7946909999999996e-9
+ kt2 = -0.028688708
+ lcit = 2.6616018e-10
+ llc = -0.039
+ lln = -1
+ voff = -0.14154522
+ lu0 = 3.253832e-9
+ lnfactor = 4.5192e-8
+ ldif = 9e-8
+ lua = -1.9124487e-16
+ lub = 4.117038e-25
+ luc = 4.038815e-17
+ nch = 3.9e+17
+ pvoff = -6.159972e-15
+ lwl = 0.0
+ lwn = 1.0
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ pub1 = -1.8996434e-32
+ puc1 = 1.3569954e-23
+ pa0 = -1.0015934e-13
+ nlx = 0.0
+ eta0 = 5e-5
+ pk1 = -1.457495e-14
+ pk2 = 2.2122807e-15
+ pvag = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ etab = -5e-5
+ peta0 = 4.148964422023837e-25
+ vsat = 87007.25
+ wint = 3e-9
+ pu0 = 1.6856667e-15
+ pute = -3.577514e-14
+ pvsat = 1.2437262e-9
+ vth0 = 0.45254382
+ prt = 0
+ pua = 4.758471e-23
+ pub = -5.695533e-32
+ puc = -9.239189e-24
+ lpdiblc2 = 3.0196912e-9
+ wketa = 2.8803285e-10
+ rdsw = 170.0
+ pvth0 = -4.446152000000001e-15
+ wkt1 = 6.625341e-10
+ wkt2 = -8.725676e-11
+ drout = 0.0
+ lint = 1e-8
+ rsh = 6.8
+ tpbsw = 0.001554306
+ wmax = 1.2e-6
+ tcj = 0.001040287
+ ua1 = 1.224e-9
+ ub1 = -1.5338095e-18
+ uc1 = -7.316409e-11
+ wmin = 5e-7
+ lkt1 = -3.0828107e-9
+ lkt2 = -3.866881e-9
+ tpb = 0.001554306
+ tox = 4.08e-9
+ cjswg = 3.507574e-10
+ lmax = 1e-5
+ wa0 = 8.672666e-8
+ lmin = 1.2e-6
+ ute = -1.6080947
+ mjswg = 0.43879
+ wk1 = -1.9283881e-8
+ wk2 = 4.698517e-9
+ wln = 1.0
+ wu0 = 8.670528e-10
+ wvoff = -9.715325e-10
+ wua = 1.3831368e-16
+ wub = -1.4839938e-25
+ wuc = -1.3213606e-17
+ wwl = 0.0
+ wwn = 1
+ xti = 3
+ a0 = 0.324591
+ a1 = 0.0
+ a2 = 0.99
+ b0 = 0.0
+ b1 = 0.0
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ wub1 = -5.768295e-27
+ wuc1 = -1.6068998e-17
+ weta0 = 0
+ at = 20000.0
+ cf = 0
+ cj = 0.001050279
+ ef = 0.874
+ k1 = 0.5600169
+ k2 = 0.008916168700000001
+ k3 = 0.0
+ em = 30000000.0
+ hdif = 2e-7
+ wvsat = -0.00012487893
+ js = 3.5e-7
+ pscbe1 = 173636400.0
+ pscbe2 = 1e-6
+ ll = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ u0 = 0.033019980000000004
+ pb = 0.6882682
+ lub1 = 3.243357e-25
+ lpclm = 2.9892766e-7
+ wvth0 = 2.4208780000000006e-9
+ luc1 = 4.341489e-17
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ wute = 4.195195e-8
+ ua = -8.874397e-10
+ ub = 2.2584638e-18
+ uc = 1.0315766e-10
+ mjsw = 0.2003879
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ )

.model nch_sf_11 nmos (
+ level = 49
+ lvoff = 1.025939e-8
+ wcit = 5.431231e-13
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ ags = 0.02
+ beta0 = 11.59263
+ leta0 = 3.8114300968091695e-11
+ lcit = 3.0283653e-10
+ cit = -0.0001583405
+ letab = -3.81143e-11
+ voff = -0.15427401999999998
+ ldif = 9e-8
+ lvsat = -0.0007659488
+ dlc = 3e-9
+ kt1l = 0.0
+ mobmod = 1
+ prwb = 0.0
+ lvth0 = 1.2730886999999999e-8
+ prwg = 0.0
+ pub1 = -5.874811e-31
+ puc1 = -3.67348e-23
+ a0 = -0.1914371
+ a1 = 0.0
+ a2 = 0.99
+ k3b = 0.0
+ b0 = 0.0
+ b1 = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ eta0 = 1.7142847e-5
+ at = 20000.0
+ cf = 0
+ cj = 0.001050279
+ ef = 0.874
+ k1 = 0.5552615
+ ppclm = 7.308824e-14
+ k2 = 0.010775519
+ k3 = 0.0
+ em = 30000000.0
+ pvag = 0.0
+ etab = -1.7142847e-5
+ delta = 0.01
+ js = 3.5e-7
+ vsat = 82321.77
+ ll = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ u0 = 0.03400418
+ pb = 0.6882682
+ wint = 3e-9
+ pute = -2.0303331e-13
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ua = -1.3333591e-9
+ ub = 2.969086e-18
+ uc = 1.6160392e-10
+ vth0 = 0.50065652
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ rdsw = 170.0
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ wkt1 = 1.1898274e-8
+ wkt2 = 2.0987987e-9
+ lint = 1e-8
+ wmax = 1.2e-6
+ la0 = 4.013388e-7
+ wmin = 5e-7
+ lkt1 = 9.329063e-9
+ lkt2 = 2.691467e-9
+ jsw = 1.45e-12
+ lk1 = 1.6028618e-8
+ kt1 = -0.2417087
+ lk2 = -3.9515360000000006e-9
+ kt2 = -0.03434246
+ lmax = 1.2e-6
+ llc = -0.039
+ lln = -1
+ lu0 = 2.1121620999999997e-9
+ lmin = 5e-7
+ lua = 3.260216e-16
+ lub = -4.12618e-25
+ luc = -2.7409531e-17
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ pketa = 1.4501565e-15
+ pa0 = 1.1848049e-14
+ nlx = 0.0
+ pk1 = 7.144098e-15
+ pk2 = -4.137203e-15
+ pu0 = -1.1138246e-15
+ wpclm = 3.172275e-8
+ wub1 = 4.843047e-25
+ prt = 0
+ wuc1 = 2.7297169e-17
+ pua = -1.3255767e-22
+ pub = 5.546348e-32
+ puc = -6.669366e-24
+ tcjswg = 0.000645489
+ hdif = 2e-7
+ tcjsw = 0.000645489
+ rsh = 6.8
+ lub1 = 4.951269e-25
+ luc1 = 6.070172e-17
+ tcj = 0.001040287
+ ua1 = 1.224e-9
+ ub1 = -1.6810433e-18
+ uc1 = -8.806652e-11
+ wute = 1.8614003e-7
+ mjsw = 0.2003879
+ pvoff = 1.9014135e-15
+ tpb = 0.001554306
+ tox = 4.08e-9
+ wa0 = -9.831444e-9
+ lute = 2.2508574e-7
+ ute = -1.8126432
+ wk1 = -3.80072e-8
+ wk2 = 1.0172209e-8
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 4.148964422023837e-25
+ wln = 1.0
+ wu0 = 3.280407e-9
+ wua = 2.9360883e-16
+ pvsat = 4.380818e-12
+ wub = -2.4531215e-25
+ wuc = -1.542897e-17
+ wwl = 0.0
+ wwn = 1
+ cdsc = 0.0
+ wketa = -1.5510503e-9
+ pvth0 = 2.1736318e-15
+ xti = 3
+ drout = 0.0
+ cgdo = 3.665e-10
+ tpbsw = 0.001554306
+ cgso = 3.665e-10
+ cjswg = 3.507574e-10
+ nfactor = 1.0
+ mjswg = 0.43879
+ pnfactor = 0.0
+ cjsw = 2.142574e-10
+ wnfactor = 0.0
+ wvoff = -7.921003e-9
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ weta0 = 0
+ pscbe1 = 400000100.0
+ pscbe2 = 1e-6
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0011219129
+ pdiblcb = 0.01
+ wvsat = 0.0009435224
+ ppdiblc2 = 1.2928064e-16
+ tnom = 25.0
+ lpclm = 9.659676e-8
+ wvth0 = -3.2858339999999996e-9
+ wpdiblc2 = -1.1144895e-10
+ lnfactor = 4.5192e-8
+ nqsmod = 0
+ tpbswg = 0.001554306
+ toxm = 4.08e-9
+ noimod = 2
+ pcit = -2.4980728e-19
+ binunit = 2
+ pbsw = 0.6882682
+ pclm = 0.9444105
+ lpdiblc2 = 2.1785818e-9
+ lketa = -2.9090079e-9
+ xpart = 1
+ pkt1 = -5.199821e-15
+ pkt2 = -1.5611203e-15
+ keta = -0.017824383
+ pbswg = 0.6882682
+ dsub = 0.0
+ capmod = 3
+ version = 3.24
+ )

.model nch_sf_12 nmos (
+ level = 49
+ tpb = 0.001554306
+ tox = 4.08e-9
+ wa0 = 1.7605426e-7
+ pketa = -7.367843e-16
+ cjsw = 2.142574e-10
+ nfactor = 1.0
+ ute = -1.2073984
+ wk1 = -1.7855582e-8
+ wk2 = 1.6966123e-9
+ tcjswg = 0.000645489
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ wln = 1.0
+ wu0 = -4.268465e-11
+ wpclm = 1.9327061e-7
+ wua = -1.9101984e-17
+ wub = -5.11281e-26
+ wuc = -9.012729e-18
+ wwl = 0.0
+ wwn = 1
+ xti = 3
+ tcjsw = 0.000645489
+ tnom = 25.0
+ pdiblc1 = 1e-6
+ pdiblc2 = -0.00401322
+ pags = 1.8981756e-15
+ pdiblcb = 0.01
+ pvoff = -3.1245874000000002e-15
+ toxm = 4.08e-9
+ pcit = -1.4232223e-17
+ pbsw = 0.6882682
+ pclm = 0.9948969
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = -1.1371990585103558e-17
+ petab = 1.3954016e-17
+ binunit = 2
+ pvsat = 1.606088e-11
+ wketa = 3.203169e-9
+ pvth0 = 5.427536e-15
+ drout = 0.0
+ tpbsw = 0.001554306
+ a0 = 0.5005398
+ a1 = 0.0
+ a2 = 0.99
+ b0 = 0.0
+ b1 = 0.0
+ at = 20000.0
+ cf = 0
+ cj = 0.001050279
+ ef = 0.874
+ k1 = 0.489967
+ k2 = 0.036529204
+ k3 = 0.0
+ em = 30000000.0
+ js = 3.5e-7
+ cjswg = 3.507574e-10
+ ll = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ u0 = 0.03799784
+ pb = 0.6882682
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ua = -5.274002e-10
+ ub = 2.0039751e-18
+ uc = 7.914647e-11
+ mjswg = 0.43879
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ pkt1 = 2.3961372e-15
+ pkt2 = 8.832021e-16
+ keta = -0.027587207
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ wvoff = 3.005086e-9
+ wags = -4.12647e-9
+ dsub = 0.0
+ pscbe1 = 400000000.0
+ pscbe2 = 1e-6
+ weta0 = 2.4721704e-11
+ lags = -9.594464e-9
+ wetab = -3.0334849e-11
+ wcit = 3.093965e-11
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ wvsat = 0.000918131
+ version = 3.24
+ nqsmod = 0
+ lpclm = 7.337301e-8
+ wvth0 = -1.0359539e-8
+ tpbswg = 0.001554306
+ noimod = 2
+ lcit = 1.2733804e-10
+ voff = -0.12912402
+ ldif = 9e-8
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ pub1 = 1.6165291e-31
+ puc1 = 2.0250814e-23
+ eta0 = -0.00031223928
+ pvag = 0.0
+ etab = 0.0014101875
+ vsat = 81120.94
+ wint = 3e-9
+ pute = 4.383575e-14
+ vth0 = 0.50768662
+ rdsw = 170.0
+ wkt1 = -4.614678e-9
+ wkt2 = -3.214946e-9
+ lint = 1e-8
+ wmax = 1.2e-6
+ ags = 0.04085753
+ lketa = 1.5818911e-9
+ wmin = 5e-7
+ lkt1 = 1.6202869e-9
+ lkt2 = -8.228257e-11
+ lmax = 5e-7
+ xpart = 1
+ cit = 0.00022317801
+ lmin = 1.8e-7
+ pnfactor = 0.0
+ dlc = 3e-9
+ wnfactor = 0.0
+ k3b = 0.0
+ capmod = 3
+ dwb = 0.0
+ dwg = 0.0
+ pbswg = 0.6882682
+ lvoff = -1.3096095e-9
+ wub1 = -1.1442477e-24
+ wuc1 = -9.658459e-17
+ ppdiblc2 = 3.905237e-16
+ hdif = 2e-7
+ beta0 = 11.59263
+ wpdiblc2 = -6.793707e-10
+ lub1 = -6.558089e-26
+ leta0 = 1.8963006096809171e-10
+ luc1 = -7.416688e-18
+ wute = -3.505318e-7
+ mobmod = 1
+ la0 = 8.302936e-8
+ letab = -6.946862e-10
+ lnfactor = 4.5192e-8
+ mjsw = 0.2003879
+ lvsat = -0.00021356932
+ jsw = 1.45e-12
+ lk1 = 4.606408e-8
+ kt1 = -0.2249505
+ lk2 = -1.5798233e-8
+ kt2 = -0.028312566
+ lvth0 = 9.497081e-9
+ llc = -0.039
+ lln = -1
+ lute = -5.332685e-8
+ lu0 = 2.7507449999999995e-10
+ lua = -4.471944e-17
+ lub = 3.1333025e-26
+ luc = 1.0520902e-17
+ ppclm = -1.2237712e-15
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ delta = 0.01
+ pa0 = -7.365936e-14
+ nlx = 0.0
+ lpdiblc2 = 4.540744e-9
+ cdsc = 0.0
+ pk1 = -2.1256446e-15
+ pk2 = -2.3842633e-16
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ pu0 = 4.147977e-16
+ cgdo = 3.665e-10
+ prt = 0
+ pua = 1.1289303e-23
+ pub = -3.386118e-32
+ puc = -9.620837e-24
+ cgso = 3.665e-10
+ rsh = 6.8
+ tcj = 0.001040287
+ ua1 = 1.224e-9
+ ub1 = -4.621132e-19
+ uc1 = 6.001696e-11
+ )

.model nch_sf_13 nmos (
+ level = 49
+ drout = 0.0
+ wkt1 = 5.128653e-9
+ wkt2 = 3.532295e-9
+ tpbsw = 0.001554306
+ lint = 1e-8
+ wmax = 5e-7
+ wmin = 2.2e-7
+ cjswg = 3.507574e-10
+ lmax = 2.0001e-5
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ mjswg = 0.43879
+ lmin = 1e-5
+ pscbe1 = 200000030.0
+ pscbe2 = 1e-6
+ wvoff = -2.3603662000000002e-9
+ weta0 = 0
+ nqsmod = 0
+ wub1 = -4.432931e-26
+ wuc1 = -1.7086574e-17
+ tpbswg = 0.001554306
+ wvsat = 0.0
+ noimod = 2
+ hdif = 2e-7
+ wvth0 = -9.490401e-9
+ ags = 0.02
+ wute = 2.5547985e-8
+ mjsw = 0.2003879
+ cit = -9.999998e-5
+ dlc = 3e-9
+ k3b = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ cdsc = 0.0
+ cgdo = 3.665e-10
+ cgso = 3.665e-10
+ xpart = 1
+ jsw = 1.45e-12
+ capmod = 3
+ kt1 = -0.238767
+ lk2 = 3.6153600000000002e-9
+ kt2 = -0.03620588
+ llc = -0.039
+ cjsw = 2.142574e-10
+ lln = -1
+ a0 = 0.352982
+ a1 = 0.0
+ a2 = 0.99
+ lu0 = -4.5192000000000003e-10
+ b0 = 0.0
+ b1 = 0.0
+ pbswg = 0.6882682
+ nch = 3.9e+17
+ at = 20000.0
+ cf = 0
+ cj = 0.001050279
+ lwl = 0.0
+ lwn = 1.0
+ ef = 0.874
+ k1 = 0.5220979
+ k2 = 0.023773289
+ k3 = 0.0
+ em = 30000000.0
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ nfactor = 1.0
+ js = 3.5e-7
+ ll = 0.0
+ nlx = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ lvoff = -9.038400000000001e-10
+ u0 = 0.03352974
+ pb = 0.6882682
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ua = -5.860608e-10
+ ub = 1.7266676e-18
+ uc = 7.252202e-11
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ mobmod = 1
+ beta0 = 11.59263
+ pu0 = 0.0
+ tnom = 25.0
+ leta0 = 9.680916984722288e-19
+ prt = 0
+ toxm = 4.08e-9
+ rsh = 6.8
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0006999999
+ lvth0 = 2.621136e-9
+ tcj = 0.001040287
+ ua1 = 1.224e-9
+ ub1 = -1.4270478e-18
+ uc1 = -6.39873e-11
+ pdiblcb = 0.01
+ pbsw = 0.6882682
+ pclm = 0.7999999
+ tpb = 0.001554306
+ tox = 4.08e-9
+ delta = 0.01
+ wa0 = 5.286186e-8
+ ute = -1.5833832
+ wk1 = -1.4938487e-9
+ wk2 = -2.6871128e-9
+ dvt0w = 0.0
+ dvt1w = 0.0
+ wln = 1.0
+ dvt2w = 0.0
+ wu0 = 9.682726e-10
+ binunit = 2
+ wua = -1.5275344e-17
+ wub = 1.2900942e-25
+ wuc = 2.9959555e-18
+ wwl = 0.0
+ wwn = 1
+ xti = 3
+ pnfactor = 0.0
+ keta = 0.002064252
+ tcjswg = 0.000645489
+ wnfactor = 0.0
+ dsub = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ tcjsw = 0.000645489
+ lnfactor = 4.5192e-8
+ voff = -0.14016372
+ version = 3.24
+ pvoff = -9.038400000000001e-16
+ ldif = 9e-8
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ eta0 = 5e-5
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 4.148964422023837e-25
+ pvag = 0.0
+ etab = -5e-5
+ vsat = 86384.63
+ wint = 3e-9
+ vth0 = 0.48181952
+ wketa = -2.9874625e-10
+ pvth0 = 2.71152e-15
+ rdsw = 170.0
+ )

.model nch_sf_14 nmos (
+ level = 49
+ la0 = -2.4964379e-7
+ pcit = 1.5653096e-18
+ pbsw = 0.6882682
+ pclm = 0.7606163
+ jsw = 1.45e-12
+ lk1 = -6.331243e-8
+ kt1 = -0.2407974
+ lk2 = 2.4414092e-8
+ kt2 = -0.03589625
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0003968183
+ pdiblcb = 0.01
+ lpscbe1 = 262.58182
+ llc = -0.039
+ lln = -1
+ lu0 = 9.442635e-9
+ lpdiblc2 = 3.0196909e-9
+ lua = -1.2876533e-16
+ lub = 7.836163e-25
+ luc = 7.064626e-17
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ pa0 = -7.427873e-14
+ nlx = 0.0
+ pk1 = 2.1894499e-14
+ pk2 = -1.0734859e-14
+ lketa = -3.0377027e-8
+ binunit = 2
+ pu0 = -1.3716021e-15
+ capmod = 3
+ prt = 0
+ pua = 1.6719826e-23
+ pub = -2.4068014e-31
+ xpart = 1
+ puc = -2.4186704e-23
+ pkt1 = -3.679308e-15
+ pkt2 = 5.879336e-16
+ rsh = 6.8
+ keta = 0.005114151
+ tcj = 0.001040287
+ ua1 = 1.224e-9
+ ub1 = -1.4513121e-18
+ uc1 = -6.991786e-11
+ pbswg = 0.6882682
+ tpb = 0.001554306
+ tox = 4.08e-9
+ dsub = 0.0
+ wa0 = 6.031956e-8
+ lvoff = -2.0631212000000003e-8
+ mobmod = 1
+ ute = -1.5785241
+ wk1 = -3.692092e-9
+ wk2 = -1.6093152e-9
+ wcit = -1.5715551e-13
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ wln = 1.0
+ beta0 = 11.59263
+ wu0 = 1.1059835e-9
+ wua = -1.6954039e-17
+ wub = 1.5317406e-25
+ wuc = 5.42434e-18
+ leta0 = 9.680916984722288e-19
+ wwl = 0.0
+ wwn = 1
+ lcit = 2.6386249e-10
+ xti = 3
+ voff = -0.13818312
+ lvsat = -0.005267757
+ ldif = 9e-8
+ lvth0 = 5.8899376e-8
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ pub1 = 2.1839324e-32
+ puc1 = 5.837128e-24
+ version = 3.24
+ ppclm = 7.826515e-14
+ eta0 = 5e-5
+ delta = 0.01
+ pvag = 0.0
+ etab = -5e-5
+ vsat = 86913.52
+ wint = 3e-9
+ pute = -1.7889165e-14
+ vth0 = 0.47616912
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ rdsw = 170.0
+ wkt1 = 5.498062e-9
+ wkt2 = 3.473265e-9
+ lint = 1e-8
+ wmax = 5e-7
+ wmin = 2.2e-7
+ lkt1 = 2.0222748e-8
+ lkt2 = -3.0839447e-9
+ lmax = 1e-5
+ tcjswg = 0.000645489
+ lmin = 1.2e-6
+ pketa = 4.776125e-16
+ wpclm = -7.857923e-9
+ wub1 = -4.652201e-26
+ wuc1 = -1.7672629e-17
+ tcjsw = 0.000645489
+ hdif = 2e-7
+ lub1 = 2.4167225e-25
+ a0 = 0.3780467
+ a1 = 0.0
+ a2 = 0.99
+ luc1 = 5.906839e-17
+ b0 = 0.0
+ b1 = 0.0
+ wute = 2.7344081e-8
+ mjsw = 0.2003879
+ at = 20000.0
+ pvoff = 1.8058529e-15
+ cf = 0
+ cj = 0.001050279
+ ef = 0.874
+ k1 = 0.5284545
+ k2 = 0.021685062
+ k3 = 0.0
+ em = 30000000.0
+ js = 3.5e-7
+ ll = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ u0 = 0.03253632
+ pb = 0.6882682
+ w0 = 0.0
+ rd = 0
+ lute = -4.839696e-8
+ rs = 0
+ ua = -5.731325e-10
+ ub = 1.6479914e-18
+ uc = 6.542903e-11
+ cdscb = 0.0
+ cdscd = 0.0
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -2e-8
+ ww = 0.0
+ peta0 = 4.148964422023837e-25
+ xw = 0.0
+ pvsat = 7.826533e-10
+ wketa = -3.466991e-10
+ pvth0 = 3.1711749999999997e-16
+ cdsc = 0.0
+ drout = 0.0
+ tpbsw = 0.001554306
+ cgdo = 3.665e-10
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ cgso = 3.665e-10
+ cjswg = 3.507574e-10
+ pscbe1 = 173636400.0
+ pscbe2 = 1e-6
+ mjswg = 0.43879
+ ags = 0.02
+ pnfactor = 0.0
+ wnfactor = 0.0
+ wvoff = -2.6324233e-9
+ cjsw = 2.142574e-10
+ cit = -0.00012649217
+ nqsmod = 0
+ dlc = 3e-9
+ tpbswg = 0.001554306
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ noimod = 2
+ k3b = 0.0
+ weta0 = 0
+ dwb = 0.0
+ dwg = 0.0
+ wvsat = -7.857954e-5
+ nfactor = 1.0
+ lpclm = 3.92261e-7
+ wvth0 = -9.25e-9
+ tnom = 25.0
+ lnfactor = 4.5192e-8
+ toxm = 4.08e-9
+ )

.model nch_sf_15 nmos (
+ level = 49
+ wub1 = -1.0574451e-25
+ wuc1 = -4.040928e-17
+ ppdiblc2 = 4.703685e-16
+ beta0 = 11.59263
+ hdif = 2e-7
+ wpdiblc2 = -4.054901e-10
+ leta0 = 3.8114280968091696e-11
+ lub1 = -8.773805e-25
+ luc1 = -7.886598e-17
+ letab = -3.811428e-11
+ lnfactor = 4.5192e-8
+ wute = 1.9757099e-8
+ lvsat = -0.0007893788
+ mjsw = 0.2003879
+ lvth0 = 1.1480395e-8
+ lute = -1.6751561e-7
+ ppclm = 4.863229e-14
+ delta = 0.01
+ lpdiblc2 = 1.4881204e-9
+ dvt0w = 0.0
+ cdsc = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ cgdo = 3.665e-10
+ tcjswg = 0.000645489
+ cgso = 3.665e-10
+ pketa = 3.1429577e-15
+ cjsw = 2.142574e-10
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ wpclm = 1.7687656e-8
+ tcjsw = 0.000645489
+ tnom = 25.0
+ nfactor = 1.0
+ pvoff = -2.2875942e-15
+ toxm = 4.08e-9
+ ags = 0.02
+ pcit = -9.088336e-19
+ pbsw = 0.6882682
+ pclm = 0.9728217
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 4.148964422023837e-25
+ pvsat = 1.5955267e-11
+ cit = -0.00016124053
+ wketa = -2.6444102e-9
+ pvth0 = 2.7913746499999998e-15
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0017171376
+ dlc = 3e-9
+ drout = 0.0
+ pdiblcb = 0.01
+ k3b = 0.0
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ tpbsw = 0.001554306
+ dwb = 0.0
+ dwg = 0.0
+ pscbe1 = 400000100.0
+ pscbe2 = 1e-6
+ cjswg = 3.507574e-10
+ mjswg = 0.43879
+ binunit = 2
+ pkt1 = -1.1651986e-14
+ pkt2 = -1.4582807e-15
+ keta = -0.015611105
+ nqsmod = 0
+ wvoff = 8.9641e-10
+ tpbswg = 0.001554306
+ la0 = 2.7901473e-7
+ noimod = 2
+ jsw = 1.45e-12
+ dsub = 0.0
+ lk1 = 6.936774e-8
+ kt1 = -0.2426658
+ lk2 = -2.7913247000000003e-8
+ kt2 = -0.04069558
+ llc = -0.039
+ lln = -1
+ weta0 = 0
+ lu0 = -2.1965306e-9
+ lua = 6.135559e-17
+ lub = -2.9489129e-25
+ luc = -2.7169401e-17
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ wvsat = 0.0005823669
+ wcit = 1.975718e-12
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ pa0 = 7.227613e-14
+ nlx = 0.0
+ lpclm = 1.4610272e-7
+ wvth0 = -1.138298e-8
+ pk1 = -1.920543e-14
+ pk2 = 7.699883e-15
+ lcit = 3.0417063e-10
+ voff = -0.17212312
+ pu0 = 1.0146696e-15
+ ldif = 9e-8
+ prt = 0
+ pua = -1.8126578e-24
+ pub = -2.6935e-33
+ puc = -6.78799e-24
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ pub1 = 9.053745e-32
+ puc1 = 3.221165e-23
+ eta0 = 1.7142866e-5
+ rsh = 6.8
+ pvag = 0.0
+ etab = -1.7142866e-5
+ tcj = 0.001040287
+ ua1 = 1.224e-9
+ ub1 = -4.866116e-19
+ uc1 = 4.899104e-11
+ vsat = 83052.85
+ version = 3.24
+ a0 = -0.07769345
+ wint = 3e-9
+ a1 = 0.0
+ a2 = 0.99
+ pute = -9.088265e-15
+ b0 = 0.0
+ b1 = 0.0
+ tpb = 0.001554306
+ vth0 = 0.51704752
+ tox = 4.08e-9
+ at = 20000.0
+ cf = 0
+ cj = 0.001050279
+ ef = 0.874
+ k1 = 0.4140751
+ k2 = 0.06679484
+ k3 = 0.0
+ rdsw = 170.0
+ wa0 = -6.602082e-8
+ em = 30000000.0
+ js = 3.5e-7
+ wkt1 = 1.2371058e-8
+ wkt2 = 5.237243e-9
+ ute = -1.4758356
+ ll = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ lint = 1e-8
+ u0 = 0.04257008
+ pb = 0.6882682
+ wk1 = 3.173889e-8
+ wk2 = -1.7501334e-8
+ w0 = 0.0
+ rd = 0
+ wmax = 5e-7
+ lketa = -6.33573e-9
+ capmod = 3
+ rs = 0
+ ua = -7.370299e-10
+ ub = 2.5777392e-18
+ uc = 1.4975288e-10
+ wln = 1.0
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -2e-8
+ ww = 0.0
+ wmin = 2.2e-7
+ wu0 = -9.511471e-10
+ xw = 0.0
+ lkt1 = 2.2390124e-8
+ wua = -9.777621e-19
+ lkt2 = 2.4832894e-9
+ wub = -5.19868e-26
+ wuc = -9.57455e-18
+ xpart = 1
+ wwl = 0.0
+ wwn = 1
+ lmax = 1.2e-6
+ xti = 3
+ lmin = 5e-7
+ pnfactor = 0.0
+ wnfactor = 0.0
+ pbswg = 0.6882682
+ mobmod = 1
+ lvoff = 1.8739164e-8
+ )

.model nch_sf_16 nmos (
+ level = 49
+ at = 20000.0
+ cf = 0
+ cj = 0.001050279
+ ef = 0.874
+ k1 = 0.4942783
+ k2 = 0.030748973
+ k3 = 0.0
+ em = 30000000.0
+ pketa = -1.9609824e-16
+ pkt1 = 3.435378e-15
+ pkt2 = -8.505888e-17
+ wnfactor = 0.0
+ keta = -0.030443965
+ js = 3.5e-7
+ ll = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ ags = 0.0548038
+ u0 = 0.03529582
+ pb = 0.6882682
+ w0 = 0.0
+ binunit = 2
+ rd = 0
+ rs = 0
+ ua = -6.614348e-10
+ ub = 2.1301375e-18
+ uc = 1.2526492e-10
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ wags = -1.1015922e-8
+ xl = -2e-8
+ ww = 0.0
+ dsub = 0.0
+ xw = 0.0
+ wpclm = 1.2379924e-7
+ cit = 0.00029138371
+ lags = -1.6009743e-8
+ dlc = 3e-9
+ wcit = -2.7539906e-12
+ ppdiblc2 = -1.1422951e-16
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ tcjsw = 0.000645489
+ k3b = 0.0
+ wpdiblc2 = 8.65375e-10
+ dwb = 0.0
+ dwg = 0.0
+ lnfactor = 4.5192e-8
+ lcit = 9.596344e-11
+ pvoff = -1.4007737000000002e-15
+ voff = -0.12095291999999999
+ ldif = 9e-8
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ pub1 = -3.181536e-32
+ puc1 = -1.1609298e-23
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 4.148964422023837e-25
+ eta0 = -0.00026219533
+ pvag = 0.0
+ etab = 0.0013487812
+ pvsat = 1.2452966e-11
+ la0 = 1.1871046e-7
+ vsat = 81785.22
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ wint = 3e-9
+ pute = -6.731688e-15
+ wketa = 4.614407e-9
+ lpdiblc2 = 5.562512e-9
+ pvth0 = 1.6693625999999999e-15
+ jsw = 1.45e-12
+ vth0 = 0.50482072
+ lk1 = 3.247429e-8
+ kt1 = -0.1929406
+ lk2 = -1.1332151999999999e-8
+ kt2 = -0.03937921
+ drout = 0.0
+ rdsw = 170.0
+ llc = -0.039
+ lln = -1
+ tpbsw = 0.001554306
+ pscbe1 = 400000000.0
+ pscbe2 = 1e-6
+ lu0 = 1.1496252e-9
+ version = 3.24
+ wkt1 = -2.0427562e-8
+ wkt2 = 2.2519782e-9
+ lint = 1e-8
+ lua = 2.6581833e-17
+ lub = -8.899446e-26
+ luc = -1.5904941e-17
+ nch = 3.9e+17
+ wmax = 5e-7
+ lwl = 0.0
+ lwn = 1.0
+ wmin = 2.2e-7
+ pa0 = -9.128582e-14
+ nlx = 0.0
+ cjswg = 3.507574e-10
+ lkt1 = -4.834396e-10
+ lkt2 = 1.8777602e-9
+ mjswg = 0.43879
+ pk1 = 4.587708e-15
+ pk2 = -2.4446703e-15
+ lmax = 5e-7
+ nqsmod = 0
+ tpbswg = 0.001554306
+ lmin = 1.8e-7
+ noimod = 2
+ pu0 = -1.7230291e-17
+ prt = 0
+ pua = -2.3933522e-23
+ pub = 2.5580594e-32
+ puc = 3.433529e-24
+ wvoff = -1.031461e-9
+ rsh = 6.8
+ tcj = 0.001040287
+ ua1 = 1.224e-9
+ ub1 = -3.1027764e-18
+ uc1 = -2.4653823e-10
+ weta0 = 0
+ tpb = 0.001554306
+ wub1 = 1.602399e-25
+ wuc1 = 5.485366e-17
+ tox = 4.08e-9
+ wvsat = 0.0005899806
+ wa0 = 2.8954867e-7
+ hdif = 2e-7
+ lpclm = 7.125815e-8
+ wvth0 = -8.94382e-9
+ ute = -1.9466008
+ wk1 = -1.9985334e-8
+ wk2 = 4.552045e-9
+ lub1 = 3.260553e-25
+ luc1 = 5.707747e-17
+ wute = 1.4634106e-8
+ wln = 1.0
+ mjsw = 0.2003879
+ wu0 = 1.2921135e-9
+ wua = 4.711108e-17
+ wub = -1.1345223e-25
+ wuc = -3.179524e-17
+ wwl = 0.0
+ wwn = 1
+ xti = 3
+ lute = 4.90364e-8
+ cdsc = 0.0
+ capmod = 3
+ cgdo = 3.665e-10
+ lketa = 4.87385e-10
+ cgso = 3.665e-10
+ xpart = 1
+ mobmod = 1
+ cjsw = 2.142574e-10
+ pbswg = 0.6882682
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ lvoff = -4.7991109999999995e-9
+ beta0 = 11.59263
+ leta0 = 1.666098409680917e-10
+ tnom = 25.0
+ letab = -6.664392e-10
+ lvsat = -0.00020626588
+ pags = 5.067323e-15
+ lvth0 = 1.7104719e-8
+ toxm = 4.08e-9
+ nfactor = 1.0
+ pcit = 1.266836e-18
+ ppclm = -1.7902992e-16
+ pbsw = 0.6882682
+ pclm = 1.1355271
+ delta = 0.01
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ tcjswg = 0.000645489
+ pdiblc1 = 1e-6
+ pdiblc2 = -0.007140237
+ pdiblcb = 0.01
+ a0 = 0.270794
+ a1 = 0.0
+ a2 = 0.99
+ b0 = 0.0
+ b1 = 0.0
+ pnfactor = 0.0
+ )

.model nch_mc_1 nmos (
+ level = 49
+ cjsw = 2.040547e-10
+ drout = 0.0
+ tpbsw = 0.001554306
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ cjswg = 3.340547e-10
+ pnfactor = 0.0
+ mjswg = 0.43879
+ wnfactor = 0.0
+ tnom = 25.0
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ wvoff = 0.0
+ pscbe1 = 200000030.0
+ pscbe2 = 1e-6
+ toxm = 4.08e-9
+ version = 3.24
+ pbsw = 0.6882682
+ pclm = 0.8000001
+ weta0 = 0
+ wvsat = 0.0
+ nqsmod = 0
+ lnfactor = 0.0
+ tpbswg = 0.001554306
+ wvth0 = 0.0
+ noimod = 2
+ ags = 0.02
+ keta = 0.009263485
+ cit = -0.00010000001
+ a0 = 0.3700794
+ a1 = 0.0
+ a2 = 0.99
+ b0 = 0.0
+ b1 = 0.0
+ dlc = 3e-9
+ dsub = 0.0
+ k3b = 0.0
+ at = 20000.0
+ cf = 0
+ cj = 0.001000266
+ ef = 0.874
+ k1 = 0.5142301
+ k2 = 0.014797844
+ k3 = 0.0
+ em = 30000000.0
+ dwb = 0.0
+ dwg = 0.0
+ js = 3.5e-7
+ ll = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ u0 = 0.04220339
+ pb = 0.6882682
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ dvt0 = 0.0
+ ua = -6.12274e-10
+ dvt1 = 0.0
+ ub = 2.3135539e-18
+ xpart = 1
+ dvt2 = 0.0
+ uc = 1.0876087e-10
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ voff = -0.140578
+ capmod = 3
+ ldif = 9e-8
+ pbswg = 0.6882682
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ jsw = 1.45e-12
+ kt1 = -0.2240464
+ lk2 = 0.0
+ kt2 = -0.030266136
+ lvoff = 0.0
+ eta0 = 5e-5
+ llc = -0.039
+ lln = -1
+ pvag = 0.0
+ etab = -5e-5
+ lu0 = 0.0
+ vsat = 90000.01
+ beta0 = 11.59263
+ nch = 3.9e+17
+ wint = 3e-9
+ lwl = 0.0
+ lwn = 1.0
+ vth0 = 0.4365561
+ leta0 = 8e-15
+ mobmod = 1
+ nlx = 0.0
+ rdsw = 170.0
+ lint = 1e-8
+ wmax = 0.000900001
+ lvth0 = 0.0
+ pu0 = 0.0
+ wmin = 1e-5
+ prt = 0
+ lmax = 2.0001e-5
+ delta = 0.01
+ lmin = 1e-5
+ rsh = 6.8
+ tcj = 0.001040287
+ ua1 = 1.224e-9
+ ub1 = -1.1209314e-18
+ uc1 = 1.1643822e-11
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ tpb = 0.001554306
+ tox = 4.08e-9
+ ute = -1.5799998
+ wln = 1.0
+ wu0 = 0.0
+ nfactor = 1.0
+ hdif = 2e-7
+ wwl = 0.0
+ wwn = 1
+ xti = 3
+ mjsw = 0.2003879
+ tcjswg = 0.000645489
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0006999999
+ pdiblcb = 0.01
+ tcjsw = 0.000645489
+ cdsc = 0.0
+ pvoff = 0.0
+ cgdo = 3.665e-10
+ binunit = 2
+ cgso = 3.665e-10
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 1.0000000000000001e-20
+ pvth0 = 0.0
+ )

.model nch_mc_2 nmos (
+ level = 49
+ wmax = 0.000900001
+ wmin = 1e-5
+ lkt2 = -4.553491e-12
+ lmax = 1e-5
+ lmin = 1.2e-6
+ la0 = -3.496093e-7
+ jsw = 1.45e-12
+ kt1 = -0.2240468
+ lk1 = 1.4908844e-8
+ kt2 = -0.03026568
+ lk2 = -1.111338e-8
+ llc = -0.039
+ lln = -1
+ lketa = -4.320781e-8
+ lu0 = 3.291809e-9
+ lua = -4.643216e-16
+ lub = 7.375677e-25
+ luc = 3.898355e-17
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ xpart = 1
+ pnfactor = 0.0
+ nlx = 0.0
+ hdif = 2e-7
+ wnfactor = 0.0
+ capmod = 3
+ lub1 = 4.527317e-28
+ luc1 = 7.827772e-20
+ nfactor = 1.0
+ pu0 = 0.0
+ mjsw = 0.2003879
+ prt = 0
+ pbswg = 0.6882682
+ lute = -5.743953e-11
+ lvoff = -1.0471328e-8
+ rsh = 6.8
+ tcj = 0.001040287
+ ua1 = 1.224e-9
+ ub1 = -1.1209769e-18
+ uc1 = 1.1635963e-11
+ mobmod = 1
+ beta0 = 11.59263
+ tpb = 0.001554306
+ tox = 4.08e-9
+ lnfactor = 0.0
+ leta0 = 8e-15
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0003968181
+ cdsc = 0.0
+ pdiblcb = 0.01
+ lpscbe1 = 262.58185
+ ute = -1.5799941
+ lvsat = -0.006562638
+ cgdo = 3.665e-10
+ wln = 1.0
+ lvth0 = 6.061287e-8
+ wu0 = 0.0
+ wwl = 0.0
+ wwn = 1
+ cgso = 3.665e-10
+ xti = 3
+ delta = 0.01
+ lpdiblc2 = 3.0196912e-9
+ binunit = 2
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ cjsw = 2.040547e-10
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ tnom = 25.0
+ tcjswg = 0.000645489
+ a0 = 0.4051808
+ a1 = 0.0
+ a2 = 0.99
+ b0 = 0.0
+ b1 = 0.0
+ at = 20000.0
+ cf = 0
+ cj = 0.001000266
+ ef = 0.874
+ k1 = 0.5127332
+ k2 = 0.015913647
+ k3 = 0.0
+ em = 30000000.0
+ toxm = 4.08e-9
+ js = 3.5e-7
+ ll = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ u0 = 0.04187289
+ pb = 0.6882682
+ w0 = 0.0
+ pbsw = 0.6882682
+ rd = 0
+ pclm = 0.7736172
+ rs = 0
+ ua = -5.656554e-10
+ ub = 2.2395009e-18
+ uc = 1.0484686e-10
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ tcjsw = 0.000645489
+ version = 3.24
+ pvoff = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 1.0000000000000001e-20
+ pvth0 = 0.0
+ keta = 0.013601619
+ drout = 0.0
+ tpbsw = 0.001554306
+ dsub = 0.0
+ cjswg = 3.340547e-10
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ mjswg = 0.43879
+ pscbe1 = 173636400.0
+ pscbe2 = 1e-6
+ lcit = 2.6652053e-10
+ wvoff = 0.0
+ voff = -0.1395267
+ ldif = 9e-8
+ ags = 0.02
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ weta0 = 0
+ nqsmod = 0
+ eta0 = 5e-5
+ tpbswg = 0.001554306
+ pvag = 0.0
+ etab = -5e-5
+ cit = -0.00012675911
+ noimod = 2
+ wvsat = 0.0
+ vsat = 90658.91
+ wint = 3e-9
+ dlc = 3e-9
+ lpclm = 2.6277317e-7
+ wvth0 = 0.0
+ vth0 = 0.4304705
+ k3b = 0.0
+ rdsw = 170.0
+ dwb = 0.0
+ dwg = 0.0
+ lint = 1e-8
+ )

.model nch_mc_3 nmos (
+ level = 49
+ beta0 = 11.59263
+ leta0 = 3.812228e-11
+ letab = -3.811428e-11
+ lvsat = -0.0007622857
+ version = 3.24
+ lvth0 = 3.942757e-9
+ delta = 0.01
+ keta = -0.015927497
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ dsub = 0.0
+ pnfactor = 0.0
+ lags = -3.044698e-8
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ tcjswg = 0.000645489
+ wnfactor = 0.0
+ lcit = 3.0262734e-10
+ voff = -0.1621186
+ ldif = 9e-8
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ eta0 = 1.7142866e-5
+ pvag = 0.0
+ etab = -1.7142866e-5
+ vsat = 85658.6
+ tcjsw = 0.000645489
+ lnfactor = 0.0
+ wint = 3e-9
+ vth0 = 0.479324
+ rdsw = 170.0
+ pvoff = 0.0
+ lint = 1e-8
+ wmax = 0.000900001
+ wmin = 1e-5
+ cdscb = 0.0
+ cdscd = 0.0
+ lkt1 = 5.782678e-9
+ lkt2 = 1.5570838e-9
+ peta0 = 1.0000000000000001e-20
+ lmax = 1.2e-6
+ lpdiblc2 = 1.525682e-9
+ lmin = 5e-7
+ pvth0 = 0.0
+ ags = 0.0462474
+ drout = 0.0
+ tpbsw = 0.001554306
+ cit = -0.00015788565
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ dlc = 3e-9
+ cjswg = 3.340547e-10
+ k3b = 0.0
+ pscbe1 = 400000100.0
+ pscbe2 = 1e-6
+ mjswg = 0.43879
+ dwb = 0.0
+ dwg = 0.0
+ hdif = 2e-7
+ lua1 = -3.0446746e-18
+ lub1 = -1.2004175e-24
+ luc1 = -6.517273e-17
+ wvoff = 0.0
+ mjsw = 0.2003879
+ nqsmod = 0
+ tpbswg = 0.001554306
+ noimod = 2
+ nfactor = 1.0
+ lute = -2.6630502e-7
+ weta0 = 0
+ la0 = 4.581426e-7
+ wvsat = 0.0
+ jsw = 1.45e-12
+ kt1 = -0.2290285
+ lk1 = -7.214246e-9
+ kt2 = -0.031611919
+ lk2 = 1.703151e-9
+ lpclm = 1.5245718e-7
+ wvth0 = 0.0
+ a0 = -0.2911571
+ a1 = 0.0
+ a2 = 0.99
+ b0 = 0.0
+ b1 = 0.0
+ llc = -0.039
+ cdsc = 0.0
+ lln = -1
+ lu0 = 1.0406079e-9
+ at = 20000.0
+ cf = 0
+ cj = 0.001000266
+ ef = 0.874
+ k1 = 0.5318048
+ k2 = 0.004864913
+ k3 = 0.0
+ em = 30000000.0
+ lua = 7.982966e-17
+ lub = -1.5630905e-25
+ luc = -9.669895e-18
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ js = 3.5e-7
+ cgdo = 3.665e-10
+ ll = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0016847569
+ u0 = 0.04381358
+ pb = 0.6882682
+ w0 = 0.0
+ rd = 0
+ nlx = 0.0
+ rs = 0
+ pdiblcb = 0.01
+ ua = -1.0347512e-9
+ ub = 3.0100842e-18
+ uc = 1.4678947e-10
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ cgso = 3.665e-10
+ pu0 = 0.0
+ prt = 0
+ cjsw = 2.040547e-10
+ binunit = 2
+ rsh = 6.8
+ tcj = 0.001040287
+ ua1 = 1.2266247e-9
+ ub1 = -8.574386e-20
+ uc1 = 6.788683e-11
+ lketa = -8.954029e-9
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ tpb = 0.001554306
+ tox = 4.08e-9
+ capmod = 3
+ xpart = 1
+ ute = -1.3504703
+ tnom = 25.0
+ wln = 1.0
+ wu0 = 0.0
+ pbswg = 0.6882682
+ wwl = 0.0
+ wwn = 1
+ xti = 3
+ toxm = 4.08e-9
+ mobmod = 1
+ lvoff = 1.5735258e-8
+ pbsw = 0.6882682
+ pclm = 0.8687172
+ )

.model nch_mc_4 nmos (
+ level = 49
+ lua1 = 8.039099e-19
+ lub1 = 3.824101e-25
+ luc1 = 2.9606131e-17
+ mjsw = 0.2003879
+ lute = 7.030476e-8
+ ags = -0.019916179
+ tcjsw = 0.000645489
+ nfactor = 1.0
+ cdsc = 0.0
+ cit = 0.000271889
+ pvoff = 0.0
+ dlc = 3e-9
+ cgdo = 3.665e-10
+ k3b = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cgso = 3.665e-10
+ peta0 = 1.0000000000000001e-20
+ pdiblc1 = 1e-6
+ pdiblc2 = -0.00593541
+ pdiblcb = 0.01
+ pvth0 = 0.0
+ drout = 0.0
+ alpha0 = 0.0
+ cjsw = 2.040547e-10
+ alpha1 = 0.448150714
+ tpbsw = 0.001554306
+ la0 = 7.545271e-8
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ pscbe1 = 400000000.0
+ pscbe2 = 1e-6
+ binunit = 2
+ jsw = 1.45e-12
+ kt1 = -0.22715
+ lk1 = 4.899558e-8
+ kt2 = -0.029537767
+ lk2 = -2.3341336e-8
+ cjswg = 3.340547e-10
+ pnfactor = 0.0
+ llc = -0.039
+ lln = -1
+ mjswg = 0.43879
+ lu0 = 1.2517989e-9
+ wnfactor = 0.0
+ lua = -1.0530929e-18
+ lub = 5.559478e-27
+ luc = 4.133919e-18
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ tnom = 25.0
+ nqsmod = 0
+ tpbswg = 0.001554306
+ wvoff = 0.0
+ nlx = 0.0
+ noimod = 2
+ toxm = 4.08e-9
+ pu0 = 0.0
+ weta0 = 0
+ pbsw = 0.6882682
+ pclm = 1.1076791
+ prt = 0
+ wvsat = 0.0
+ lnfactor = 0.0
+ lpclm = 4.253467e-8
+ wvth0 = 0.0
+ rsh = 6.8
+ tcj = 0.001040287
+ ua1 = 1.2182583e-9
+ ub1 = -3.526674e-18
+ uc1 = -1.381542e-10
+ tpb = 0.001554306
+ tox = 4.08e-9
+ ute = -2.0822308
+ version = 3.24
+ wln = 1.0
+ wu0 = 0.0
+ lpdiblc2 = 5.030957e-9
+ wwl = 0.0
+ wwn = 1
+ xti = 3
+ keta = -0.04182327
+ capmod = 3
+ dsub = 0.0
+ lketa = 2.9580252e-9
+ xpart = 1
+ lags = -1.1735286e-11
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ lcit = 1.0493098e-10
+ voff = -0.1245498
+ pbswg = 0.6882682
+ mobmod = 1
+ ldif = 9e-8
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ lvoff = -1.5463618e-9
+ eta0 = -0.0002937502
+ pvag = 0.0
+ etab = 0.0013875004
+ beta0 = 11.59263
+ vsat = 84438.96
+ wint = 3e-9
+ leta0 = 1.8113305999999998e-10
+ vth0 = 0.4752311
+ letab = -6.842502e-10
+ rdsw = 170.0
+ lvsat = -0.00020125005
+ lint = 1e-8
+ lvth0 = 5.825501e-9
+ wmax = 0.000900001
+ wmin = 1e-5
+ lkt1 = 4.918561e-9
+ lkt2 = 6.029743e-10
+ delta = 0.01
+ lmax = 5e-7
+ a0 = 0.5407774
+ a1 = 0.0
+ a2 = 0.99
+ b0 = 0.0
+ b1 = 0.0
+ lmin = 1.8e-7
+ at = 20000.0
+ cf = 0
+ cj = 0.001000266
+ ef = 0.874
+ k1 = 0.4096095
+ k2 = 0.05930946
+ k3 = 0.0
+ em = 30000000.0
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ js = 3.5e-7
+ ll = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ u0 = 0.04335447
+ pb = 0.6882682
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ua = -8.589192e-10
+ ub = 2.6581962e-18
+ uc = 1.1678118e-10
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ tcjswg = 0.000645489
+ hdif = 2e-7
+ )

.model nch_mc_5 nmos (
+ level = 49
+ pu0 = 0.0
+ pscbe1 = 200000030.0
+ pscbe2 = 1e-6
+ tpbsw = 0.001554306
+ prt = 0
+ dsub = 0.0
+ cjswg = 3.340547e-10
+ rsh = 6.8
+ tcj = 0.001040287
+ ua1 = 1.224e-9
+ ub1 = -1.0684574e-18
+ a0 = 0.3702259
+ a1 = 0.0
+ a2 = 0.99
+ uc1 = 2.4230474e-11
+ b0 = 0.0
+ b1 = 0.0
+ mjswg = 0.43879
+ nqsmod = 0
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ tpbswg = 0.001554306
+ at = 20000.0
+ cf = 0
+ cj = 0.001000266
+ ef = 0.874
+ k1 = 0.5102321
+ k2 = 0.016091494
+ k3 = 0.0
+ tpb = 0.001554306
+ noimod = 2
+ em = 30000000.0
+ tox = 4.08e-9
+ js = 3.5e-7
+ wa0 = -1.4643313e-9
+ ll = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ wvoff = 8.907224e-10
+ u0 = 0.0430359
+ pb = 0.6882682
+ w0 = 0.0
+ rd = 0
+ ute = -1.5803809
+ rs = 0
+ ua = -5.885942e-10
+ ub = 2.3329335e-18
+ uc = 1.1057788e-10
+ voff = -0.1406671
+ wk1 = 3.995606e-8
+ wk2 = -1.2928737e-8
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -2e-8
+ ww = 0.0
+ ldif = 9e-8
+ xw = 0.0
+ wln = 1.0
+ wu0 = -8.320099e-9
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ puc1 = -1.4905616e-28
+ weta0 = 0
+ wua = -2.3665659e-16
+ wub = -1.936796e-25
+ wuc = -1.815927e-17
+ wwl = 0.0
+ wwn = 1
+ eta0 = 5e-5
+ xti = 3
+ wvsat = 0.0
+ pvag = 0.0
+ etab = -5e-5
+ vsat = 90000.01
+ wvth0 = 6.876114e-10
+ wint = 3e-9
+ vth0 = 0.4364873
+ rdsw = 170.0
+ wkt1 = -8.215166e-9
+ wkt2 = 1.6245854e-9
+ lint = 1e-8
+ wmax = 1e-5
+ wmin = 1.2e-6
+ lmax = 2.0001e-5
+ lmin = 1e-5
+ capmod = 3
+ xpart = 1
+ wub1 = -5.244247e-25
+ pnfactor = 0.0
+ wuc1 = -1.257911e-16
+ wnfactor = 0.0
+ hdif = 2e-7
+ mobmod = 1
+ wute = 3.808433e-9
+ pbswg = 0.6882682
+ mjsw = 0.2003879
+ lvoff = 0.0
+ beta0 = 11.59263
+ lnfactor = 0.0
+ leta0 = 8e-15
+ cdsc = 0.0
+ nfactor = 1.0
+ lvth0 = 0.0
+ cgdo = 3.665e-10
+ cgso = 3.665e-10
+ delta = 0.01
+ dvt0w = 0.0
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0006999999
+ dvt1w = 0.0
+ dvt2w = 0.0
+ pdiblcb = 0.01
+ cjsw = 2.040547e-10
+ tcjswg = 0.000645489
+ ags = 0.02
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ cit = -0.00010000001
+ binunit = 2
+ dlc = 3e-9
+ tnom = 25.0
+ k3b = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ toxm = 4.08e-9
+ pbsw = 0.6882682
+ pclm = 0.8000001
+ tcjsw = 0.000645489
+ pvoff = 0.0
+ jsw = 1.45e-12
+ kt1 = -0.2232244
+ kt2 = -0.030428693
+ lk2 = 0.0
+ llc = -0.039
+ lln = -1
+ lu0 = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ nch = 3.9e+17
+ peta0 = 1.0000000000000001e-20
+ lwl = 0.0
+ lwn = 1.0
+ nlx = 0.0
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ version = 3.24
+ wketa = -1.0935369e-8
+ pvth0 = 0.0
+ keta = 0.010357677
+ drout = 0.0
+ )

.model nch_mc_6 nmos (
+ level = 49
+ nfactor = 1.0
+ cgso = 3.665e-10
+ capmod = 3
+ cjsw = 2.040547e-10
+ lketa = -4.518989e-8
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0003968181
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ pdiblcb = 0.01
+ lpscbe1 = 262.58185
+ xpart = 1
+ mobmod = 1
+ tnom = 25.0
+ pbswg = 0.6882682
+ binunit = 2
+ toxm = 4.08e-9
+ lvoff = -1.0806052e-8
+ a0 = 0.40626
+ a1 = 0.0
+ a2 = 0.99
+ b0 = 0.0
+ b1 = 0.0
+ pbsw = 0.6882682
+ pclm = 0.7755287
+ at = 20000.0
+ cf = 0
+ cj = 0.001000266
+ ef = 0.874
+ k1 = 0.508509
+ beta0 = 11.59263
+ k2 = 0.01731023
+ k3 = 0.0
+ em = 30000000.0
+ js = 3.5e-7
+ ll = 0.0
+ leta0 = 8e-15
+ mj = 0.3595262
+ lw = 0.0
+ u0 = 0.04273027
+ pb = 0.6882682
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ags = 0.02
+ ua = -5.377125e-10
+ ub = 2.2537915e-18
+ uc = 1.0657759e-10
+ lvsat = -0.006753025
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ lvth0 = 6.070609e-8
+ cit = -0.00012675911
+ ppclm = 1.9027247e-13
+ delta = 0.01
+ dlc = 3e-9
+ k3b = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ tcjswg = 0.000645489
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ pkt1 = 4.710912e-15
+ pkt2 = -4.130377e-15
+ keta = 0.014894814
+ version = 3.24
+ dsub = 0.0
+ pnfactor = 0.0
+ la0 = -3.588995e-7
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ wnfactor = 0.0
+ jsw = 1.45e-12
+ lk1 = 1.7161611e-8
+ kt1 = -0.2231775
+ lk2 = -1.2138612e-8
+ kt2 = -0.030469729
+ pketa = 1.9809019e-14
+ llc = -0.039
+ lln = -1
+ lu0 = 3.0440912e-9
+ lcit = 2.6652053e-10
+ voff = -0.1395822
+ lua = -5.067804e-16
+ lub = 7.882536e-25
+ luc = 3.984287e-17
+ nch = 3.9e+17
+ ldif = 9e-8
+ lwl = 0.0
+ lwn = 1.0
+ wpclm = -1.9103656e-8
+ kt1l = 0.0
+ pa0 = 9.284546e-14
+ prwb = 0.0
+ prwg = 0.0
+ pub1 = 4.176128e-31
+ nlx = 0.0
+ puc1 = 7.417578e-23
+ eta0 = 5e-5
+ pk1 = -2.2514154e-14
+ pk2 = 1.0246181e-14
+ pvag = 0.0
+ etab = -5e-5
+ tcjsw = 0.000645489
+ pu0 = 2.4756895e-15
+ vsat = 90678.02
+ lnfactor = 0.0
+ wint = 3e-9
+ pute = -5.708167e-14
+ prt = 0
+ pua = 4.243342e-22
+ pub = -5.065558e-31
+ puc = -8.588134e-24
+ vth0 = 0.4303924
+ rdsw = 170.0
+ pvoff = 3.345241e-15
+ wkt1 = -8.688151e-9
+ wkt2 = 2.0392819e-9
+ rsh = 6.8
+ lint = 1e-8
+ tcj = 0.001040287
+ ua1 = 1.224e-9
+ ub1 = -1.0643074e-18
+ uc1 = 2.4967807e-11
+ wmax = 1e-5
+ wmin = 1.2e-6
+ cdscb = 0.0
+ cdscd = 0.0
+ tpb = 0.001554306
+ peta0 = 1.0000000000000001e-20
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ tox = 4.08e-9
+ lkt1 = -4.674615e-10
+ lkt2 = 4.087321e-10
+ wa0 = -1.0786144e-8
+ lpdiblc2 = 3.0196912e-9
+ lmax = 1e-5
+ pvsat = 1.9027204e-9
+ ute = -1.5809486
+ pscbe1 = 173636400.0
+ pscbe2 = 1e-6
+ wk1 = 4.221652e-8
+ wk2 = -1.3957471e-8
+ lmin = 1.2e-6
+ wketa = -1.292423e-8
+ pvth0 = -9.316875e-16
+ wln = 1.0
+ drout = 0.0
+ wu0 = -8.568663e-9
+ tpbsw = 0.001554306
+ wua = -2.7926046e-16
+ wub = -1.4282058e-25
+ wuc = -1.7297008e-17
+ wwl = 0.0
+ wwn = 1
+ xti = 3
+ nqsmod = 0
+ tpbswg = 0.001554306
+ cjswg = 3.340547e-10
+ noimod = 2
+ wub1 = -5.663537e-25
+ wuc1 = -1.3323848e-16
+ mjswg = 0.43879
+ hdif = 2e-7
+ wvoff = 5.548539e-10
+ lub1 = -4.133362e-26
+ luc1 = -7.343755e-18
+ wute = 9.539526e-9
+ mjsw = 0.2003879
+ weta0 = 0
+ lute = 5.654154e-9
+ wvsat = -0.00019104627
+ lpclm = 2.4373449e-7
+ wvth0 = 7.811502e-10
+ cdsc = 0.0
+ cgdo = 3.665e-10
+ )

.model nch_mc_7 nmos (
+ level = 49
+ beta0 = 11.59263
+ pvag = 0.0
+ etab = -1.7142869e-5
+ vsat = 85513.59
+ leta0 = 3.812228e-11
+ wint = 3e-9
+ pute = 4.357466e-13
+ letab = -3.811428e-11
+ vth0 = 0.4799949
+ lvsat = -0.0007622865
+ rdsw = 170.0
+ lvth0 = 3.167132e-9
+ wkt1 = -3.681822e-9
+ wkt2 = -1.3190541e-9
+ lint = 1e-8
+ wmax = 1e-5
+ la0 = 4.645035e-7
+ ppclm = 7.258032e-15
+ wmin = 1.2e-6
+ jsw = 1.45e-12
+ lk1 = -1.1179709e-8
+ kt1 = -0.2286601
+ lk2 = 3.431065e-9
+ kt2 = -0.031479932
+ delta = 0.01
+ tcjswg = 0.000645489
+ lkt1 = 5.892387e-9
+ lkt2 = 1.5805686e-9
+ llc = -0.039
+ lln = -1
+ lmax = 1.2e-6
+ lu0 = 9.604713e-10
+ lmin = 5e-7
+ lua = 6.148926e-17
+ lub = -1.2783527e-25
+ luc = -6.505068e-18
+ nch = 3.9e+17
+ dvt0w = 0.0
+ lwl = 0.0
+ lwn = 1.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ pa0 = -6.357063e-14
+ nlx = 0.0
+ pk1 = 3.963084e-14
+ pk2 = -1.7268767e-14
+ pu0 = 8.008865e-16
+ prt = 0
+ pua = 1.8329395e-22
+ pub = -2.8456703e-31
+ puc = -3.16293e-23
+ wua1 = -3.55913e-18
+ wub1 = -1.6132161e-24
+ wuc1 = -1.8047248e-16
+ hdif = 2e-7
+ rsh = 6.8
+ pketa = 9.843987e-15
+ tcj = 0.001040287
+ ua1 = 1.2269809e-9
+ ub1 = 7.567455e-20
+ lua1 = -3.457781e-18
+ uc1 = 8.594492e-11
+ lub1 = -1.3637128e-24
+ luc1 = -7.807721e-17
+ wute = -4.153124e-7
+ mjsw = 0.2003879
+ tpb = 0.001554306
+ tox = 4.08e-9
+ wa0 = 1.2405528e-7
+ wpclm = 1.3866737e-7
+ ute = -1.3089141
+ lute = -3.0990586e-7
+ wk1 = -1.1356744e-8
+ wk2 = 9.762311e-9
+ wln = 1.0
+ tcjsw = 0.000645489
+ wu0 = -7.124867e-9
+ wua = -7.146715e-17
+ wub = -3.341902e-25
+ wuc = 2.5660584e-18
+ wwl = 0.0
+ wwn = 1
+ xti = 3
+ cdsc = 0.0
+ pvoff = -3.013814e-15
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ cgdo = 3.665e-10
+ a0 = -0.3035701
+ a1 = 0.0
+ a2 = 0.99
+ b0 = 0.0
+ b1 = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 1.0000000000000001e-20
+ at = 20000.0
+ cf = 0
+ cj = 0.001000266
+ pscbe1 = 400000100.0
+ pscbe2 = 1e-6
+ ef = 0.874
+ k1 = 0.5329412
+ k2 = 0.003888095
+ k3 = 0.0
+ em = 30000000.0
+ cgso = 3.665e-10
+ js = 3.5e-7
+ ll = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ u0 = 0.04452649
+ pb = 0.6882682
+ nfactor = 1.0
+ w0 = 0.0
+ rd = 0
+ wketa = -4.333682e-9
+ rs = 0
+ ua = -1.0276002e-9
+ ub = 3.0435232e-18
+ uc = 1.4653272e-10
+ pvth0 = 7.751598e-15
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ drout = 0.0
+ tpbsw = 0.001554306
+ nqsmod = 0
+ cjsw = 2.040547e-10
+ tpbswg = 0.001554306
+ noimod = 2
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ cjswg = 3.340547e-10
+ pnfactor = 0.0
+ mjswg = 0.43879
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0017737894
+ pdiblcb = 0.01
+ wnfactor = 0.0
+ tnom = 25.0
+ wvoff = 6.036798e-9
+ pags = 4.128623e-14
+ toxm = 4.08e-9
+ weta0 = 0
+ ppdiblc2 = 1.0321563e-15
+ binunit = 2
+ pbsw = 0.6882682
+ pclm = 0.8548421
+ wvsat = 0.0014492224
+ wpdiblc2 = -8.897895e-10
+ lpclm = 1.5173094e-7
+ wvth0 = -6.704436e-9
+ lnfactor = 0.0
+ capmod = 3
+ lpdiblc2 = 1.4224044e-9
+ pkt1 = -1.0964308e-15
+ pkt2 = -2.3470743e-16
+ keta = -0.01549387
+ lketa = -9.939018e-9
+ mobmod = 1
+ wags = -3.559157e-8
+ dsub = 0.0
+ version = 3.24
+ xpart = 1
+ ags = 0.04980868
+ lags = -3.457808e-8
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ cit = -0.00015788565
+ pbswg = 0.6882682
+ lcit = 3.0262734e-10
+ voff = -0.1627226
+ ldif = 9e-8
+ dlc = 3e-9
+ k3b = 0.0
+ kt1l = 0.0
+ lvoff = 1.6036822e-8
+ pua1 = 4.128591e-24
+ prwb = 0.0
+ prwg = 0.0
+ pub1 = 1.6319734e-30
+ puc1 = 1.2896722e-22
+ dwb = 0.0
+ dwg = 0.0
+ eta0 = 1.7142869e-5
+ )

.model nch_mc_8 nmos (
+ level = 49
+ pketa = -2.7027957e-15
+ tnom = 25.0
+ pdiblc1 = 1e-6
+ pdiblc2 = -0.006119013
+ pdiblcb = 0.01
+ pags = -1.0838496e-14
+ toxm = 4.08e-9
+ wpclm = 6.656068e-8
+ pcit = 1.4220811e-17
+ pbsw = 0.6882682
+ pclm = 1.1010191
+ tcjsw = 0.000645489
+ binunit = 2
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ pvoff = -9.75415e-16
+ pscbe1 = 400000000.0
+ pscbe2 = 1e-6
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = -1.3721218e-18
+ petab = 1.6959704e-18
+ pvsat = 1.5350395e-12
+ wketa = 2.2941933e-8
+ nqsmod = 0
+ pvth0 = 4.508938e-15
+ tpbswg = 0.001554306
+ drout = 0.0
+ noimod = 2
+ pkt1 = -1.7512235e-15
+ pkt2 = 7.382567e-17
+ keta = -0.04411884
+ tpbsw = 0.001554306
+ wags = 7.772305e-8
+ dsub = 0.0
+ cjswg = 3.340547e-10
+ mjswg = 0.43879
+ lags = 1.0727657e-9
+ wcit = -3.0914837e-11
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ version = 3.24
+ wvoff = 1.6054964e-9
+ lcit = 1.0350804e-10
+ voff = -0.1247105
+ ldif = 9e-8
+ weta0 = 3.0046217e-12
+ kt1l = 0.0
+ pua1 = -1.0901051e-24
+ prwb = 0.0
+ prwg = 0.0
+ pub1 = -4.238914e-31
+ puc1 = -2.7204607e-23
+ wetab = -3.686654e-12
+ wvsat = 0.0014459029
+ eta0 = -0.00029405078
+ pvag = 0.0
+ etab = 0.0013878694
+ lpclm = 3.848953e-8
+ wvth0 = 3.448236e-10
+ vsat = 84294.28
+ wint = 3e-9
+ pute = -1.178615e-13
+ vth0 = 0.4751966
+ rdsw = 170.0
+ capmod = 3
+ wkt1 = -2.2583577e-9
+ wkt2 = -1.9897783e-9
+ lint = 1e-8
+ ags = -0.027693154
+ wmax = 1e-5
+ wmin = 1.2e-6
+ lkt1 = 5.093789e-9
+ lkt2 = 5.955873e-10
+ lmax = 5e-7
+ cit = 0.00027498236
+ lmin = 1.8e-7
+ dlc = 3e-9
+ mobmod = 1
+ k3b = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ a0 = 0.5262308
+ a1 = 0.0
+ a2 = 0.99
+ lketa = 3.228467e-9
+ b0 = 0.0
+ b1 = 0.0
+ at = 20000.0
+ cf = 0
+ cj = 0.001000266
+ ef = 0.874
+ k1 = 0.4007356
+ k2 = 0.0631886
+ k3 = 0.0
+ em = 30000000.0
+ xpart = 1
+ js = 3.5e-7
+ ll = 0.0
+ pnfactor = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ u0 = 0.04384084
+ wua1 = 7.785862e-18
+ pb = 0.6882682
+ wub1 = 2.8560549e-24
+ w0 = 0.0
+ wuc1 = 1.5903152e-16
+ rd = 0
+ rs = 0
+ ua = -9.017296e-10
+ ub = 2.7527719e-18
+ uc = 1.2291169e-10
+ wnfactor = 0.0
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ hdif = 2e-7
+ lua1 = 9.129858e-19
+ lub1 = 4.248247e-25
+ la0 = 8.279508e-8
+ luc1 = 3.232822e-17
+ pbswg = 0.6882682
+ wute = 7.881835e-7
+ mjsw = 0.2003879
+ jsw = 1.45e-12
+ lk1 = 4.963488e-8
+ kt1 = -0.226924
+ lk2 = -2.3847164e-8
+ kt2 = -0.029338669
+ llc = -0.039
+ lvoff = -1.4487617e-9
+ lln = -1
+ lu0 = 1.2758692e-9
+ ppdiblc2 = -2.2121929e-16
+ lute = 8.209799e-8
+ lua = 3.588764e-18
+ lub = 5.910339e-27
+ luc = 4.360599e-18
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ wpdiblc2 = 1.8349379e-9
+ beta0 = 11.59263
+ pa0 = -7.337964e-14
+ lnfactor = 0.0
+ nlx = 0.0
+ leta0 = 1.8127133999999998e-10
+ letab = -6.844199e-10
+ pk1 = -6.389182e-15
+ pk2 = 5.055259e-15
+ lvsat = -0.00020140363
+ cdsc = 0.0
+ pu0 = -2.4055863e-16
+ lvth0 = 5.374336e-9
+ prt = 0
+ pua = -4.639069e-23
+ pub = -3.506499e-33
+ puc = -2.2654354e-24
+ cgdo = 3.665e-10
+ tcjswg = 0.000645489
+ ppclm = 4.042711e-14
+ delta = 0.01
+ cgso = 3.665e-10
+ rsh = 6.8
+ tcj = 0.001040287
+ lpdiblc2 = 5.053093e-9
+ ua1 = 1.2174792e-9
+ ub1 = -3.81245e-18
+ uc1 = -1.540669e-10
+ tpb = 0.001554306
+ tox = 4.08e-9
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ wa0 = 1.4537927e-7
+ nfactor = 1.0
+ ute = -2.1610963
+ cjsw = 2.040547e-10
+ wk1 = 8.868675e-8
+ wk2 = -3.876818e-8
+ wln = 1.0
+ wu0 = -4.860856e-9
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ wua = 4.278473e-16
+ wub = -9.451913e-25
+ wuc = -6.126842e-17
+ wwl = 0.0
+ wwn = 1
+ xti = 3
+ )

.model nch_mc_9 nmos (
+ level = 49
+ cjswg = 3.340547e-10
+ mjswg = 0.43879
+ wub1 = -7.675553e-27
+ wuc1 = -1.4706552e-17
+ hdif = 2e-7
+ wvoff = -8.66569e-10
+ ags = 0.02
+ wute = 3.836007e-8
+ mjsw = 0.2003879
+ weta0 = 0
+ cit = -0.00010000004
+ wvsat = 0.0
+ dlc = 3e-9
+ k3b = 0.0
+ wvth0 = -4.263109e-9
+ dwb = 0.0
+ dwg = 0.0
+ capmod = 3
+ cdsc = 0.0
+ cgdo = 3.665e-10
+ cgso = 3.665e-10
+ mobmod = 1
+ jsw = 1.45e-12
+ kt1 = -0.2313184
+ lk2 = 0.0
+ kt2 = -0.029076951
+ llc = -0.039
+ lln = -1
+ lu0 = 0.0
+ cjsw = 2.040547e-10
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ nlx = 0.0
+ nfactor = 1.0
+ xpart = 1
+ pu0 = 0.0
+ prt = 0
+ tnom = 25.0
+ pbswg = 0.6882682
+ rsh = 6.8
+ tcj = 0.001040287
+ ua1 = 1.224e-9
+ pdiblc1 = 1e-6
+ toxm = 4.08e-9
+ pdiblc2 = 0.0007000003
+ ub1 = -1.5012456e-18
+ lvoff = 0.0
+ uc1 = -6.880516e-11
+ pdiblcb = 0.01
+ pbsw = 0.6882682
+ tpb = 0.001554306
+ pclm = 0.8000001
+ tox = 4.08e-9
+ beta0 = 11.59263
+ wa0 = 7.667051e-8
+ leta0 = 8e-15
+ ute = -1.6093186
+ wk1 = -2.074723e-8
+ wk2 = 4.920634e-9
+ tcjswg = 0.000645489
+ wln = 1.0
+ wu0 = 1.0362965e-9
+ lvth0 = 0.0
+ binunit = 2
+ wua = 1.4309126e-16
+ wub = -1.5411778e-25
+ wuc = -1.4141237e-17
+ wwl = 0.0
+ wwn = 1
+ xti = 3
+ delta = 0.01
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ keta = 0.0010152902
+ dsub = 0.0
+ pnfactor = 0.0
+ wnfactor = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ a0 = 0.3047864
+ a1 = 0.0
+ a2 = 0.99
+ b0 = 0.0
+ b1 = 0.0
+ voff = -0.1391954
+ version = 3.24
+ at = 20000.0
+ cf = 0
+ cj = 0.001000266
+ ldif = 9e-8
+ ef = 0.874
+ k1 = 0.5610723
+ k2 = 0.0011422717
+ k3 = 0.0
+ em = 30000000.0
+ kt1l = 0.0
+ js = 3.5e-7
+ prwb = 0.0
+ ll = 0.0
+ prwg = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ u0 = 0.03519972
+ pb = 0.6882682
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ua = -9.066409e-10
+ ub = 2.2997995e-18
+ uc = 1.072127e-10
+ eta0 = 5e-5
+ wl = 0.0
+ tcjsw = 0.000645489
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -2e-8
+ ww = 0.0
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ xw = 0.0
+ pvag = 0.0
+ etab = -5e-5
+ lnfactor = 0.0
+ vsat = 90000.01
+ wint = 3e-9
+ pscbe1 = 200000030.0
+ pscbe2 = 1e-6
+ vth0 = 0.4406337
+ pvoff = 0.0
+ rdsw = 170.0
+ wkt1 = 1.4490446e-9
+ wkt2 = 1.0605161e-11
+ lint = 1e-8
+ wmax = 1.2e-6
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 1.0000000000000001e-20
+ wmin = 5e-7
+ nqsmod = 0
+ tpbswg = 0.001554306
+ noimod = 2
+ lmax = 2.0001e-5
+ wketa = 2.1944087e-10
+ pvth0 = 0.0
+ lmin = 1e-5
+ drout = 0.0
+ tpbsw = 0.001554306
+ )

.model nch_mc_10 nmos (
+ level = 49
+ lute = -1.2190513e-8
+ nqsmod = 0
+ tpbswg = 0.001554306
+ noimod = 2
+ cdsc = 0.0
+ cgdo = 3.665e-10
+ nfactor = 1.0
+ lketa = -2.8027248e-8
+ cgso = 3.665e-10
+ xpart = 1
+ cjsw = 2.040547e-10
+ pbswg = 0.6882682
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0003968185
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ pdiblcb = 0.01
+ lpscbe1 = 262.58185
+ lvoff = -3.602222e-9
+ capmod = 3
+ beta0 = 11.59263
+ tnom = 25.0
+ leta0 = 8e-15
+ binunit = 2
+ lvsat = -0.006201102
+ toxm = 4.08e-9
+ lvth0 = 6.592048e-8
+ pcit = 4.302753e-19
+ pbsw = 0.6882682
+ pclm = 0.7699873
+ ppclm = 1.243718e-13
+ mobmod = 1
+ delta = 0.01
+ ags = 0.02
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ cit = -0.00012672294
+ dlc = 3e-9
+ k3b = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ pnfactor = 0.0
+ pkt1 = 7.833639e-15
+ pkt2 = 9.747044e-16
+ keta = 0.00382927
+ wnfactor = 0.0
+ pketa = -6.831802e-16
+ version = 3.24
+ dsub = 0.0
+ wpclm = -1.2487239e-8
+ wcit = -4.317371e-14
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ la0 = -1.9725388e-7
+ tcjsw = 0.000645489
+ jsw = 1.45e-12
+ tcjswg = 0.000645489
+ lk1 = 1.0512358e-8
+ kt1 = -0.2310088
+ lk2 = -5.410051e-9
+ kt2 = -0.028688708
+ lcit = 2.6616018e-10
+ llc = -0.039
+ lln = -1
+ voff = -0.1388337
+ lu0 = 3.705752e-9
+ lnfactor = 0.0
+ ldif = 9e-8
+ lua = -1.9124487e-16
+ lub = 4.117038e-25
+ luc = 4.038815e-17
+ nch = 3.9e+17
+ pvoff = -5.256132e-15
+ lwl = 0.0
+ lwn = 1.0
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ pub1 = -1.8996434e-32
+ puc1 = 1.3569954e-23
+ pa0 = -1.0015934e-13
+ nlx = 0.0
+ eta0 = 5e-5
+ pk1 = -1.457495e-14
+ pk2 = 2.2122807e-15
+ pvag = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ etab = -5e-5
+ peta0 = 1.0000000000000001e-20
+ vsat = 90622.61
+ wint = 3e-9
+ pu0 = 1.6856667e-15
+ pute = -3.577514e-14
+ pvsat = 1.2437262e-9
+ vth0 = 0.4340151
+ prt = 0
+ pua = 4.758471e-23
+ pub = -5.695533e-32
+ puc = -9.239189e-24
+ lpdiblc2 = 3.0196912e-9
+ wketa = 2.8803285e-10
+ rdsw = 170.0
+ pvth0 = -7.157672e-15
+ wkt1 = 6.625341e-10
+ wkt2 = -8.725676e-11
+ drout = 0.0
+ lint = 1e-8
+ rsh = 6.8
+ tpbsw = 0.001554306
+ wmax = 1.2e-6
+ tcj = 0.001040287
+ ua1 = 1.224e-9
+ ub1 = -1.5338095e-18
+ uc1 = -7.316409e-11
+ wmin = 5e-7
+ lkt1 = -3.0828107e-9
+ lkt2 = -3.866881e-9
+ tpb = 0.001554306
+ tox = 4.08e-9
+ cjswg = 3.340547e-10
+ lmax = 1e-5
+ wa0 = 8.672666e-8
+ lmin = 1.2e-6
+ ute = -1.6080947
+ mjswg = 0.43879
+ wk1 = -1.9283881e-8
+ wk2 = 4.698517e-9
+ wln = 1.0
+ wu0 = 8.670528e-10
+ wvoff = -3.388445e-10
+ wua = 1.3831368e-16
+ wub = -1.4839938e-25
+ wuc = -1.3213606e-17
+ wwl = 0.0
+ wwn = 1
+ xti = 3
+ a0 = 0.324591
+ a1 = 0.0
+ a2 = 0.99
+ b0 = 0.0
+ b1 = 0.0
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ wub1 = -5.768295e-27
+ wuc1 = -1.6068998e-17
+ weta0 = 0
+ at = 20000.0
+ cf = 0
+ cj = 0.001000266
+ ef = 0.874
+ k1 = 0.5600169
+ k2 = 0.0016854487
+ k3 = 0.0
+ em = 30000000.0
+ hdif = 2e-7
+ wvsat = -0.00012487893
+ js = 3.5e-7
+ pscbe1 = 173636400.0
+ pscbe2 = 1e-6
+ ll = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ u0 = 0.03482766
+ pb = 0.6882682
+ lub1 = 3.243357e-25
+ lpclm = 2.9892766e-7
+ wvth0 = -3.544466e-9
+ luc1 = 4.341489e-17
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ wute = 4.195195e-8
+ ua = -8.874397e-10
+ ub = 2.2584638e-18
+ uc = 1.0315766e-10
+ mjsw = 0.2003879
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ )

.model nch_mc_11 nmos (
+ level = 49
+ lvoff = 1.116323e-8
+ wcit = 5.431231e-13
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ ags = 0.02
+ beta0 = 11.59263
+ leta0 = 3.8122299999999996e-11
+ lcit = 3.0283653e-10
+ cit = -0.0001583405
+ letab = -3.81143e-11
+ voff = -0.1515625
+ ldif = 9e-8
+ lvsat = -0.0007659488
+ dlc = 3e-9
+ kt1l = 0.0
+ mobmod = 1
+ prwb = 0.0
+ lvth0 = 1.0109751e-8
+ prwg = 0.0
+ pub1 = -5.874811e-31
+ puc1 = -3.67348e-23
+ a0 = -0.1914371
+ a1 = 0.0
+ a2 = 0.99
+ k3b = 0.0
+ b0 = 0.0
+ b1 = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ eta0 = 1.7142847e-5
+ at = 20000.0
+ cf = 0
+ cj = 0.001000266
+ ef = 0.874
+ k1 = 0.5552615
+ ppclm = 7.308824e-14
+ k2 = 0.003544799
+ k3 = 0.0
+ em = 30000000.0
+ pvag = 0.0
+ etab = -1.7142847e-5
+ delta = 0.01
+ js = 3.5e-7
+ vsat = 85937.13
+ ll = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ u0 = 0.03581186
+ pb = 0.6882682
+ wint = 3e-9
+ pute = -2.0303331e-13
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ua = -1.3333591e-9
+ ub = 2.969086e-18
+ uc = 1.6160392e-10
+ vth0 = 0.4821278
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ rdsw = 170.0
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ wkt1 = 1.1898274e-8
+ wkt2 = 2.0987987e-9
+ lint = 1e-8
+ wmax = 1.2e-6
+ la0 = 4.013388e-7
+ wmin = 5e-7
+ lkt1 = 9.329063e-9
+ lkt2 = 2.691467e-9
+ jsw = 1.45e-12
+ lk1 = 1.6028618e-8
+ kt1 = -0.2417087
+ lk2 = -7.566896e-9
+ kt2 = -0.03434246
+ lmax = 1.2e-6
+ llc = -0.039
+ lln = -1
+ lu0 = 2.5640821e-9
+ lmin = 5e-7
+ lua = 3.260216e-16
+ lub = -4.12618e-25
+ luc = -2.7409531e-17
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ pketa = 1.4501565e-15
+ pa0 = 1.1848049e-14
+ nlx = 0.0
+ pk1 = 7.144098e-15
+ pk2 = -4.137203e-15
+ pu0 = -1.1138246e-15
+ wpclm = 3.172275e-8
+ wub1 = 4.843047e-25
+ prt = 0
+ wuc1 = 2.7297169e-17
+ pua = -1.3255767e-22
+ pub = 5.546348e-32
+ puc = -6.669366e-24
+ tcjswg = 0.000645489
+ hdif = 2e-7
+ tcjsw = 0.000645489
+ rsh = 6.8
+ lub1 = 4.951269e-25
+ luc1 = 6.070172e-17
+ tcj = 0.001040287
+ ua1 = 1.224e-9
+ ub1 = -1.6810433e-18
+ uc1 = -8.806652e-11
+ wute = 1.8614003e-7
+ mjsw = 0.2003879
+ pvoff = 2.8052535e-15
+ tpb = 0.001554306
+ tox = 4.08e-9
+ wa0 = -9.831444e-9
+ lute = 2.2508574e-7
+ ute = -1.8126432
+ wk1 = -3.80072e-8
+ wk2 = 1.0172209e-8
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 1.0000000000000001e-20
+ wln = 1.0
+ wu0 = 3.280407e-9
+ wua = 2.9360883e-16
+ pvsat = 4.380818e-12
+ wub = -2.4531215e-25
+ wuc = -1.542897e-17
+ wwl = 0.0
+ wwn = 1
+ cdsc = 0.0
+ wketa = -1.5510503e-9
+ pvth0 = -5.378882e-16
+ xti = 3
+ drout = 0.0
+ cgdo = 3.665e-10
+ tpbsw = 0.001554306
+ cgso = 3.665e-10
+ cjswg = 3.340547e-10
+ nfactor = 1.0
+ mjswg = 0.43879
+ pnfactor = 0.0
+ cjsw = 2.040547e-10
+ wnfactor = 0.0
+ wvoff = -7.288315e-9
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ weta0 = 0
+ pscbe1 = 400000100.0
+ pscbe2 = 1e-6
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0011219129
+ pdiblcb = 0.01
+ wvsat = 0.0009435224
+ ppdiblc2 = 1.2928064e-16
+ tnom = 25.0
+ lpclm = 9.659676e-8
+ wvth0 = -9.251178e-9
+ wpdiblc2 = -1.1144895e-10
+ lnfactor = 0.0
+ nqsmod = 0
+ tpbswg = 0.001554306
+ toxm = 4.08e-9
+ noimod = 2
+ pcit = -2.4980728e-19
+ binunit = 2
+ pbsw = 0.6882682
+ pclm = 0.9444105
+ lpdiblc2 = 2.1785818e-9
+ lketa = -2.9090079e-9
+ xpart = 1
+ pkt1 = -5.199821e-15
+ pkt2 = -1.5611203e-15
+ keta = -0.017824383
+ pbswg = 0.6882682
+ dsub = 0.0
+ capmod = 3
+ version = 3.24
+ )

.model nch_mc_12 nmos (
+ level = 49
+ tpb = 0.001554306
+ tox = 4.08e-9
+ wa0 = 1.7605426e-7
+ pketa = -7.367843e-16
+ cjsw = 2.040547e-10
+ nfactor = 1.0
+ ute = -1.2073984
+ wk1 = -1.7855582e-8
+ wk2 = 1.6966123e-9
+ tcjswg = 0.000645489
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ wln = 1.0
+ wu0 = -4.268465e-11
+ wpclm = 1.9327061e-7
+ wua = -1.9101984e-17
+ wub = -5.11281e-26
+ wuc = -9.012729e-18
+ wwl = 0.0
+ wwn = 1
+ xti = 3
+ tcjsw = 0.000645489
+ tnom = 25.0
+ pdiblc1 = 1e-6
+ pdiblc2 = -0.00401322
+ pags = 1.8981756e-15
+ pdiblcb = 0.01
+ pvoff = -2.2207474e-15
+ toxm = 4.08e-9
+ pcit = -1.4232223e-17
+ pbsw = 0.6882682
+ pclm = 0.9948969
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = -1.1361991e-17
+ petab = 1.3954016e-17
+ binunit = 2
+ pvsat = 1.606088e-11
+ wketa = 3.203169e-9
+ pvth0 = 2.716016e-15
+ drout = 0.0
+ tpbsw = 0.001554306
+ a0 = 0.5005398
+ a1 = 0.0
+ a2 = 0.99
+ b0 = 0.0
+ b1 = 0.0
+ at = 20000.0
+ cf = 0
+ cj = 0.001000266
+ ef = 0.874
+ k1 = 0.489967
+ k2 = 0.029298484
+ k3 = 0.0
+ em = 30000000.0
+ js = 3.5e-7
+ cjswg = 3.340547e-10
+ ll = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ u0 = 0.03980552
+ pb = 0.6882682
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ua = -5.274002e-10
+ ub = 2.0039751e-18
+ uc = 7.914647e-11
+ mjswg = 0.43879
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ pkt1 = 2.3961372e-15
+ pkt2 = 8.832021e-16
+ keta = -0.027587207
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ wvoff = 3.637774e-9
+ wags = -4.12647e-9
+ dsub = 0.0
+ pscbe1 = 400000000.0
+ pscbe2 = 1e-6
+ weta0 = 2.4721704e-11
+ lags = -9.594464e-9
+ wetab = -3.0334849e-11
+ wcit = 3.093965e-11
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ wvsat = 0.000918131
+ version = 3.24
+ nqsmod = 0
+ lpclm = 7.337301e-8
+ wvth0 = -1.6324883e-8
+ tpbswg = 0.001554306
+ noimod = 2
+ lcit = 1.2733804e-10
+ voff = -0.1264125
+ ldif = 9e-8
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ pub1 = 1.6165291e-31
+ puc1 = 2.0250814e-23
+ eta0 = -0.00031223928
+ pvag = 0.0
+ etab = 0.0014101875
+ vsat = 84736.3
+ wint = 3e-9
+ pute = 4.383575e-14
+ vth0 = 0.4891579
+ rdsw = 170.0
+ wkt1 = -4.614678e-9
+ wkt2 = -3.214946e-9
+ lint = 1e-8
+ wmax = 1.2e-6
+ ags = 0.04085753
+ lketa = 1.5818911e-9
+ wmin = 5e-7
+ lkt1 = 1.6202869e-9
+ lkt2 = -8.228257e-11
+ lmax = 5e-7
+ xpart = 1
+ cit = 0.00022317801
+ lmin = 1.8e-7
+ pnfactor = 0.0
+ dlc = 3e-9
+ wnfactor = 0.0
+ k3b = 0.0
+ capmod = 3
+ dwb = 0.0
+ dwg = 0.0
+ pbswg = 0.6882682
+ lvoff = -4.057695e-10
+ wub1 = -1.1442477e-24
+ wuc1 = -9.658459e-17
+ ppdiblc2 = 3.905237e-16
+ hdif = 2e-7
+ beta0 = 11.59263
+ wpdiblc2 = -6.793707e-10
+ lub1 = -6.558089e-26
+ leta0 = 1.8963806e-10
+ luc1 = -7.416688e-18
+ wute = -3.505318e-7
+ mobmod = 1
+ la0 = 8.302936e-8
+ letab = -6.946862e-10
+ lnfactor = 0.0
+ mjsw = 0.2003879
+ lvsat = -0.00021356932
+ jsw = 1.45e-12
+ lk1 = 4.606408e-8
+ kt1 = -0.2249505
+ lk2 = -1.9413593e-8
+ kt2 = -0.028312566
+ lvth0 = 6.875945e-9
+ llc = -0.039
+ lln = -1
+ lute = -5.332685e-8
+ lu0 = 7.269945e-10
+ lua = -4.471944e-17
+ lub = 3.1333025e-26
+ luc = 1.0520902e-17
+ ppclm = -1.2237712e-15
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ delta = 0.01
+ pa0 = -7.365936e-14
+ nlx = 0.0
+ lpdiblc2 = 4.540744e-9
+ cdsc = 0.0
+ pk1 = -2.1256446e-15
+ pk2 = -2.3842633e-16
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ pu0 = 4.147977e-16
+ cgdo = 3.665e-10
+ prt = 0
+ pua = 1.1289303e-23
+ pub = -3.386118e-32
+ puc = -9.620837e-24
+ cgso = 3.665e-10
+ rsh = 6.8
+ tcj = 0.001040287
+ ua1 = 1.224e-9
+ ub1 = -4.621132e-19
+ uc1 = 6.001696e-11
+ )

.model nch_mc_13 nmos (
+ level = 49
+ drout = 0.0
+ wkt1 = 5.128653e-9
+ wkt2 = 3.532295e-9
+ tpbsw = 0.001554306
+ lint = 1e-8
+ wmax = 5e-7
+ wmin = 2.2e-7
+ cjswg = 3.340547e-10
+ lmax = 2.0001e-5
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ mjswg = 0.43879
+ lmin = 1e-5
+ pscbe1 = 200000030.0
+ pscbe2 = 1e-6
+ wvoff = -1.7276782e-9
+ weta0 = 0
+ nqsmod = 0
+ wub1 = -4.432931e-26
+ wuc1 = -1.7086574e-17
+ tpbswg = 0.001554306
+ wvsat = 0.0
+ noimod = 2
+ hdif = 2e-7
+ wvth0 = -1.5455745e-8
+ ags = 0.02
+ wute = 2.5547985e-8
+ mjsw = 0.2003879
+ cit = -9.999998e-5
+ dlc = 3e-9
+ k3b = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ cdsc = 0.0
+ cgdo = 3.665e-10
+ cgso = 3.665e-10
+ xpart = 1
+ jsw = 1.45e-12
+ capmod = 3
+ kt1 = -0.238767
+ lk2 = 0.0
+ kt2 = -0.03620588
+ llc = -0.039
+ cjsw = 2.040547e-10
+ lln = -1
+ a0 = 0.352982
+ a1 = 0.0
+ a2 = 0.99
+ lu0 = 0.0
+ b0 = 0.0
+ b1 = 0.0
+ pbswg = 0.6882682
+ nch = 3.9e+17
+ at = 20000.0
+ cf = 0
+ cj = 0.001000266
+ lwl = 0.0
+ lwn = 1.0
+ ef = 0.874
+ k1 = 0.5220979
+ k2 = 0.016542569
+ k3 = 0.0
+ em = 30000000.0
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ nfactor = 1.0
+ js = 3.5e-7
+ ll = 0.0
+ nlx = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ lvoff = 0.0
+ u0 = 0.03533742
+ pb = 0.6882682
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ua = -5.860608e-10
+ ub = 1.7266676e-18
+ uc = 7.252202e-11
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ mobmod = 1
+ beta0 = 11.59263
+ pu0 = 0.0
+ tnom = 25.0
+ leta0 = 8e-15
+ prt = 0
+ toxm = 4.08e-9
+ rsh = 6.8
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0006999999
+ lvth0 = 0.0
+ tcj = 0.001040287
+ ua1 = 1.224e-9
+ ub1 = -1.4270478e-18
+ uc1 = -6.39873e-11
+ pdiblcb = 0.01
+ pbsw = 0.6882682
+ pclm = 0.7999999
+ tpb = 0.001554306
+ tox = 4.08e-9
+ delta = 0.01
+ wa0 = 5.286186e-8
+ ute = -1.5833832
+ wk1 = -1.4938487e-9
+ wk2 = -2.6871128e-9
+ dvt0w = 0.0
+ dvt1w = 0.0
+ wln = 1.0
+ dvt2w = 0.0
+ wu0 = 9.682726e-10
+ binunit = 2
+ wua = -1.5275344e-17
+ wub = 1.2900942e-25
+ wuc = 2.9959555e-18
+ wwl = 0.0
+ wwn = 1
+ xti = 3
+ pnfactor = 0.0
+ keta = 0.002064252
+ tcjswg = 0.000645489
+ wnfactor = 0.0
+ dsub = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ tcjsw = 0.000645489
+ lnfactor = 0.0
+ voff = -0.1374522
+ version = 3.24
+ pvoff = 0.0
+ ldif = 9e-8
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ eta0 = 5e-5
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 1.0000000000000001e-20
+ pvag = 0.0
+ etab = -5e-5
+ vsat = 89999.99
+ wint = 3e-9
+ vth0 = 0.4632908
+ wketa = -2.9874625e-10
+ pvth0 = 0.0
+ rdsw = 170.0
+ )

.model nch_mc_14 nmos (
+ level = 49
+ la0 = -2.4964379e-7
+ pcit = 1.5653096e-18
+ pbsw = 0.6882682
+ pclm = 0.7606163
+ jsw = 1.45e-12
+ lk1 = -6.331243e-8
+ kt1 = -0.2407974
+ lk2 = 2.0798732e-8
+ kt2 = -0.03589625
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0003968183
+ pdiblcb = 0.01
+ lpscbe1 = 262.58182
+ llc = -0.039
+ lln = -1
+ lu0 = 9.894555e-9
+ lpdiblc2 = 3.0196909e-9
+ lua = -1.2876533e-16
+ lub = 7.836163e-25
+ luc = 7.064626e-17
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ pa0 = -7.427873e-14
+ nlx = 0.0
+ pk1 = 2.1894499e-14
+ pk2 = -1.0734859e-14
+ lketa = -3.0377027e-8
+ binunit = 2
+ pu0 = -1.3716021e-15
+ capmod = 3
+ prt = 0
+ pua = 1.6719826e-23
+ pub = -2.4068014e-31
+ xpart = 1
+ puc = -2.4186704e-23
+ pkt1 = -3.679308e-15
+ pkt2 = 5.879336e-16
+ rsh = 6.8
+ keta = 0.005114151
+ tcj = 0.001040287
+ ua1 = 1.224e-9
+ ub1 = -1.4513121e-18
+ uc1 = -6.991786e-11
+ pbswg = 0.6882682
+ tpb = 0.001554306
+ tox = 4.08e-9
+ dsub = 0.0
+ wa0 = 6.031956e-8
+ lvoff = -1.9727372e-8
+ mobmod = 1
+ ute = -1.5785241
+ wk1 = -3.692092e-9
+ wk2 = -1.6093152e-9
+ wcit = -1.5715551e-13
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ wln = 1.0
+ beta0 = 11.59263
+ wu0 = 1.1059835e-9
+ wua = -1.6954039e-17
+ wub = 1.5317406e-25
+ wuc = 5.42434e-18
+ leta0 = 8e-15
+ wwl = 0.0
+ wwn = 1
+ lcit = 2.6386249e-10
+ xti = 3
+ voff = -0.1354716
+ lvsat = -0.005267757
+ ldif = 9e-8
+ lvth0 = 5.627824e-8
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ pub1 = 2.1839324e-32
+ puc1 = 5.837128e-24
+ version = 3.24
+ ppclm = 7.826515e-14
+ eta0 = 5e-5
+ delta = 0.01
+ pvag = 0.0
+ etab = -5e-5
+ vsat = 90528.88
+ wint = 3e-9
+ pute = -1.7889165e-14
+ vth0 = 0.4576404
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ rdsw = 170.0
+ wkt1 = 5.498062e-9
+ wkt2 = 3.473265e-9
+ lint = 1e-8
+ wmax = 5e-7
+ wmin = 2.2e-7
+ lkt1 = 2.0222748e-8
+ lkt2 = -3.0839447e-9
+ lmax = 1e-5
+ tcjswg = 0.000645489
+ lmin = 1.2e-6
+ pketa = 4.776125e-16
+ wpclm = -7.857923e-9
+ wub1 = -4.652201e-26
+ wuc1 = -1.7672629e-17
+ tcjsw = 0.000645489
+ hdif = 2e-7
+ lub1 = 2.4167225e-25
+ a0 = 0.3780467
+ a1 = 0.0
+ a2 = 0.99
+ luc1 = 5.906839e-17
+ b0 = 0.0
+ b1 = 0.0
+ wute = 2.7344081e-8
+ mjsw = 0.2003879
+ at = 20000.0
+ pvoff = 2.7096929e-15
+ cf = 0
+ cj = 0.001000266
+ ef = 0.874
+ k1 = 0.5284545
+ k2 = 0.014454342
+ k3 = 0.0
+ em = 30000000.0
+ js = 3.5e-7
+ ll = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ u0 = 0.034344
+ pb = 0.6882682
+ w0 = 0.0
+ rd = 0
+ lute = -4.839696e-8
+ rs = 0
+ ua = -5.731325e-10
+ ub = 1.6479914e-18
+ uc = 6.542903e-11
+ cdscb = 0.0
+ cdscd = 0.0
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -2e-8
+ ww = 0.0
+ peta0 = 1.0000000000000001e-20
+ xw = 0.0
+ pvsat = 7.826533e-10
+ wketa = -3.466991e-10
+ pvth0 = -2.3944025e-15
+ cdsc = 0.0
+ drout = 0.0
+ tpbsw = 0.001554306
+ cgdo = 3.665e-10
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ cgso = 3.665e-10
+ cjswg = 3.340547e-10
+ pscbe1 = 173636400.0
+ pscbe2 = 1e-6
+ mjswg = 0.43879
+ ags = 0.02
+ pnfactor = 0.0
+ wnfactor = 0.0
+ wvoff = -1.9997353e-9
+ cjsw = 2.040547e-10
+ cit = -0.00012649217
+ nqsmod = 0
+ dlc = 3e-9
+ tpbswg = 0.001554306
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ noimod = 2
+ k3b = 0.0
+ weta0 = 0
+ dwb = 0.0
+ dwg = 0.0
+ wvsat = -7.857954e-5
+ nfactor = 1.0
+ lpclm = 3.92261e-7
+ wvth0 = -1.5215344e-8
+ tnom = 25.0
+ lnfactor = 0.0
+ toxm = 4.08e-9
+ )

.model nch_mc_15 nmos (
+ level = 49
+ wub1 = -1.0574451e-25
+ wuc1 = -4.040928e-17
+ ppdiblc2 = 4.703685e-16
+ beta0 = 11.59263
+ hdif = 2e-7
+ wpdiblc2 = -4.054901e-10
+ leta0 = 3.812228e-11
+ lub1 = -8.773805e-25
+ luc1 = -7.886598e-17
+ letab = -3.811428e-11
+ lnfactor = 0.0
+ wute = 1.9757099e-8
+ lvsat = -0.0007893788
+ mjsw = 0.2003879
+ lvth0 = 8.859259e-9
+ lute = -1.6751561e-7
+ ppclm = 4.863229e-14
+ delta = 0.01
+ lpdiblc2 = 1.4881204e-9
+ dvt0w = 0.0
+ cdsc = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ cgdo = 3.665e-10
+ tcjswg = 0.000645489
+ cgso = 3.665e-10
+ pketa = 3.1429577e-15
+ cjsw = 2.040547e-10
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ wpclm = 1.7687656e-8
+ tcjsw = 0.000645489
+ tnom = 25.0
+ nfactor = 1.0
+ pvoff = -1.3837542e-15
+ toxm = 4.08e-9
+ ags = 0.02
+ pcit = -9.088336e-19
+ pbsw = 0.6882682
+ pclm = 0.9728217
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 1.0000000000000001e-20
+ pvsat = 1.5955267e-11
+ cit = -0.00016124053
+ wketa = -2.6444102e-9
+ pvth0 = 7.985465e-17
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0017171376
+ dlc = 3e-9
+ drout = 0.0
+ pdiblcb = 0.01
+ k3b = 0.0
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ tpbsw = 0.001554306
+ dwb = 0.0
+ dwg = 0.0
+ pscbe1 = 400000100.0
+ pscbe2 = 1e-6
+ cjswg = 3.340547e-10
+ mjswg = 0.43879
+ binunit = 2
+ pkt1 = -1.1651986e-14
+ pkt2 = -1.4582807e-15
+ keta = -0.015611105
+ nqsmod = 0
+ wvoff = 1.529098e-9
+ tpbswg = 0.001554306
+ la0 = 2.7901473e-7
+ noimod = 2
+ jsw = 1.45e-12
+ dsub = 0.0
+ lk1 = 6.936774e-8
+ kt1 = -0.2426658
+ lk2 = -3.1528607e-8
+ kt2 = -0.04069558
+ llc = -0.039
+ lln = -1
+ weta0 = 0
+ lu0 = -1.7446106e-9
+ lua = 6.135559e-17
+ lub = -2.9489129e-25
+ luc = -2.7169401e-17
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ wvsat = 0.0005823669
+ wcit = 1.975718e-12
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ pa0 = 7.227613e-14
+ nlx = 0.0
+ lpclm = 1.4610272e-7
+ wvth0 = -1.7348324e-8
+ pk1 = -1.920543e-14
+ pk2 = 7.699883e-15
+ lcit = 3.0417063e-10
+ voff = -0.1694116
+ pu0 = 1.0146696e-15
+ ldif = 9e-8
+ prt = 0
+ pua = -1.8126578e-24
+ pub = -2.6935e-33
+ puc = -6.78799e-24
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ pub1 = 9.053745e-32
+ puc1 = 3.221165e-23
+ eta0 = 1.7142866e-5
+ rsh = 6.8
+ pvag = 0.0
+ etab = -1.7142866e-5
+ tcj = 0.001040287
+ ua1 = 1.224e-9
+ ub1 = -4.866116e-19
+ uc1 = 4.899104e-11
+ vsat = 86668.21
+ version = 3.24
+ a0 = -0.07769345
+ wint = 3e-9
+ a1 = 0.0
+ a2 = 0.99
+ pute = -9.088265e-15
+ b0 = 0.0
+ b1 = 0.0
+ tpb = 0.001554306
+ vth0 = 0.4985188
+ tox = 4.08e-9
+ at = 20000.0
+ cf = 0
+ cj = 0.001000266
+ ef = 0.874
+ k1 = 0.4140751
+ k2 = 0.05956412
+ k3 = 0.0
+ rdsw = 170.0
+ wa0 = -6.602082e-8
+ em = 30000000.0
+ js = 3.5e-7
+ wkt1 = 1.2371058e-8
+ wkt2 = 5.237243e-9
+ ute = -1.4758356
+ ll = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ lint = 1e-8
+ u0 = 0.04437776
+ pb = 0.6882682
+ wk1 = 3.173889e-8
+ wk2 = -1.7501334e-8
+ w0 = 0.0
+ rd = 0
+ wmax = 5e-7
+ lketa = -6.33573e-9
+ capmod = 3
+ rs = 0
+ ua = -7.370299e-10
+ ub = 2.5777392e-18
+ uc = 1.4975288e-10
+ wln = 1.0
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ xl = -2e-8
+ ww = 0.0
+ wmin = 2.2e-7
+ wu0 = -9.511471e-10
+ xw = 0.0
+ lkt1 = 2.2390124e-8
+ wua = -9.777621e-19
+ lkt2 = 2.4832894e-9
+ wub = -5.19868e-26
+ wuc = -9.57455e-18
+ xpart = 1
+ wwl = 0.0
+ wwn = 1
+ lmax = 1.2e-6
+ xti = 3
+ lmin = 5e-7
+ pnfactor = 0.0
+ wnfactor = 0.0
+ pbswg = 0.6882682
+ mobmod = 1
+ lvoff = 1.9643004e-8
+ )

.model nch_mc_16 nmos (
+ level = 49
+ at = 20000.0
+ cf = 0
+ cj = 0.001000266
+ ef = 0.874
+ k1 = 0.4942783
+ k2 = 0.023518253
+ k3 = 0.0
+ em = 30000000.0
+ pketa = -1.9609824e-16
+ pkt1 = 3.435378e-15
+ pkt2 = -8.505888e-17
+ wnfactor = 0.0
+ keta = -0.030443965
+ js = 3.5e-7
+ ll = 0.0
+ mj = 0.3595262
+ lw = 0.0
+ ags = 0.0548038
+ u0 = 0.0371035
+ pb = 0.6882682
+ w0 = 0.0
+ binunit = 2
+ rd = 0
+ rs = 0
+ ua = -6.614348e-10
+ ub = 2.1301375e-18
+ uc = 1.2526492e-10
+ wl = 0.0
+ wr = 1.0
+ xj = 1.6e-7
+ wags = -1.1015922e-8
+ xl = -2e-8
+ ww = 0.0
+ dsub = 0.0
+ xw = 0.0
+ wpclm = 1.2379924e-7
+ cit = 0.00029138371
+ lags = -1.6009743e-8
+ dlc = 3e-9
+ wcit = -2.7539906e-12
+ ppdiblc2 = -1.1422951e-16
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ tcjsw = 0.000645489
+ k3b = 0.0
+ wpdiblc2 = 8.65375e-10
+ dwb = 0.0
+ dwg = 0.0
+ lnfactor = 0.0
+ lcit = 9.596344e-11
+ pvoff = -4.969337e-16
+ voff = -0.1182414
+ ldif = 9e-8
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ pub1 = -3.181536e-32
+ puc1 = -1.1609298e-23
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 1.0000000000000001e-20
+ eta0 = -0.00026219533
+ pvag = 0.0
+ etab = 0.0013487812
+ pvsat = 1.2452966e-11
+ la0 = 1.1871046e-7
+ vsat = 85400.58
+ alpha0 = 0.0
+ alpha1 = 0.448150714
+ wint = 3e-9
+ pute = -6.731688e-15
+ wketa = 4.614407e-9
+ lpdiblc2 = 5.562512e-9
+ pvth0 = -1.0421574e-15
+ jsw = 1.45e-12
+ vth0 = 0.486292
+ lk1 = 3.247429e-8
+ kt1 = -0.1929406
+ lk2 = -1.4947512e-8
+ kt2 = -0.03937921
+ drout = 0.0
+ rdsw = 170.0
+ llc = -0.039
+ lln = -1
+ tpbsw = 0.001554306
+ pscbe1 = 400000000.0
+ pscbe2 = 1e-6
+ lu0 = 1.6015452e-9
+ version = 3.24
+ wkt1 = -2.0427562e-8
+ wkt2 = 2.2519782e-9
+ lint = 1e-8
+ lua = 2.6581833e-17
+ lub = -8.899446e-26
+ luc = -1.5904941e-17
+ nch = 3.9e+17
+ wmax = 5e-7
+ lwl = 0.0
+ lwn = 1.0
+ wmin = 2.2e-7
+ pa0 = -9.128582e-14
+ nlx = 0.0
+ cjswg = 3.340547e-10
+ lkt1 = -4.834396e-10
+ lkt2 = 1.8777602e-9
+ mjswg = 0.43879
+ pk1 = 4.587708e-15
+ pk2 = -2.4446703e-15
+ lmax = 5e-7
+ nqsmod = 0
+ tpbswg = 0.001554306
+ lmin = 1.8e-7
+ noimod = 2
+ pu0 = -1.7230291e-17
+ prt = 0
+ pua = -2.3933522e-23
+ pub = 2.5580594e-32
+ puc = 3.433529e-24
+ wvoff = -3.98773e-10
+ rsh = 6.8
+ tcj = 0.001040287
+ ua1 = 1.224e-9
+ ub1 = -3.1027764e-18
+ uc1 = -2.4653823e-10
+ weta0 = 0
+ tpb = 0.001554306
+ wub1 = 1.602399e-25
+ wuc1 = 5.485366e-17
+ tox = 4.08e-9
+ wvsat = 0.0005899806
+ wa0 = 2.8954867e-7
+ hdif = 2e-7
+ lpclm = 7.125815e-8
+ wvth0 = -1.4909164e-8
+ ute = -1.9466008
+ wk1 = -1.9985334e-8
+ wk2 = 4.552045e-9
+ lub1 = 3.260553e-25
+ luc1 = 5.707747e-17
+ wute = 1.4634106e-8
+ wln = 1.0
+ mjsw = 0.2003879
+ wu0 = 1.2921135e-9
+ wua = 4.711108e-17
+ wub = -1.1345223e-25
+ wuc = -3.179524e-17
+ wwl = 0.0
+ wwn = 1
+ xti = 3
+ lute = 4.90364e-8
+ cdsc = 0.0
+ capmod = 3
+ cgdo = 3.665e-10
+ lketa = 4.87385e-10
+ cgso = 3.665e-10
+ xpart = 1
+ mobmod = 1
+ cjsw = 2.040547e-10
+ pbswg = 0.6882682
+ noia = 2e+19
+ noib = 12000.0
+ noic = 2.5e-13
+ lvoff = -3.895271e-9
+ beta0 = 11.59263
+ leta0 = 1.6661783999999998e-10
+ tnom = 25.0
+ letab = -6.664392e-10
+ lvsat = -0.00020626588
+ pags = 5.067323e-15
+ lvth0 = 1.4483583e-8
+ toxm = 4.08e-9
+ nfactor = 1.0
+ pcit = 1.266836e-18
+ ppclm = -1.7902992e-16
+ pbsw = 0.6882682
+ pclm = 1.1355271
+ delta = 0.01
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ tcjswg = 0.000645489
+ pdiblc1 = 1e-6
+ pdiblc2 = -0.007140237
+ pdiblcb = 0.01
+ a0 = 0.270794
+ a1 = 0.0
+ a2 = 0.99
+ b0 = 0.0
+ b1 = 0.0
+ pnfactor = 0.0
+ )

.model pch_ss_1 pmos (
+ level = 49
+ lvth0 = -3.9543e-9
+ cdsc = 0.0
+ binunit = 2
+ pnfactor = 0
+ cgdo = 3.116e-10
+ delta = 0.01
+ wnfactor = 0.0
+ cgso = 3.116e-10
+ dvt0w = 0.0
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ dvt1w = 0.0
+ dvt2w = 0.0
+ pscbe1 = 199999970.0
+ pscbe2 = 5e-7
+ cjsw = 2.60505e-10
+ ags = 0.02
+ lnfactor = -3.9543e-9
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ nqsmod = 0
+ tpbswg = 0.001572025
+ noimod = 2
+ cit = -0.0001
+ dlc = 2e-9
+ tnom = 25.0
+ version = 3.24
+ k3b = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ toxm = 4.08e-9
+ tcjsw = 0.0004130718
+ pbsw = 0.895226
+ pclm = 0.6000001
+ pvoff = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ jsw = 1.2e-12
+ peta0 = 1.8966694548261387e-25
+ kt1 = -0.2311294
+ lk2 = 1.18629e-9
+ kt2 = -0.02433992
+ llc = -0.039
+ lln = -1
+ lu0 = -7.9086e-11
+ nch = 3.9e+17
+ pvth0 = -1.18629e-15
+ lwl = 0.0
+ lwn = 1.0
+ drout = 0.0
+ nlx = 0.0
+ tpbsw = 0.001572025
+ capmod = 3
+ keta = 0.026632193
+ pu0 = 0.0
+ cjswg = 4.43205e-10
+ prt = 0
+ dsub = 0.0
+ mjswg = 0.3683619
+ rsh = 7.2
+ tcj = 0.0009739001
+ ua1 = 1.224e-9
+ ub1 = -1.3928839e-18
+ uc1 = -4.59467e-12
+ wvoff = 0.0
+ mobmod = 1
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ tpb = 0.001572025
+ tox = 4.13259219e-9
+ ute = -0.8288856
+ voff = -0.1275921
+ weta0 = 0
+ ldif = 9e-8
+ wvsat = 0.0
+ wln = 1.0
+ kt1l = 0.0
+ prwb = 0.0
+ wu0 = -1.97715e-11
+ prwg = 0.0
+ wvth0 = -1.18629e-9
+ wwl = 0.0
+ wwn = 1.0
+ eta0 = 5e-5
+ xti = 3
+ pvag = 0.0
+ etab = -5e-5
+ vsat = 149999.98
+ wint = 5e-9
+ vth0 = -0.46220690000000003
+ rdsw = 530.0
+ lint = 1.4999999e-8
+ wmax = 0.000900001
+ wmin = 1.000869946e-5
+ a0 = 1.0461572
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ lmax = 2.0001e-5
+ at = 10000.0
+ cf = 0
+ cj = 0.00117705
+ lmin = 9.994740781e-6
+ ef = 1.064
+ k1 = 0.5375325
+ k2 = 0.04056858
+ k3 = 0.0
+ em = 30000000.0
+ tcjswg = 0.0004130718
+ js = 2.5e-7
+ ll = 0.0
+ mj = 0.4476
+ lw = 0.0
+ u0 = 0.0108097578
+ pb = 0.895226
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ua = 8.23294e-10
+ ub = 6.854322e-19
+ uc = -8.655411e-11
+ wl = 0.0
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -1.4740781e-8
+ ww = 0.0
+ xw = -8.69946e-9
+ xpart = 1
+ nfactor = 1.0
+ pbswg = 0.895226
+ hdif = 2e-7
+ lvoff = -1.5817200000000002e-9
+ mjsw = 0.3683619
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0010000003
+ pdiblcb = 0.01
+ beta0 = 22.67827
+ leta0 = 1.8966694548261387e-18
+ )

.model pch_ss_2 pmos (
+ level = 49
+ mj = 0.4476
+ lw = 0.0
+ kt1 = -0.2295883
+ lk1 = 1.8783622e-8
+ kt2 = -0.024031118
+ lk2 = -4.300882e-9
+ u0 = 0.0109398048
+ pb = 0.895226
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ua = 8.625313e-10
+ ub = 6.401998e-19
+ uc = -8.855145e-11
+ llc = -0.039
+ lln = -1
+ wl = 0.0
+ lu0 = -1.3730549e-9
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -1.4740781e-8
+ ww = 0.0
+ xw = -8.69946e-9
+ voff = -0.1274002
+ lua = -3.904111e-16
+ lub = 4.500626e-25
+ luc = 1.9873557e-17
+ ldif = 9e-8
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ kt1l = 0.0
+ tcjsw = 0.0004130718
+ prwb = 0.0
+ prwg = 0.0
+ nlx = 0.0
+ eta0 = 5e-5
+ pvag = 0.0
+ etab = -5e-5
+ pvoff = 0.0
+ vsat = 151306.8
+ pu0 = 0.0
+ wint = 5e-9
+ prt = 0
+ vth0 = -0.45971300000000004
+ rdsw = 530.0
+ pnfactor = 0
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 1.8966694548261387e-25
+ lint = 1.4999999e-8
+ rsh = 7.2
+ tcj = 0.0009739001
+ ua1 = 1.224e-9
+ wnfactor = 0.0
+ wmax = 0.000900001
+ ub1 = -1.3977103e-18
+ uc1 = -6.694918e-12
+ wmin = 1.000869946e-5
+ tpb = 0.001572025
+ capmod = 3
+ pvth0 = -1.18629e-15
+ tox = 4.13259219e-9
+ lkt1 = -1.5333228e-8
+ lkt2 = -3.0725886e-9
+ drout = 0.0
+ lmax = 9.994740781e-6
+ tpbsw = 0.001572025
+ ute = -0.8385549
+ lmin = 1.194740781e-6
+ wln = 1.0
+ wu0 = -1.97715e-11
+ cjswg = 4.43205e-10
+ wwl = 0.0
+ wwn = 1.0
+ mjswg = 0.3683619
+ lnfactor = -3.9543e-9
+ xti = 3
+ mobmod = 1
+ nfactor = 1.0
+ wvoff = 0.0
+ hdif = 2e-7
+ lub1 = 4.802326e-26
+ luc1 = 2.0897466e-17
+ weta0 = 0
+ mjsw = 0.3683619
+ lpdiblc2 = 5.201137e-9
+ wvsat = 0.0
+ lute = 9.620972e-8
+ lpclm = 2.6005682e-7
+ wvth0 = -1.18629e-9
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0004772727
+ pdiblcb = 0.01
+ lpscbe1 = 195.04263
+ cdsc = 0.0
+ cgdo = 3.116e-10
+ binunit = 2
+ cgso = 3.116e-10
+ tcjswg = 0.0004130718
+ lketa = -2.0462676e-9
+ cjsw = 2.60505e-10
+ xpart = 1
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ pbswg = 0.895226
+ tnom = 25.0
+ lvoff = -3.4908509e-9
+ toxm = 4.08e-9
+ beta0 = 22.67827
+ version = 3.24
+ pbsw = 0.895226
+ pclm = 0.5738637
+ leta0 = 1.8966694548261387e-18
+ lvsat = -0.013002843
+ lvth0 = -2.8768353e-8
+ ags = 0.02
+ delta = 0.01
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ cit = -0.0001
+ dlc = 2e-9
+ dvt0w = 0.0
+ dvt1w = 0.0
+ pscbe1 = 180397680.0
+ pscbe2 = 5e-7
+ dvt2w = 0.0
+ k3b = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ keta = 0.026837848
+ nqsmod = 0
+ tpbswg = 0.001572025
+ dsub = 0.0
+ noimod = 2
+ a0 = 1.0385712
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ at = 10000.0
+ cf = 0
+ cj = 0.00117705
+ la0 = 7.548124e-8
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ ef = 1.064
+ k1 = 0.5356447
+ k2 = 0.041120050000000005
+ k3 = 0.0
+ em = 30000000.0
+ js = 2.5e-7
+ jsw = 1.2e-12
+ ll = 0.0
+ )

.model pch_ss_3 pmos (
+ level = 49
+ cjswg = 4.43205e-10
+ mjswg = 0.3683619
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ wvoff = 0.0
+ tnom = 25.0
+ weta0 = 0
+ wvsat = 0.0
+ toxm = 4.08e-9
+ a0 = 1.0045335
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ lpclm = 1.4785704e-7
+ wvth0 = -1.18629e-9
+ pbsw = 0.895226
+ pclm = 0.6714287
+ at = 10000.0
+ cf = 0
+ cj = 0.00117705
+ ef = 1.064
+ k1 = 0.5405614
+ k2 = 0.04043759
+ k3 = 0.0
+ em = 30000000.0
+ js = 2.5e-7
+ version = 3.24
+ ll = 0.0
+ mj = 0.4476
+ lw = 0.0
+ u0 = 0.0101692238
+ pb = 0.895226
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ua = 5.26694e-10
+ ub = 1.1734415e-18
+ uc = -4.332115e-11
+ wl = 0.0
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -1.4740781e-8
+ ww = 0.0
+ xw = -8.69946e-9
+ pnfactor = 0
+ wnfactor = 0.0
+ tcjswg = 0.0004130718
+ lketa = -8.158225e-9
+ keta = 0.03215259
+ xpart = 1
+ dsub = 0.0
+ lnfactor = -3.9543e-9
+ ags = 0.02
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ pbswg = 0.895226
+ lvoff = -2.5305025000000003e-9
+ lcit = 2.2402701e-10
+ cit = -0.00029480609
+ voff = -0.1282353
+ lpdiblc2 = 3.696428e-9
+ ldif = 9e-8
+ dlc = 2e-9
+ beta0 = 22.67827
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ k3b = 0.0
+ dwb = 0.0
+ leta0 = 3.6964281896669455e-11
+ dwg = 0.0
+ eta0 = 1.7857143e-5
+ letab = -3.696428e-11
+ pvag = 0.0
+ etab = -1.7857143e-5
+ lvsat = -0.007392833
+ vsat = 146428.53
+ wint = 5e-9
+ lvth0 = -1.0643742e-8
+ vth0 = -0.4754736
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ rdsw = 530.0
+ delta = 0.01
+ lint = 1.4999999e-8
+ wmax = 0.000900001
+ pscbe1 = 349999900.0
+ pscbe2 = 5e-7
+ la0 = 1.146246e-7
+ wmin = 1.000869946e-5
+ jsw = 1.2e-12
+ lkt1 = 1.5747348e-9
+ lkt2 = 9.740028e-10
+ kt1 = -0.2442909
+ lk1 = 1.3129389e-8
+ kt2 = -0.027549893
+ lk2 = -3.5160449999999997e-9
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ lmax = 1.194740781e-6
+ llc = -0.039
+ lln = -1
+ lu0 = -4.868866e-10
+ lmin = 4.94740781e-7
+ lua = -4.198125e-18
+ lub = -1.631654e-25
+ luc = -3.214129e-17
+ nch = 3.9e+17
+ nqsmod = 0
+ lwl = 0.0
+ lwn = 1.0
+ tpbswg = 0.001572025
+ noimod = 2
+ nlx = 0.0
+ pu0 = 0.0
+ prt = 0
+ hdif = 2e-7
+ rsh = 7.2
+ tcj = 0.0009739001
+ nfactor = 1.0
+ ua1 = 1.224e-9
+ lub1 = 3.0810812e-26
+ ub1 = -1.3827429e-18
+ luc1 = 2.9752128e-17
+ uc1 = -1.4394627e-11
+ mjsw = 0.3683619
+ tpb = 0.001572025
+ tox = 4.13259219e-9
+ tcjsw = 0.0004130718
+ lute = 3.654092e-8
+ ute = -0.786669
+ wln = 1.0
+ pvoff = 0.0
+ wu0 = -1.97715e-11
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0017857148
+ wwl = 0.0
+ wwn = 1.0
+ pdiblcb = 0.01
+ cdsc = 0.0
+ xti = 3
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 1.8966694548261387e-25
+ capmod = 3
+ cgdo = 3.116e-10
+ pvth0 = -1.18629e-15
+ cgso = 3.116e-10
+ drout = 0.0
+ binunit = 2
+ tpbsw = 0.001572025
+ cjsw = 2.60505e-10
+ mobmod = 1
+ )

.model pch_ss_4 pmos (
+ level = 49
+ wmin = 1.000869946e-5
+ lkt1 = -2.665e-9
+ lkt2 = -2.325577e-10
+ lmax = 4.94740781e-7
+ cit = -4.054396e-5
+ lmin = 1.8e-7
+ lketa = -8.307595e-10
+ dlc = 2e-9
+ k3b = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ xpart = 1
+ pbswg = 0.895226
+ hdif = 2e-7
+ lub1 = 2.883988e-26
+ luc1 = -6.846759e-18
+ lvoff = -1.6174359200000002e-9
+ la0 = 1.6196543e-8
+ mjsw = 0.3683619
+ jsw = 1.2e-12
+ kt1 = -0.2348693
+ lk1 = 1.6807924e-8
+ kt2 = -0.024868647
+ lk2 = -4.689925e-9
+ beta0 = 22.67827
+ nfactor = 1.0
+ llc = -0.039
+ lln = -1
+ lu0 = -1.7803381e-10
+ lute = 1.6013461e-9
+ leta0 = 2.559375218966695e-10
+ lua = -1.5999061e-16
+ lub = 1.2197973e-25
+ luc = 1.8500639e-17
+ nch = 3.9e+17
+ letab = -5.298917e-10
+ lwl = 0.0
+ lwn = 1.0
+ lvsat = -0.0003656265
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ nlx = 0.0
+ lvth0 = -1.2194852e-8
+ cdsc = 0.0
+ pscbe1 = 350000000.0
+ pscbe2 = 5e-7
+ pnfactor = 0
+ pu0 = 0.0
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.00796875
+ delta = 0.01
+ a0 = 1.2232625
+ a1 = 0.0
+ a2 = 0.4
+ prt = 0
+ b0 = 0.0
+ b1 = 0.0
+ cgdo = 3.116e-10
+ wnfactor = 0.0
+ pdiblcb = 0.01
+ at = 10000.0
+ cf = 0
+ cj = 0.00117705
+ ef = 1.064
+ k1 = 0.5323869
+ k2 = 0.04304621
+ k3 = 0.0
+ em = 30000000.0
+ cgso = 3.116e-10
+ js = 2.5e-7
+ dvt0w = 0.0
+ dvt1w = 0.0
+ ll = 0.0
+ rsh = 7.2
+ mj = 0.4476
+ dvt2w = 0.0
+ lw = 0.0
+ u0 = 0.0094828838
+ tcj = 0.0009739001
+ nqsmod = 0
+ pb = 0.895226
+ ua1 = 1.224e-9
+ w0 = 0.0
+ ub1 = -1.3783631e-18
+ rd = 0
+ uc1 = 6.693623e-11
+ tpbswg = 0.001572025
+ rs = 0
+ ua = 8.728995e-10
+ ub = 5.397856e-19
+ uc = -1.5585878e-10
+ noimod = 2
+ wl = 0.0
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -1.4740781e-8
+ ww = 0.0
+ xw = -8.69946e-9
+ tpb = 0.001572025
+ tox = 4.13259219e-9
+ binunit = 2
+ cjsw = 2.60505e-10
+ ute = -0.7090256
+ lnfactor = -3.9543e-9
+ wln = 1.0
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ wu0 = -1.97715e-11
+ wwl = 0.0
+ wwn = 1.0
+ xti = 3
+ tnom = 25.0
+ lcdscd = 3.65625e-11
+ lpdiblc2 = 9.140626e-10
+ toxm = 4.08e-9
+ tcjsw = 0.0004130718
+ pbsw = 0.895226
+ pclm = 0.9102259
+ pvoff = 0.0
+ capmod = 3
+ version = 3.24
+ cdscb = 0.0
+ cdscd = -8.125e-5
+ peta0 = 1.8966694548261387e-25
+ pvth0 = -1.18629e-15
+ drout = 0.0
+ tpbsw = 0.001572025
+ mobmod = 1
+ keta = 0.015869336
+ cjswg = 4.43205e-10
+ mjswg = 0.3683619
+ dsub = 0.0
+ wvoff = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ weta0 = 0
+ lcit = 1.0960905e-10
+ voff = -0.1302643
+ ldif = 9e-8
+ wvsat = 0.0
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ lpclm = 4.03983e-8
+ wvth0 = -1.18629e-9
+ eta0 = -0.0004687502
+ pvag = 0.0
+ etab = 0.0010775371
+ vsat = 130812.52
+ wint = 5e-9
+ vth0 = -0.4720267
+ rdsw = 530.0
+ tcjswg = 0.0004130718
+ lint = 1.4999999e-8
+ wmax = 0.000900001
+ ags = 0.02
+ )

.model pch_ss_5 pmos (
+ level = 49
+ wa0 = -4.787191e-8
+ pscbe1 = 199999970.0
+ pscbe2 = 5e-7
+ ute = -0.8394966
+ lvth0 = -3.9543e-9
+ wk1 = 1.2456701e-8
+ wk2 = -5.940143e-9
+ wln = 1.0
+ wu0 = -1.2692462000000002e-9
+ delta = 0.01
+ wua = 1.7543858e-16
+ wub = -6.530953e-25
+ wuc = -7.950096e-17
+ wwl = 0.0
+ wwn = 1.0
+ nqsmod = 0
+ xti = 3
+ version = 3.24
+ tpbswg = 0.001572025
+ noimod = 2
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ keta = 0.02600144
+ dsub = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ voff = -0.1274889
+ ldif = 9e-8
+ tcjsw = 0.0004130718
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ eta0 = 5e-5
+ pvoff = 0.0
+ capmod = 3
+ pvag = 0.0
+ etab = -5e-5
+ vsat = 149999.98
+ wint = 5e-9
+ vth0 = -0.4634952
+ cdscb = 0.0
+ rdsw = 530.0
+ cdscd = 0.0
+ pnfactor = 0
+ peta0 = 1.8966694548261387e-25
+ wkt1 = 8.228274e-9
+ wkt2 = 1.4868883e-9
+ lint = 1.4999999e-8
+ wnfactor = 0.0
+ wmax = 1.000869946e-5
+ wketa = 6.301227e-9
+ wmin = 1.20869946e-6
+ pvth0 = -1.18629e-15
+ mobmod = 1
+ drout = 0.0
+ tpbsw = 0.001572025
+ lmax = 2.0001e-5
+ lmin = 9.994740781e-6
+ cjswg = 4.43205e-10
+ a0 = 1.0509492
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ at = 10000.0
+ mjswg = 0.3683619
+ cf = 0
+ cj = 0.00117705
+ lnfactor = -3.9543e-9
+ ef = 1.064
+ k1 = 0.5362856
+ k2 = 0.04116319
+ k3 = 0.0
+ em = 30000000.0
+ js = 2.5e-7
+ ll = 0.0
+ mj = 0.4476
+ lw = 0.0
+ u0 = 0.0109348308
+ pb = 0.895226
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ wvoff = -1.0305298e-9
+ ua = 8.057326e-10
+ ub = 7.508071e-19
+ uc = -7.859605e-11
+ wub1 = 6.909715e-26
+ wuc1 = 3.0354498e-17
+ wl = 0.0
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -1.4740781e-8
+ ww = 0.0
+ xw = -8.69946e-9
+ hdif = 2e-7
+ weta0 = 0
+ ags = 0.02
+ wute = 1.0600407e-7
+ mjsw = 0.3683619
+ wvsat = 0.0
+ wvth0 = 1.1684168e-8
+ cit = -0.0001
+ dlc = 2e-9
+ nfactor = 1.0
+ k3b = 0.0
+ tcjswg = 0.0004130718
+ dwb = 0.0
+ dwg = 0.0
+ cdsc = 0.0
+ cgdo = 3.116e-10
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0010000004
+ cgso = 3.116e-10
+ pdiblcb = 0.01
+ jsw = 1.2e-12
+ kt1 = -0.231953
+ kt2 = -0.024488758
+ lk2 = 1.18629e-9
+ llc = -0.039
+ lln = -1
+ cjsw = 2.60505e-10
+ lu0 = -7.9086e-11
+ xpart = 1
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ binunit = 2
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ nlx = 0.0
+ pbswg = 0.895226
+ pu0 = 0.0
+ prt = 0
+ tnom = 25.0
+ lvoff = -1.5817200000000002e-9
+ rsh = 7.2
+ beta0 = 22.67827
+ toxm = 4.08e-9
+ tcj = 0.0009739001
+ ua1 = 1.224e-9
+ ub1 = -1.3998005e-18
+ uc1 = -7.633158e-12
+ leta0 = 1.8966694548261387e-18
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ pbsw = 0.895226
+ pclm = 0.6000001
+ tpb = 0.001572025
+ tox = 4.13259219e-9
+ )

.model pch_ss_6 pmos (
+ level = 49
+ lub1 = 5.442727e-26
+ luc1 = 1.8276951e-17
+ wute = 1.0644106e-7
+ mjsw = 0.3683619
+ tcjsw = 0.0004130718
+ capmod = 3
+ lute = 9.664497e-8
+ pvoff = -4.403278e-15
+ nfactor = 1.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 1.8966694548261387e-25
+ mobmod = 1
+ cgdo = 3.116e-10
+ wketa = 7.084359e-9
+ pvth0 = -6.522762e-15
+ cgso = 3.116e-10
+ drout = 0.0
+ tpbsw = 0.001572025
+ ags = 0.02
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0004772728
+ pdiblcb = 0.01
+ lpscbe1 = 195.04262
+ cjswg = 4.43205e-10
+ cit = -0.0001
+ cjsw = 2.60505e-10
+ mjswg = 0.3683619
+ dlc = 2e-9
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ k3b = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ wvoff = -5.879894e-10
+ binunit = 2
+ tnom = 25.0
+ weta0 = 0
+ wvsat = 0.0
+ toxm = 4.08e-9
+ lpclm = 2.6005682e-7
+ wvth0 = 1.2220496e-8
+ la0 = 6.878132e-8
+ pbsw = 0.895226
+ tcjswg = 0.0004130718
+ pclm = 0.5738637
+ jsw = 1.2e-12
+ kt1 = -0.2303147
+ lk1 = 1.8184398e-8
+ kt2 = -0.024155809
+ lk2 = -4.094344999999999e-9
+ llc = -0.039
+ lln = -1
+ lu0 = -1.3846097e-9
+ lua = -3.935608e-16
+ lub = 4.219459e-25
+ luc = 1.8883157e-17
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ pnfactor = 0
+ pa0 = 6.693222e-14
+ nlx = 0.0
+ wnfactor = 0.0
+ pk1 = 5.986243e-15
+ pk2 = -2.063307e-15
+ pu0 = 1.1543239e-16
+ prt = 0
+ pua = 3.1465633e-23
+ pub = 2.8088595e-31
+ puc = 9.8941e-24
+ version = 3.24
+ lketa = -1.2662711e-9
+ rsh = 7.2
+ pkt1 = 9.666697e-15
+ tcj = 0.0009739001
+ pkt2 = 2.4000725e-15
+ ua1 = 1.224e-9
+ keta = 0.026128704
+ ub1 = -1.4052706e-18
+ uc1 = -9.470036e-12
+ xpart = 1
+ tpb = 0.001572025
+ lnfactor = -3.9543e-9
+ tox = 4.13259219e-9
+ dsub = 0.0
+ wa0 = -5.459876e-8
+ ute = -0.8492097
+ wk1 = 1.185507e-8
+ wk2 = -5.732776e-9
+ pbswg = 0.895226
+ wln = 1.0
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ wu0 = -1.2808475e-9
+ wua = 1.7227619e-16
+ wub = -6.81325e-25
+ wuc = -8.049533e-17
+ wwl = 0.0
+ wwn = 1.0
+ a0 = 1.0440365
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ lvoff = -3.0500824000000002e-9
+ xti = 3
+ at = 10000.0
+ cf = 0
+ lpdiblc2 = 5.201137e-9
+ cj = 0.00117705
+ voff = -0.1273414
+ ef = 1.064
+ k1 = 0.534458
+ k2 = 0.04169391
+ k3 = 0.0
+ em = 30000000.0
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ ldif = 9e-8
+ beta0 = 22.67827
+ js = 2.5e-7
+ ll = 0.0
+ mj = 0.4476
+ lw = 0.0
+ u0 = 0.0110660398
+ pb = 0.895226
+ kt1l = 0.0
+ w0 = 0.0
+ prwb = 0.0
+ rd = 0
+ pub1 = -6.397619e-32
+ prwg = 0.0
+ leta0 = 1.8966694548261387e-18
+ puc1 = 2.6178952e-23
+ rs = 0
+ ua = 8.452865e-10
+ ub = 7.084005e-19
+ uc = -8.049386e-11
+ pscbe1 = 180397700.0
+ pscbe2 = 5e-7
+ wl = 0.0
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -1.4740781e-8
+ ww = 0.0
+ xw = -8.69946e-9
+ eta0 = 5e-5
+ lvsat = -0.013002842
+ pvag = 0.0
+ etab = -5e-5
+ vsat = 151306.8
+ lvth0 = -2.8234169e-8
+ wint = 5e-9
+ pute = -4.348101e-15
+ vth0 = -0.4610551
+ nqsmod = 0
+ rdsw = 530.0
+ tpbswg = 0.001572025
+ delta = 0.01
+ wkt1 = 7.256747e-9
+ wkt2 = 1.245675e-9
+ noimod = 2
+ lint = 1.4999999e-8
+ wmax = 1.000869946e-5
+ wmin = 1.20869946e-6
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ lkt1 = -1.6300865e-8
+ lkt2 = -3.312836e-9
+ lmax = 9.994740781e-6
+ lmin = 1.194740781e-6
+ pketa = -7.792167e-15
+ wub1 = 7.552692e-26
+ wuc1 = 2.7723443e-17
+ hdif = 2e-7
+ )

.model pch_ss_7 pmos (
+ level = 49
+ mjswg = 0.3683619
+ jsw = 1.2e-12
+ kt1 = -0.2459144
+ lk1 = 8.371453e-9
+ kt2 = -0.027846618
+ lk2 = -2.029564e-9
+ dsub = 0.0
+ llc = -0.039
+ lln = -1
+ lu0 = -4.248086e-10
+ wvoff = -7.866491e-9
+ lua = 3.0792715e-17
+ lub = -1.9665828e-25
+ luc = -3.700045e-17
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ wcit = -1.788104e-11
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ pa0 = -1.2519753e-13
+ nlx = 0.0
+ weta0 = 0
+ pk1 = 4.753178e-14
+ pk2 = -1.4849934e-14
+ lcit = 2.2196864e-10
+ voff = -0.1274479
+ pu0 = -6.201592e-16
+ wvsat = 0.0
+ ldif = 9e-8
+ tcjswg = 0.0004130718
+ prt = 0
+ pua = -3.495584e-22
+ pub = 3.345938e-31
+ puc = 4.854297e-23
+ lpclm = 1.4785702e-7
+ wvth0 = 8.94442e-9
+ kt1l = 0.0
+ prwb = 0.0
+ pub1 = -1.382964e-31
+ prwg = 0.0
+ puc1 = -5.043768e-23
+ eta0 = 1.7857139e-5
+ rsh = 7.2
+ tcj = 0.0009739001
+ ua1 = 1.224e-9
+ pvag = 0.0
+ ub1 = -1.3967723e-18
+ etab = -1.7857139e-5
+ uc1 = -2.3838735e-11
+ vsat = 146428.53
+ wint = 5e-9
+ pute = 2.0900147e-14
+ tpb = 0.001572025
+ tox = 4.13259219e-9
+ vth0 = -0.4764877
+ wa0 = 1.1247056e-7
+ rdsw = 530.0
+ ute = -0.7951261
+ wkt1 = 1.6218328e-8
+ wkt2 = 2.9642964e-9
+ wk1 = -2.4271484e-8
+ wk2 = 5.386031e-9
+ lint = 1.4999999e-8
+ wmax = 1.000869946e-5
+ wln = 1.0
+ wu0 = -6.412026e-10
+ wmin = 1.20869946e-6
+ wua = 5.036014e-16
+ wub = -7.280275e-25
+ wuc = -1.1410304e-16
+ lkt1 = 1.6387112e-9
+ lkt2 = 9.315946e-10
+ wwl = 0.0
+ wwn = 1.0
+ xti = 3
+ lmax = 1.194740781e-6
+ lketa = -8.380984e-9
+ lmin = 4.94740781e-7
+ xpart = 1
+ wub1 = 1.4015321e-25
+ pbswg = 0.895226
+ wuc1 = 9.434661e-17
+ hdif = 2e-7
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ lvoff = -2.9275995000000004e-9
+ lub1 = 4.46543e-26
+ luc1 = 3.480094e-17
+ wute = 8.448607e-8
+ mjsw = 0.3683619
+ pscbe1 = 349999900.0
+ pscbe2 = 5e-7
+ beta0 = 22.67827
+ leta0 = 3.6964291896669454e-11
+ lute = 3.444881e-8
+ letab = -3.696429e-11
+ lvsat = -0.007392833
+ lvth0 = -1.0486687e-8
+ nqsmod = 0
+ tpbswg = 0.001572025
+ noimod = 2
+ cdsc = 0.0
+ pnfactor = 0
+ delta = 0.01
+ wnfactor = 0.0
+ cgdo = 3.116e-10
+ nfactor = 1.0
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ cgso = 3.116e-10
+ cjsw = 2.60505e-10
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0017857144
+ lnfactor = -3.9543e-9
+ pdiblcb = 0.01
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ pketa = 2.2253538e-15
+ tnom = 25.0
+ binunit = 2
+ capmod = 3
+ lpdiblc2 = 3.696428e-9
+ tcjsw = 0.0004130718
+ toxm = 4.08e-9
+ ags = 0.02
+ pcit = 2.0563189e-17
+ pbsw = 0.895226
+ pclm = 0.6714287
+ pvoff = 3.966999e-15
+ cit = -0.0002930162
+ a0 = 0.9932752
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ at = 10000.0
+ mobmod = 1
+ cf = 0
+ dlc = 2e-9
+ cj = 0.00117705
+ ef = 1.064
+ k1 = 0.542991
+ k2 = 0.03989844
+ k3 = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ em = 30000000.0
+ peta0 = 1.8966694548261387e-25
+ k3b = 0.0
+ js = 2.5e-7
+ ll = 0.0
+ mj = 0.4476
+ lw = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ u0 = 0.0102314288
+ pb = 0.895226
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ua = 4.762835e-10
+ ub = 1.2463172e-18
+ uc = -3.189942e-11
+ wl = 0.0
+ wr = 1.0
+ xj = 1.7000001e-7
+ wketa = -1.6265284e-9
+ xl = -1.4740781e-8
+ ww = 0.0
+ xw = -8.69946e-9
+ pvth0 = -2.7552727999999998e-15
+ drout = 0.0
+ tpbsw = 0.001572025
+ pkt1 = -6.391237e-16
+ pkt2 = 4.236579e-16
+ keta = 0.03231541
+ cjswg = 4.43205e-10
+ version = 3.24
+ la0 = 1.2715688e-7
+ )

.model pch_ss_8 pmos (
+ level = 49
+ cgso = 3.116e-10
+ nfactor = 1.0
+ a0 = 1.2640158
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ lketa = -5.872592e-10
+ at = 10000.0
+ cf = 0
+ cj = 0.00117705
+ ef = 1.064
+ k1 = 0.5203763
+ k2 = 0.04747528
+ k3 = 0.0
+ em = 30000000.0
+ pcdscd = -7.408954e-18
+ js = 2.5e-7
+ ll = 0.0
+ mj = 0.4476
+ lw = 0.0
+ u0 = 0.0097404008
+ pb = 0.895226
+ xpart = 1
+ w0 = 0.0
+ rd = 0
+ cjsw = 2.60505e-10
+ rs = 0
+ ua = 9.357863e-10
+ ub = 5.091257e-19
+ uc = -1.5731644e-10
+ wl = 0.0
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -1.4740781e-8
+ ww = 0.0
+ xw = -8.69946e-9
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.007987866
+ pbswg = 0.895226
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ pdiblcb = 0.01
+ pscbe1 = 350000000.0
+ pscbe2 = 5e-7
+ lvoff = -1.4181850500000001e-9
+ tnom = 25.0
+ pags = -6.875222e-16
+ beta0 = 22.67827
+ toxm = 4.08e-9
+ binunit = 2
+ leta0 = 2.559375218966695e-10
+ letab = -5.545772e-10
+ nqsmod = 0
+ pcit = -7.907631e-17
+ pbsw = 0.895226
+ pclm = 0.9107697
+ tpbswg = 0.001572025
+ lvsat = -0.0003656271
+ noimod = 2
+ lvth0 = -1.2082326e-8
+ ppclm = 2.4445072e-15
+ delta = 0.01
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ lcdscd = 3.730414e-11
+ pkt1 = -1.8229216e-15
+ pkt2 = -1.2254391e-15
+ keta = 0.014996022
+ ags = 0.019847063
+ wags = 1.5278273e-9
+ dsub = 0.0
+ version = 3.24
+ cit = -6.09184e-5
+ pketa = -2.4325694e-15
+ dlc = 2e-9
+ lags = 6.882101e-11
+ wcit = 2.0354016e-10
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ k3b = 0.0
+ capmod = 3
+ dwb = 0.0
+ dwg = 0.0
+ wpclm = -5.432238e-9
+ lcit = 1.1752459e-10
+ voff = -0.1308021
+ tcjsw = 0.0004130718
+ ldif = 9e-8
+ kt1l = 0.0
+ prwb = 0.0
+ pub1 = 2.7781507e-32
+ prwg = 0.0
+ puc1 = 8.113434e-24
+ pvoff = -1.9905158e-15
+ eta0 = -0.0004687502
+ mobmod = 1
+ pvag = 0.0
+ etab = 0.0011323938
+ la0 = 5.323636e-9
+ vsat = 130812.52
+ wint = 5e-9
+ pute = 9.798417e-15
+ jsw = 1.2e-12
+ kt1 = -0.2367561
+ lk1 = 1.854804e-8
+ kt2 = -0.025532207
+ lk2 = -5.439136e-9
+ vth0 = -0.4729418
+ cdscb = 0.0
+ cdscd = -8.289813e-5
+ pnfactor = 0
+ peta0 = 1.8966694548261387e-25
+ llc = -0.039
+ rdsw = 530.0
+ lln = -1
+ lu0 = -2.0384533e-10
+ petab = 2.4660761e-16
+ wnfactor = 0.0
+ wkt1 = 1.8848993e-8
+ wkt2 = 6.628956e-9
+ lua = -1.759835e-16
+ lub = 1.3507784e-25
+ luc = 1.9437196e-17
+ lint = 1.4999999e-8
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ wmax = 1.000869946e-5
+ wketa = 8.724413e-9
+ pvth0 = -2.3104256e-15
+ pa0 = 1.0862038e-13
+ nlx = 0.0
+ wmin = 1.20869946e-6
+ drout = 0.0
+ lkt1 = -2.4825255e-9
+ lkt2 = -1.0989117e-10
+ tpbsw = 0.001572025
+ pk1 = -1.7383759e-14
+ pk2 = 7.484627e-15
+ lmax = 4.94740781e-7
+ pu0 = 2.5785697e-16
+ lmin = 1.8e-7
+ ppdiblc2 = 8.594017e-17
+ prt = 0
+ pua = 1.5976873e-22
+ pub = -1.3085017e-31
+ puc = -9.356197e-24
+ cjswg = 4.43205e-10
+ wpdiblc2 = -1.9097854e-10
+ mjswg = 0.3683619
+ lnfactor = -3.9543e-9
+ rsh = 7.2
+ tcj = 0.0009739001
+ ua1 = 1.224e-9
+ ub1 = -1.3554493e-18
+ uc1 = 7.051652e-11
+ wvoff = 5.372431e-9
+ tpb = 0.001572025
+ tox = 4.13259219e-9
+ wub1 = -2.2890885e-25
+ wuc1 = -3.576699e-17
+ wa0 = -4.071248e-7
+ hdif = 2e-7
+ ute = -0.7199521
+ wk1 = 1.1998529e-7
+ wk2 = -4.424634e-8
+ weta0 = 0
+ tcjswg = 0.0004130718
+ lub1 = 2.6058948e-26
+ luc1 = -7.658915e-18
+ wln = 1.0
+ wetab = -5.480169e-10
+ lpdiblc2 = 9.0546e-10
+ wu0 = -2.5923497e-9
+ wute = 1.0915658e-7
+ mjsw = 0.3683619
+ wvsat = 0.0
+ wua = -6.282368e-16
+ wub = 3.0629255e-25
+ wuc = 1.4561782e-17
+ wwl = 0.0
+ wwn = 1.0
+ lpclm = 4.015361e-8
+ wvth0 = 7.955874e-9
+ xti = 3
+ lute = 6.205235e-10
+ cdsc = 0.0
+ wcdscd = 1.6464351e-11
+ cgdo = 3.116e-10
+ )

.model pch_ss_9 pmos (
+ level = 49
+ pvag = 0.0
+ etab = -5e-5
+ lvth0 = -3.9543e-9
+ ags = 0.02
+ vsat = 149999.98
+ wint = 5e-9
+ vth0 = -0.4523646
+ delta = 0.01
+ rdsw = 530.0
+ cit = -0.0001
+ wkt1 = 6.74333e-9
+ wkt2 = 1.2948118e-10
+ lint = 1.4999999e-8
+ dlc = 2e-9
+ wmax = 1.20869946e-6
+ dvt0w = 0.0
+ k3b = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ wmin = 5.086994599999999e-7
+ dwb = 0.0
+ dwg = 0.0
+ lmax = 2.0001e-5
+ lmin = 9.994740781e-6
+ capmod = 3
+ a0 = 0.9810578
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ jsw = 1.2e-12
+ kt1 = -0.2307052
+ kt2 = -0.02334808
+ lk2 = 1.18629e-9
+ wub1 = 3.495163e-26
+ wuc1 = 1.9335648e-17
+ at = 10000.0
+ cf = 0
+ cj = 0.00117705
+ ef = 1.064
+ k1 = 0.5449055
+ k2 = 0.0393854
+ k3 = 0.0
+ em = 30000000.0
+ llc = -0.039
+ lln = -1
+ lu0 = -7.9086e-11
+ hdif = 2e-7
+ js = 2.5e-7
+ ll = 0.0
+ mj = 0.4476
+ lw = 0.0
+ u0 = 0.0100768048
+ nch = 3.9e+17
+ pb = 0.895226
+ w0 = 0.0
+ rd = 0
+ lwl = 0.0
+ lwn = 1.0
+ rs = 0
+ ua = 1.0698959e-9
+ ub = 3.0837888e-19
+ uc = -1.1659398e-10
+ wl = 0.0
+ wute = -2.7886795e-9
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -1.4740781e-8
+ ww = 0.0
+ xw = -8.69946e-9
+ mjsw = 0.3683619
+ nlx = 0.0
+ tcjsw = 0.0004130718
+ mobmod = 1
+ pu0 = 0.0
+ pvoff = 0.0
+ prt = 0
+ rsh = 7.2
+ cdscb = 0.0
+ cdscd = 0.0
+ tcj = 0.0009739001
+ peta0 = 1.8966694548261387e-25
+ cdsc = 0.0
+ ua1 = 1.224e-9
+ ub1 = -1.3711068e-18
+ uc1 = 1.6263793e-12
+ tpb = 0.001572025
+ tox = 4.13259219e-9
+ cgdo = 3.116e-10
+ wketa = -1.0458587e-9
+ wa0 = 3.529885e-8
+ pvth0 = -1.18629e-15
+ drout = 0.0
+ ute = -0.7480742
+ wk1 = 2.1990281e-9
+ cgso = 3.116e-10
+ wk2 = -3.824582e-9
+ tpbsw = 0.001572025
+ wln = 1.0
+ wu0 = -2.481951e-10
+ wua = -1.3891575e-16
+ wub = -1.2660565e-25
+ wuc = -3.428342e-17
+ wwl = 0.0
+ wwn = 1.0
+ cjswg = 4.43205e-10
+ nfactor = 1.0
+ xti = 3
+ cjsw = 2.60505e-10
+ mjswg = 0.3683619
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ wvoff = -4.105241e-10
+ tcjswg = 0.0004130718
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0009999998
+ weta0 = 0
+ tnom = 25.0
+ pdiblcb = 0.01
+ wvsat = 0.0
+ wvth0 = -1.5613511000000001e-9
+ toxm = 4.08e-9
+ pbsw = 0.895226
+ pclm = 0.6
+ binunit = 2
+ pnfactor = 0
+ wnfactor = 0.0
+ keta = 0.03217546
+ xpart = 1
+ lnfactor = -3.9543e-9
+ alpha0 = 0.0
+ dsub = 0.0
+ alpha1 = 6.8730453846
+ pbswg = 0.895226
+ pscbe1 = 199999970.0
+ pscbe2 = 5e-7
+ dvt0 = 0.0
+ version = 3.24
+ dvt1 = 0.0
+ dvt2 = 0.0
+ lvoff = -1.5817200000000002e-9
+ voff = -0.12801
+ beta0 = 22.67827
+ nqsmod = 0
+ ldif = 9e-8
+ tpbswg = 0.001572025
+ noimod = 2
+ leta0 = 1.8966694548261387e-18
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ eta0 = 5e-5
+ )

.model pch_ss_10 pmos (
+ level = 49
+ dsub = 0.0
+ wk1 = 1.7598129e-9
+ wk2 = -3.600003e-9
+ wln = 1.0
+ wu0 = -2.1789574e-10
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ wua = -1.6455617e-16
+ wub = -7.150721e-26
+ wuc = -2.8652769e-17
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ wwl = 0.0
+ wwn = 1.0
+ xti = 3
+ pscbe1 = 180397680.0
+ pscbe2 = 5e-7
+ voff = -0.1269095
+ ldif = 9e-8
+ nfactor = 1.0
+ kt1l = 0.0
+ prwb = 0.0
+ pub1 = -8.629597e-32
+ prwg = 0.0
+ puc1 = 1.5034668e-23
+ nqsmod = 0
+ tpbswg = 0.001572025
+ lketa = -6.417587e-9
+ eta0 = 5e-5
+ noimod = 2
+ pvag = 0.0
+ etab = -5e-5
+ vsat = 151306.8
+ wint = 5e-9
+ pute = 3.909688e-14
+ xpart = 1
+ vth0 = -0.4482969
+ rdsw = 530.0
+ wkt1 = 6.495125e-9
+ wkt2 = 2.3726165e-10
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0004772722
+ lint = 1.4999999e-8
+ pdiblcb = 0.01
+ lpscbe1 = 195.04263
+ wmax = 1.20869946e-6
+ pbswg = 0.895226
+ wmin = 5.086994599999999e-7
+ lkt1 = -1.0252924e-8
+ lkt2 = -3.947785e-10
+ lmax = 9.994740781e-6
+ lvoff = -1.2530685e-8
+ lmin = 1.194740781e-6
+ beta0 = 22.67827
+ binunit = 2
+ leta0 = 1.8966694548261387e-18
+ lvsat = -0.013002842
+ lvth0 = -4.442723e-8
+ wub1 = 4.362458e-26
+ wuc1 = 1.7824627e-17
+ capmod = 3
+ hdif = 2e-7
+ delta = 0.01
+ lub1 = 7.318341e-26
+ luc1 = 2.7641896e-17
+ pnfactor = 0
+ wute = -6.718015e-9
+ mjsw = 0.3683619
+ wnfactor = 0.0
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ lute = 6.013659e-8
+ mobmod = 1
+ cdsc = 0.0
+ version = 3.24
+ lnfactor = -3.9543e-9
+ pketa = -1.6621007e-15
+ cgdo = 3.116e-10
+ ags = 0.02
+ cgso = 3.116e-10
+ cit = -0.0001
+ tcjsw = 0.0004130718
+ dlc = 2e-9
+ lpdiblc2 = 5.201137e-9
+ cjsw = 2.60505e-10
+ k3b = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ pvoff = 6.87864e-15
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 1.8966694548261387e-25
+ tcjswg = 0.0004130718
+ tnom = 25.0
+ wketa = -8.788133e-10
+ pvth0 = 1.274698e-14
+ la0 = 1.2176828e-7
+ drout = 0.0
+ toxm = 4.08e-9
+ jsw = 1.2e-12
+ kt1 = -0.2296747
+ lk1 = 1.9542425e-8
+ kt2 = -0.023308404
+ lk2 = -3.950429e-9
+ tpbsw = 0.001572025
+ pbsw = 0.895226
+ llc = -0.039
+ pclm = 0.5738636
+ lln = -1
+ lu0 = -1.0342642e-9
+ lua = -5.815077e-16
+ lub = 1.1186816e-24
+ luc = 7.427734e-17
+ nch = 3.9e+17
+ a0 = 0.9688198
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ lwl = 0.0
+ lwn = 1.0
+ cjswg = 4.43205e-10
+ at = 10000.0
+ cf = 0
+ cj = 0.00117705
+ pa0 = 3.87773e-15
+ nlx = 0.0
+ ef = 1.064
+ k1 = 0.5429414
+ k2 = 0.039901660000000005
+ k3 = 0.0
+ em = 30000000.0
+ mjswg = 0.3683619
+ js = 2.5e-7
+ ll = 0.0
+ mj = 0.4476
+ lw = 0.0
+ pk1 = 4.370194e-15
+ pk2 = -2.2345663e-15
+ u0 = 0.0101728028
+ pb = 0.895226
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ua = 1.1283389e-9
+ ub = 1.9594849e-19
+ uc = -1.2405904e-10
+ wvoff = -1.1018445e-9
+ wl = 0.0
+ pu0 = -3.0147877e-16
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -1.4740781e-8
+ ww = 0.0
+ xw = -8.69946e-9
+ prt = 0
+ pua = 2.5512236e-22
+ pub = -5.482294e-31
+ puc = -5.602498e-23
+ weta0 = 0
+ rsh = 7.2
+ tcj = 0.0009739001
+ ua1 = 1.224e-9
+ ub1 = -1.3784619e-18
+ uc1 = -1.1517035e-12
+ wvsat = 0.0
+ pkt1 = 2.469645e-15
+ pkt2 = -1.0724159e-15
+ keta = 0.03282044
+ tpb = 0.001572025
+ tox = 4.13259219e-9
+ lpclm = 2.6005682e-7
+ wvth0 = -2.9616815e-9
+ wa0 = 3.490912e-8
+ ute = -0.754118
+ )

.model pch_ss_11 pmos (
+ level = 49
+ cgso = 3.116e-10
+ a0 = 1.1936638
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ lvoff = 3.655491e-9
+ at = 10000.0
+ cf = 0
+ cj = 0.00117705
+ ef = 1.064
+ k1 = 0.4715038
+ k2 = 0.06532277
+ k3 = 0.0
+ em = 30000000.0
+ js = 2.5e-7
+ ll = 0.0
+ mj = 0.4476
+ lw = 0.0
+ beta0 = 22.67827
+ u0 = 0.0106717438
+ pb = 0.895226
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ua = 1.036115e-9
+ ub = 1.0523674e-18
+ uc = -7.205117e-11
+ cjsw = 2.60505e-10
+ leta0 = 3.696426189666945e-11
+ wl = 0.0
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -1.4740781e-8
+ ww = 0.0
+ xw = -8.69946e-9
+ letab = -3.696426e-11
+ lvsat = -0.007392855
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ capmod = 3
+ lvth0 = -7.517002e-9
+ delta = 0.01
+ tnom = 25.0
+ ags = 0.02
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ toxm = 4.08e-9
+ mobmod = 1
+ pcit = -1.0851648e-17
+ pbsw = 0.895226
+ pclm = 0.6714286
+ cit = -0.00031597191
+ dlc = 2e-9
+ k3b = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ pketa = 4.024799e-15
+ la0 = -1.3680231e-7
+ pkt1 = -6.051915e-15
+ pkt2 = -1.4802061e-15
+ tcjsw = 0.0004130718
+ keta = 0.03584265
+ jsw = 1.2e-12
+ kt1 = -0.2439705
+ lk1 = 1.0169572e-7
+ kt2 = -0.025852976
+ lk2 = -3.3184709999999996e-8
+ llc = -0.039
+ lln = -1
+ lu0 = -1.6080454999999999e-9
+ dsub = 0.0
+ pvoff = -3.866879e-15
+ lua = -4.754501e-16
+ lub = 1.337998e-25
+ luc = 1.4468274e-17
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ pa0 = 1.8891395e-13
+ nlx = 0.0
+ tcjswg = 0.0004130718
+ wcit = 9.436221e-12
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ pk1 = -6.35241e-14
+ pk2 = 2.2224691e-14
+ peta0 = 1.8966694548261387e-25
+ pu0 = 7.878928e-16
+ pnfactor = 0
+ prt = 0
+ lcit = 2.4836766e-10
+ pua = 2.5287059e-22
+ pub = -5.865131e-32
+ puc = -1.2704817e-23
+ wketa = -5.823942e-9
+ voff = -0.1409845
+ pvth0 = -6.289198e-15
+ wnfactor = 0.0
+ ldif = 9e-8
+ drout = 0.0
+ kt1l = 0.0
+ tpbsw = 0.001572025
+ prwb = 0.0
+ pub1 = 4.97241e-32
+ prwg = 0.0
+ rsh = 7.2
+ puc1 = 1.7282469e-23
+ tcj = 0.0009739001
+ ua1 = 1.224e-9
+ ub1 = -1.2162624e-18
+ uc1 = 4.210797e-11
+ eta0 = 1.7857154e-5
+ nfactor = 1.0
+ pvag = 0.0
+ etab = -1.7857154e-5
+ tpb = 0.001572025
+ tox = 4.13259219e-9
+ cjswg = 4.43205e-10
+ vsat = 146428.56
+ wa0 = -1.2599192e-7
+ wint = 5e-9
+ pute = -5.928695e-14
+ mjswg = 0.3683619
+ vth0 = -0.4803928
+ ute = -0.7903757
+ wk1 = 6.079834e-8
+ wk2 = -2.4868919e-8
+ rdsw = 530.0
+ wln = 1.0
+ wkt1 = 1.3905176e-8
+ wkt2 = 5.918618e-10
+ lnfactor = -3.9543e-9
+ wu0 = -1.1651754e-9
+ lint = 1.4999999e-8
+ wvoff = 8.242083e-9
+ wua = -1.625981e-16
+ wmax = 1.20869946e-6
+ wub = -4.972273e-25
+ wuc = -6.632247e-17
+ wwl = 0.0
+ wwn = 1.0
+ wmin = 5.086994599999999e-7
+ xti = 3
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0017857137
+ lkt1 = 6.187276e-9
+ lkt2 = 2.5314804e-9
+ pdiblcb = 0.01
+ weta0 = 0
+ lmax = 1.194740781e-6
+ lmin = 4.94740781e-7
+ wvsat = 0.0
+ lpclm = 1.4785714e-7
+ wvth0 = 1.3591517e-8
+ lpdiblc2 = 3.696429e-9
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ binunit = 2
+ pscbe1 = 349999900.0
+ pscbe2 = 5e-7
+ wub1 = -7.465372e-26
+ wuc1 = 1.5870021e-17
+ hdif = 2e-7
+ lub1 = -1.133461e-25
+ luc1 = -2.2106738e-17
+ wute = 7.883313e-8
+ mjsw = 0.3683619
+ nqsmod = 0
+ tpbswg = 0.001572025
+ noimod = 2
+ lute = 1.0183292e-7
+ lketa = -9.893122e-9
+ xpart = 1
+ cdsc = 0.0
+ cgdo = 3.116e-10
+ pbswg = 0.895226
+ version = 3.24
+ )

.model pch_ss_12 pmos (
+ level = 49
+ wint = 5e-9
+ llc = -0.039
+ pute = 1.3160581e-15
+ lln = -1
+ lu0 = 1.3290007e-10
+ vth0 = -0.47008160000000004
+ nfactor = 1.0
+ lua = 2.3815556e-17
+ lub = -3.425063e-26
+ luc = 8.803578e-18
+ nch = 3.9e+17
+ rdsw = 530.0
+ lwl = 0.0
+ lwn = 1.0
+ pketa = -9.609158e-16
+ wkt1 = 2.7434011e-10
+ wkt2 = -6.113567e-9
+ lint = 1.4999999e-8
+ pa0 = -8.476619e-14
+ nlx = 0.0
+ wmax = 1.20869946e-6
+ pk1 = 1.5213101e-14
+ pk2 = -6.235986e-15
+ wmin = 5.086994599999999e-7
+ lkt1 = -4.083267e-9
+ lkt2 = -2.4314675e-9
+ wpclm = 5.671285e-8
+ pu0 = -1.4287007e-16
+ lmax = 4.94740781e-7
+ prt = 0
+ pua = -7.799214e-23
+ pub = 7.065072e-32
+ puc = 3.297807e-24
+ lmin = 1.8e-7
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.009150297
+ tcjsw = 0.0004130718
+ pdiblcb = 0.01
+ rsh = 7.2
+ tcj = 0.0009739001
+ ua1 = 1.224e-9
+ ub1 = -1.6175756e-18
+ uc1 = -2.2818641e-11
+ pvoff = -1.4343533e-15
+ tcjswg = 0.0004130718
+ tpb = 0.001572025
+ tox = 4.13259219e-9
+ a0 = 0.5166956
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ wa0 = 4.821862e-7
+ at = 10000.0
+ cf = 0
+ cj = 0.00117705
+ wub1 = 8.30214e-26
+ ute = -0.5812994
+ wuc1 = 7.530186e-17
+ ef = 1.064
+ k1 = 0.7171482
+ k2 = -0.021956119
+ k3 = 0.0
+ em = 30000000.0
+ wk1 = -1.1417325e-7
+ wk2 = 3.837703e-8
+ binunit = 2
+ cdscb = 0.0
+ cdscd = -5.200001e-5
+ peta0 = 1.8966694548261387e-25
+ js = 2.5e-7
+ ll = 0.0
+ mj = 0.4476
+ hdif = 2e-7
+ lw = 0.0
+ u0 = 0.0068029748
+ wln = 1.0
+ pb = 0.895226
+ w0 = 0.0
+ wu0 = 9.031869e-10
+ rd = 0
+ rs = 0
+ ua = -7.336427e-11
+ ub = 1.4258127e-18
+ uc = -5.946296e-11
+ lub1 = 6.724484e-26
+ wua = 5.726523e-16
+ wub = -7.845651e-25
+ wuc = -1.0188386e-16
+ wl = 0.0
+ luc1 = 7.110234e-18
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -1.4740781e-8
+ ww = 0.0
+ xw = -8.69946e-9
+ wwl = 0.0
+ wwn = 1.0
+ wute = -5.584022e-8
+ wketa = 5.255423e-9
+ mjsw = 0.3683619
+ pvth0 = -2.2215402e-15
+ xti = 3
+ drout = 0.0
+ tpbsw = 0.001572025
+ lute = 7.748556e-9
+ wcdscd = -2.0304376e-11
+ cjswg = 4.43205e-10
+ mjswg = 0.3683619
+ cdsc = 0.0
+ wvoff = 2.8364715e-9
+ cgdo = 3.116e-10
+ pcdscd = 9.13697e-18
+ cgso = 3.116e-10
+ weta0 = 0
+ version = 3.24
+ wvsat = 0.0
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ lpclm = 6.365384e-8
+ wvth0 = 4.552275e-9
+ cjsw = 2.60505e-10
+ pscbe1 = 350000000.0
+ pscbe2 = 5e-7
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ nqsmod = 0
+ tpbswg = 0.001572025
+ tnom = 25.0
+ pnfactor = 0
+ noimod = 2
+ pags = -5.667374e-15
+ wnfactor = 0.0
+ toxm = 4.08e-9
+ pcit = 2.6834248e-18
+ pbsw = 0.895226
+ lketa = -1.8239428e-9
+ pclm = 0.858547
+ xpart = 1
+ ppdiblc2 = 7.08422e-16
+ wpdiblc2 = -1.5742713e-9
+ lnfactor = -3.9543e-9
+ pbswg = 0.895226
+ lcdscd = 2.3400004e-11
+ lvoff = -1.8855486300000003e-9
+ ags = 0.010547621
+ beta0 = 22.67827
+ pkt1 = 8.196091e-17
+ pkt2 = 1.5372367e-15
+ keta = 0.01791114
+ lpdiblc2 = 3.823661e-10
+ leta0 = 2.5593747189666946e-10
+ capmod = 3
+ letab = -3.473438e-10
+ cit = 0.00012746976
+ wags = 1.2594167e-8
+ lvsat = -0.0003656142
+ dsub = 0.0
+ dlc = 2e-9
+ lvth0 = -1.2157019e-8
+ k3b = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ lags = 4.253569e-9
+ wcit = -2.0641719e-11
+ ppclm = -2.5520774e-14
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ delta = 0.01
+ mobmod = 1
+ lcit = 4.881893e-11
+ voff = -0.1286711
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ ldif = 9e-8
+ kt1l = 0.0
+ prwb = 0.0
+ pub1 = -2.1229706e-32
+ prwg = 0.0
+ puc1 = -9.461855e-24
+ la0 = 1.6783336e-7
+ eta0 = -0.00046875
+ pvag = 0.0
+ jsw = 1.2e-12
+ etab = 0.0006718753
+ kt1 = -0.2211471
+ lk1 = -8.844278e-9
+ kt2 = -0.014824204
+ lk2 = 6.090789e-9
+ vsat = 130812.46
+ )

.model pch_ss_13 pmos (
+ level = 49
+ wketa = -6.403492e-9
+ pvth0 = -1.18629e-15
+ drout = 0.0
+ toxm = 4.08e-9
+ tpbsw = 0.001572025
+ pbsw = 0.895226
+ pclm = 0.5999999
+ cjswg = 4.43205e-10
+ mjswg = 0.3683619
+ wvoff = -1.320298e-9
+ weta0 = 0
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ wvsat = 0.0
+ keta = 0.04310941
+ pscbe1 = 199999970.0
+ pscbe2 = 5e-7
+ wvth0 = 8.154323e-9
+ dsub = 0.0
+ nqsmod = 0
+ tpbswg = 0.001572025
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ noimod = 2
+ voff = -0.1261533
+ ldif = 9e-8
+ a0 = 0.8704194
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ at = 10000.0
+ cf = 0
+ cj = 0.00117705
+ ef = 1.064
+ k1 = 0.5421249
+ k2 = 0.04121244
+ k3 = 0.0
+ em = 30000000.0
+ ags = 0.02
+ eta0 = 5e-5
+ js = 2.5e-7
+ ll = 0.0
+ mj = 0.4476
+ lw = 0.0
+ pvag = 0.0
+ etab = -5e-5
+ u0 = 0.0096929738
+ pb = 0.895226
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ vsat = 149999.98
+ xpart = 1
+ ua = 1.2584637e-9
+ ub = 4.999999e-20
+ uc = -1.6065008e-10
+ wint = 5e-9
+ wl = 0.0
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -1.4740781e-8
+ ww = 0.0
+ xw = -8.69946e-9
+ cit = -0.0001
+ vth0 = -0.4721925
+ rdsw = 530.0
+ dlc = 2e-9
+ wkt1 = 3.830554e-9
+ wkt2 = 1.9527771e-9
+ k3b = 0.0
+ lint = 1.4999999e-8
+ pbswg = 0.895226
+ dwb = 0.0
+ wmax = 5.086994599999999e-7
+ dwg = 0.0
+ nfactor = 1.0
+ wmin = 2.2e-7
+ lvoff = -1.5817200000000002e-9
+ lmax = 2.0001e-5
+ lmin = 9.994740781e-6
+ capmod = 3
+ beta0 = 22.67827
+ leta0 = 1.8966694548261387e-18
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.001
+ pdiblcb = 0.01
+ jsw = 1.2e-12
+ kt1 = -0.2247607
+ kt2 = -0.027069092
+ lk2 = 1.18629e-9
+ lvth0 = -3.9543e-9
+ llc = -0.039
+ lln = -1
+ lu0 = -7.9086e-11
+ wub1 = 2.1644123e-27
+ wuc1 = -1.2526765e-17
+ nch = 3.9e+17
+ mobmod = 1
+ lwl = 0.0
+ lwn = 1.0
+ delta = 0.01
+ hdif = 2e-7
+ nlx = 0.0
+ pnfactor = 0
+ binunit = 2
+ wute = 6.898109e-9
+ mjsw = 0.3683619
+ wnfactor = 0.0
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ pu0 = 0.0
+ prt = 0
+ rsh = 7.2
+ tcj = 0.0009739001
+ ua1 = 1.224e-9
+ ub1 = -1.3041941e-18
+ uc1 = 6.665171e-11
+ cdsc = 0.0
+ tpb = 0.001572025
+ tox = 4.13259219e-9
+ wa0 = 8.951166e-8
+ lnfactor = -3.9543e-9
+ cgdo = 3.116e-10
+ ute = -0.7678431
+ wk1 = 3.561511e-9
+ wk2 = -4.719829e-9
+ wln = 1.0
+ cgso = 3.116e-10
+ wu0 = -6.011836e-11
+ wua = -2.3131395e-16
+ wuc = -1.2695932e-17
+ wwl = 0.0
+ wwn = 1.0
+ xti = 3
+ tcjsw = 0.0004130718
+ tcjswg = 0.0004130718
+ version = 3.24
+ cjsw = 2.60505e-10
+ pvoff = 0.0
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 1.8966694548261387e-25
+ tnom = 25.0
+ )

.model pch_ss_14 pmos (
+ level = 49
+ tpbswg = 0.001572025
+ noimod = 2
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0004772729
+ cit = -0.0001
+ wub1 = -3.0198158e-27
+ wuc1 = -1.0513175e-17
+ pdiblcb = 0.01
+ lpscbe1 = 195.04262
+ dlc = 2e-9
+ hdif = 2e-7
+ k3b = 0.0
+ lub1 = -2.0820251e-25
+ dwb = 0.0
+ dwg = 0.0
+ luc1 = 9.921307e-17
+ wute = 1.1298283e-8
+ mjsw = 0.3683619
+ binunit = 2
+ lketa = -4.562476e-8
+ lute = 2.2927659e-7
+ xpart = 1
+ la0 = 5.081137e-7
+ cdsc = 0.0
+ jsw = 1.2e-12
+ kt1 = -0.2237138
+ lk1 = -4.88067e-8
+ kt2 = -0.026908273
+ lk2 = 2.4488488e-8
+ llc = -0.039
+ lln = -1
+ cgdo = 3.116e-10
+ lu0 = -3.7909119e-10
+ pbswg = 0.895226
+ lua = -3.24011e-17
+ lub = -3.941427e-28
+ luc = -6.882293e-17
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ cgso = 3.116e-10
+ pa0 = -1.854315e-13
+ lvoff = -3.9703229000000005e-9
+ nlx = 0.0
+ capmod = 3
+ pk1 = 3.786126e-14
+ pk2 = -1.6169635e-14
+ beta0 = 22.67827
+ pu0 = -6.225135e-16
+ leta0 = 1.8966694548261387e-18
+ prt = 0
+ pua = -1.3939852e-23
+ pub = 1.1764949e-34
+ puc = 1.4094153e-23
+ cjsw = 2.60505e-10
+ lvsat = -0.013002842
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ lvth0 = -8.562635e-9
+ version = 3.24
+ rsh = 7.2
+ tcj = 0.0009739001
+ mobmod = 1
+ ua1 = 1.224e-9
+ ub1 = -1.2832692e-18
+ uc1 = 5.668055e-11
+ tpb = 0.001572025
+ tox = 4.13259219e-9
+ delta = 0.01
+ wa0 = 1.0814799e-7
+ tnom = 25.0
+ ute = -0.790886
+ wk1 = -2.4364055e-10
+ wk2 = -3.0947396e-9
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ wln = 1.0
+ wu0 = 2.4458129999999986e-12
+ toxm = 4.08e-9
+ wua = -2.2991296e-16
+ wub = -1.1822094e-29
+ wuc = -1.4112429e-17
+ wwl = 0.0
+ wwn = 1.0
+ pbsw = 0.895226
+ xti = 3
+ pclm = 0.5738635
+ pketa = 1.7549415e-14
+ a0 = 0.8193527
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ at = 10000.0
+ cf = 0
+ cj = 0.00117705
+ ef = 1.064
+ k1 = 0.5470301
+ k2 = 0.038870510000000004
+ k3 = 0.0
+ em = 30000000.0
+ js = 2.5e-7
+ ll = 0.0
+ mj = 0.4476
+ lw = 0.0
+ u0 = 0.0097231258
+ pb = 0.895226
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ua = 1.2617201e-9
+ ub = 5.00396e-20
+ uc = -1.5373321e-10
+ wl = 0.0
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -1.4740781e-8
+ ww = 0.0
+ tcjswg = 0.0004130718
+ xw = -8.69946e-9
+ tcjsw = 0.0004130718
+ pkt1 = 2.5501714e-15
+ pkt2 = -4.817884e-16
+ keta = 0.04769481
+ pvoff = 2.6840621e-15
+ dsub = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 1.8966694548261387e-25
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ pnfactor = 0
+ wketa = -8.167253e-9
+ pvth0 = -4.826672e-15
+ wnfactor = 0.0
+ voff = -0.1259132
+ drout = 0.0
+ ldif = 9e-8
+ tpbsw = 0.001572025
+ kt1l = 0.0
+ prwb = 0.0
+ pub1 = 5.158311e-32
+ prwg = 0.0
+ puc1 = -2.0035212e-23
+ eta0 = 5e-5
+ cjswg = 4.43205e-10
+ pvag = 0.0
+ etab = -5e-5
+ vsat = 151306.8
+ mjswg = 0.3683619
+ wint = 5e-9
+ pute = -4.378173e-14
+ vth0 = -0.4717293
+ rdsw = 530.0
+ lnfactor = -3.9543e-9
+ wvoff = -1.590053e-9
+ wkt1 = 3.574256e-9
+ wkt2 = 2.0011981e-9
+ lint = 1.4999999e-8
+ wmax = 5.086994599999999e-7
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ wmin = 2.2e-7
+ lkt1 = -1.0417262e-8
+ lkt2 = -1.6001408e-9
+ weta0 = 0
+ nfactor = 1.0
+ lmax = 9.994740781e-6
+ pscbe1 = 180397700.0
+ pscbe2 = 5e-7
+ wvsat = 0.0
+ lmin = 1.194740781e-6
+ lpclm = 2.6005691e-7
+ wvth0 = 8.52019e-9
+ lpdiblc2 = 5.201136e-9
+ ags = 0.02
+ nqsmod = 0
+ )

.model pch_ss_15 pmos (
+ level = 49
+ ute = -0.5904401
+ wk1 = 4.182789e-8
+ wk2 = -2.2085489e-8
+ beta0 = 22.67827
+ wln = 1.0
+ wu0 = -4.185056e-10
+ pkt1 = -8.599671e-15
+ pkt2 = 1.9347028e-16
+ lpdiblc2 = 3.696429e-9
+ keta = 0.0004484208
+ wua = -1.9008923e-16
+ leta0 = 3.6964281896669455e-11
+ wub = 8.369847e-27
+ wuc = 5.370726e-18
+ wwl = 0.0
+ wwn = 1.0
+ letab = -3.696428e-11
+ xti = 3
+ mobmod = 1
+ lvsat = -0.007392816
+ dsub = 0.0
+ lvth0 = -1.9486833e-8
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ delta = 0.01
+ lcit = 2.2622144e-10
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ voff = -0.1186655
+ ldif = 9e-8
+ kt1l = 0.0
+ prwb = 0.0
+ pub1 = -1.2589071e-33
+ prwg = 0.0
+ puc1 = 4.27717e-24
+ eta0 = 1.7857146e-5
+ pvag = 0.0
+ etab = -1.7857146e-5
+ vsat = 146428.52
+ wint = 5e-9
+ pute = -8.783067e-15
+ vth0 = -0.46223000000000003
+ rdsw = 530.0
+ pketa = -5.090041e-15
+ wkt1 = 1.3269771e-8
+ wkt2 = 1.4140165e-9
+ lint = 1.4999999e-8
+ wmax = 5.086994599999999e-7
+ tcjswg = 0.0004130718
+ wmin = 2.2e-7
+ lkt1 = 1.1386779e-8
+ lkt2 = -8.841858e-10
+ lmax = 1.194740781e-6
+ lmin = 4.94740781e-7
+ tcjsw = 0.0004130718
+ nfactor = 1.0
+ pvoff = 3.95383e-15
+ wub1 = 4.292976e-26
+ cdscb = 0.0
+ wuc1 = -3.165437e-17
+ cdscd = 0.0
+ peta0 = 1.8966694548261387e-25
+ hdif = 2e-7
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0017857139
+ pdiblcb = 0.01
+ lub1 = -9.299159e-27
+ wketa = 1.1519229e-8
+ luc1 = 4.434689e-18
+ pvth0 = -4.239814e-16
+ wute = -1.9135335e-8
+ mjsw = 0.3683619
+ drout = 0.0
+ tpbsw = 0.001572025
+ lute = -1.2362289e-9
+ cjswg = 4.43205e-10
+ binunit = 2
+ mjswg = 0.3683619
+ ags = 0.02
+ cdsc = 0.0
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ wvoff = -2.6941984e-9
+ cit = -0.00029671428
+ cgdo = 3.116e-10
+ pscbe1 = 349999900.0
+ pscbe2 = 5e-7
+ dlc = 2e-9
+ cgso = 3.116e-10
+ k3b = 0.0
+ weta0 = 0
+ dwb = 0.0
+ dwg = 0.0
+ wvsat = 0.0
+ lpclm = 1.4785714e-7
+ wvth0 = 4.691763999999999e-9
+ nqsmod = 0
+ a0 = 1.1508681
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ tpbswg = 0.001572025
+ cjsw = 2.60505e-10
+ noimod = 2
+ at = 10000.0
+ cf = 0
+ cj = 0.00117705
+ ef = 1.064
+ k1 = 0.510219
+ k2 = 0.0596423
+ k3 = 0.0
+ em = 30000000.0
+ js = 2.5e-7
+ ll = 0.0
+ noia = 9.5e+18
+ mj = 0.4476
+ noib = 100000.0
+ noic = 1.4e-12
+ lw = 0.0
+ u0 = 0.0091479268
+ pb = 0.895226
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ua = 1.0922192e-9
+ ub = 2.0536515e-20
+ uc = -2.183638e-10
+ la0 = 1.2687106e-7
+ wl = 0.0
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -1.4740781e-8
+ ww = 0.0
+ xw = -8.69946e-9
+ jsw = 1.2e-12
+ version = 3.24
+ kt1 = -0.2426738
+ lk1 = -6.473878e-9
+ kt2 = -0.027530843
+ lk2 = 6.009272e-10
+ llc = -0.039
+ lln = -1
+ pnfactor = 0
+ lu0 = 2.823877e-10
+ tnom = 25.0
+ lua = 1.6252487e-16
+ lub = 3.353441e-26
+ luc = 5.502275e-18
+ nch = 3.9e+17
+ wnfactor = 0.0
+ lwl = 0.0
+ lwn = 1.0
+ pa0 = 5.971399e-14
+ nlx = 0.0
+ toxm = 4.08e-9
+ lketa = 8.708591e-9
+ pk1 = -1.0521005e-14
+ pk2 = 5.669729e-15
+ pbsw = 0.895226
+ pclm = 0.6714286
+ pu0 = -1.384194e-16
+ xpart = 1
+ prt = 0
+ pua = -5.973716e-23
+ pub = -9.521269e-33
+ puc = -8.311478e-24
+ rsh = 7.2
+ lnfactor = -3.9543e-9
+ tcj = 0.0009739001
+ ua1 = 1.224e-9
+ ub1 = -1.4562286e-18
+ uc1 = 1.3909653e-10
+ pbswg = 0.895226
+ capmod = 3
+ tpb = 0.001572025
+ tox = 4.13259219e-9
+ wa0 = -1.0502199e-7
+ lvoff = -1.2305139000000001e-8
+ )

.model pch_ss_16 pmos (
+ level = 49
+ cdsc = 0.0
+ binunit = 2
+ pketa = 7.45672e-16
+ lnfactor = -3.9543e-9
+ tcjswg = 0.0004130718
+ cgdo = 3.116e-10
+ wpclm = 4.634222e-9
+ cgso = 3.116e-10
+ tcjsw = 0.0004130718
+ lpdiblc2 = 1.8281252e-9
+ cjsw = 2.60505e-10
+ pvoff = 1.4541431e-15
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ wcdscd = -1.4183201e-11
+ ags = 0.03625
+ cdscb = 0.0
+ cdscd = -6.449223e-5
+ peta0 = 1.8966694548261387e-25
+ cit = 8.534377e-5
+ tnom = 25.0
+ wketa = -1.4490222e-9
+ pvth0 = -1.47043808e-15
+ version = 3.24
+ dlc = 2e-9
+ drout = 0.0
+ pcdscd = 6.382441e-18
+ tpbsw = 0.001572025
+ k3b = 0.0
+ toxm = 4.08e-9
+ dwb = 0.0
+ dwg = 0.0
+ pbsw = 0.895226
+ pclm = 0.9648299
+ cjswg = 4.43205e-10
+ mjswg = 0.3683619
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ wvoff = 2.8606606e-9
+ pscbe1 = 350000000.0
+ pscbe2 = 5e-7
+ la0 = 7.233052e-9
+ jsw = 1.2e-12
+ kt1 = -0.2130934
+ lk1 = 1.3789155e-8
+ kt2 = -0.03589084
+ lk2 = -1.920656e-9
+ llc = -0.039
+ weta0 = 0
+ lln = -1
+ lu0 = -4.357122e-10
+ nqsmod = 0
+ lua = -2.6402067e-16
+ lub = 2.6345733e-25
+ luc = 3.340897e-17
+ nch = 3.9e+17
+ wvsat = 0.0
+ tpbswg = 0.001572025
+ lwl = 0.0
+ lwn = 1.0
+ noimod = 2
+ lpclm = 1.5826547e-8
+ pa0 = -6.072043e-15
+ wvth0 = 7.017223000000001e-9
+ nlx = 0.0
+ pkt1 = -9.758805e-16
+ pkt2 = -1.0643102e-15
+ keta = 0.03159368
+ pk1 = 4.122718e-15
+ pk2 = -2.3103772e-15
+ dsub = 0.0
+ pu0 = 1.3574996e-16
+ prt = 0
+ pua = 6.304761e-23
+ pub = -7.522618e-32
+ puc = -8.758834e-24
+ lags = -7.312499e-9
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ rsh = 7.2
+ tcj = 0.0009739001
+ ua1 = 1.224e-9
+ ub1 = -1.4433942e-18
+ uc1 = 2.0396977e-10
+ tpb = 0.001572025
+ tox = 4.13259219e-9
+ lcit = 5.429531e-11
+ voff = -0.1287204
+ wa0 = 4.116919e-8
+ lcdscd = 2.9021494e-11
+ ldif = 9e-8
+ ute = -0.5893072
+ wk1 = 9.286284e-9
+ kt1l = 0.0
+ wk2 = -4.351921e-9
+ prwb = 0.0
+ pub1 = 1.9106841e-32
+ prwg = 0.0
+ lketa = -5.306775e-9
+ puc1 = 6.153712e-24
+ wln = 1.0
+ wu0 = -1.0277709000000001e-9
+ eta0 = -0.0004687502
+ wua = -4.629443e-16
+ pvag = 0.0
+ wub = 1.5438073e-25
+ wuc = 6.364847e-18
+ etab = 0.0006718753
+ xpart = 1
+ wwl = 0.0
+ wwn = 1.0
+ vsat = 130812.55
+ xti = 3
+ wint = 5e-9
+ pute = 5.968411e-15
+ vth0 = -0.47511210000000004
+ capmod = 3
+ rdsw = 530.0
+ wkt1 = -3.671987e-9
+ wkt2 = 4.209085e-9
+ pbswg = 0.895226
+ lint = 1.4999999e-8
+ wmax = 5.086994599999999e-7
+ wmin = 2.2e-7
+ lvoff = -7.780439e-9
+ lkt1 = -1.9244071e-9
+ lkt2 = 2.877812e-9
+ lmax = 4.94740781e-7
+ beta0 = 22.67827
+ lmin = 1.8e-7
+ mobmod = 1
+ leta0 = 2.559375818966695e-10
+ letab = -3.473438e-10
+ lvsat = -0.0003656336
+ nfactor = 1.0
+ lvth0 = -1.3689881e-8
+ ppclm = -2.0853998e-15
+ wub1 = -2.3274574e-27
+ wuc1 = -3.582447e-17
+ delta = 0.01
+ hdif = 2e-7
+ a0 = 1.4167303
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ pnfactor = 0
+ lub1 = -1.5074642e-26
+ luc1 = -2.4758267e-17
+ at = 10000.0
+ cf = 0
+ cj = 0.00117705
+ ef = 1.064
+ k1 = 0.46519
+ dvt0w = 0.0
+ k2 = 0.06524582
+ k3 = 0.0
+ em = 30000000.0
+ wnfactor = 0.0
+ wute = -5.191639e-8
+ dvt1w = 0.0
+ dvt2w = 0.0
+ mjsw = 0.3683619
+ js = 2.5e-7
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.005937499
+ ll = 0.0
+ mj = 0.4476
+ lw = 0.0
+ u0 = 0.0107437038
+ pb = 0.895226
+ w0 = 0.0
+ rd = 0
+ pdiblcb = 0.01
+ rs = 0
+ ua = 2.0400983e-9
+ ub = -4.904033e-19
+ uc = -2.8037866e-10
+ wl = 0.0
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -1.4740781e-8
+ ww = 0.0
+ lute = -1.7460413e-9
+ xw = -8.69946e-9
+ )

.model pch_ff_1 pmos (
+ level = 49
+ lvth0 = 3.9543e-9
+ cdsc = 0.0
+ binunit = 2
+ pnfactor = 0
+ cgdo = 3.444e-10
+ delta = 0.01
+ wnfactor = 0.0
+ cgso = 3.444e-10
+ dvt0w = 0.0
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ dvt1w = 0.0
+ dvt2w = 0.0
+ pscbe1 = 199999970.0
+ pscbe2 = 5e-7
+ cjsw = 2.35695e-10
+ ags = 0.02
+ lnfactor = 3.9543e-9
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ nqsmod = 0
+ tpbswg = 0.001572025
+ noimod = 2
+ cit = -0.0001
+ dlc = 2e-9
+ tnom = 25.0
+ version = 3.24
+ k3b = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ toxm = 4.08e-9
+ tcjsw = 0.0004130718
+ pbsw = 0.895226
+ pclm = 0.6000001
+ pvoff = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ jsw = 1.2e-12
+ peta0 = 4.7451600189666944e-17
+ kt1 = -0.2311294
+ lk2 = -1.18629e-9
+ kt2 = -0.02433992
+ llc = -0.039
+ lln = -1
+ lu0 = 7.9086e-11
+ nch = 3.9e+17
+ pvth0 = 1.18629e-15
+ lwl = 0.0
+ lwn = 1.0
+ drout = 0.0
+ nlx = 0.0
+ tpbsw = 0.001572025
+ capmod = 3
+ keta = 0.026632193
+ pu0 = 0.0
+ cjswg = 4.00995e-10
+ prt = 0
+ dsub = 0.0
+ mjswg = 0.3683619
+ rsh = 7.2
+ tcj = 0.0009739001
+ ua1 = 1.224e-9
+ ub1 = -1.3928839e-18
+ uc1 = -4.59467e-12
+ wvoff = 0.0
+ mobmod = 1
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ tpb = 0.001572025
+ tox = 4.02740781e-9
+ ute = -0.8288856
+ voff = -0.1275921
+ weta0 = 0
+ ldif = 9e-8
+ wvsat = 0.0
+ wln = 1.0
+ kt1l = 0.0
+ prwb = 0.0
+ wu0 = 1.97715e-11
+ prwg = 0.0
+ wvth0 = 1.18629e-9
+ wwl = 0.0
+ wwn = 1.0
+ eta0 = 5e-5
+ xti = 3
+ pvag = 0.0
+ etab = -5e-5
+ vsat = 149999.98
+ wint = 5e-9
+ vth0 = -0.4147553
+ rdsw = 530.0
+ lint = 1.4999999e-8
+ wmax = 0.000900001
+ wmin = 9.991300540000001e-6
+ a0 = 1.0461572
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ lmax = 2.0001e-5
+ at = 10000.0
+ cf = 0
+ cj = 0.00106495
+ lmin = 1.0005259219000001e-5
+ ef = 1.064
+ k1 = 0.5375325
+ k2 = 0.029496539999999998
+ k3 = 0.0
+ em = 30000000.0
+ tcjswg = 0.0004130718
+ js = 2.5e-7
+ ll = 0.0
+ mj = 0.4476
+ lw = 0.0
+ u0 = 0.0109204782
+ pb = 0.895226
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ua = 8.23294e-10
+ ub = 6.854322e-19
+ uc = -8.655411e-11
+ wl = 0.0
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -2.5259219000000002e-8
+ ww = 0.0
+ xw = 8.69946e-9
+ xpart = 1
+ nfactor = 1.0
+ pbswg = 0.895226
+ hdif = 2e-7
+ lvoff = 1.5817200000000002e-9
+ mjsw = 0.3683619
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0010000003
+ pdiblcb = 0.01
+ beta0 = 22.67827
+ leta0 = 4.745160018966694e-10
+ )

.model pch_ff_2 pmos (
+ level = 49
+ mj = 0.4476
+ lw = 0.0
+ kt1 = -0.2295883
+ lk1 = 1.8783622e-8
+ kt2 = -0.024031118
+ lk2 = -6.673462e-9
+ u0 = 0.0110505252
+ pb = 0.895226
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ua = 8.625313e-10
+ ub = 6.401998e-19
+ uc = -8.855145e-11
+ llc = -0.039
+ lln = -1
+ wl = 0.0
+ lu0 = -1.2148829000000001e-9
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -2.5259219000000002e-8
+ ww = 0.0
+ xw = 8.69946e-9
+ voff = -0.1274002
+ lua = -3.904111e-16
+ lub = 4.500626e-25
+ luc = 1.9873557e-17
+ ldif = 9e-8
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ kt1l = 0.0
+ tcjsw = 0.0004130718
+ prwb = 0.0
+ prwg = 0.0
+ nlx = 0.0
+ eta0 = 5e-5
+ pvag = 0.0
+ etab = -5e-5
+ pvoff = 0.0
+ vsat = 151306.8
+ pu0 = 0.0
+ wint = 5e-9
+ prt = 0
+ vth0 = -0.4122614
+ rdsw = 530.0
+ pnfactor = 0
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 4.7451600189666944e-17
+ lint = 1.4999999e-8
+ rsh = 7.2
+ tcj = 0.0009739001
+ ua1 = 1.224e-9
+ wnfactor = 0.0
+ wmax = 0.000900001
+ ub1 = -1.3977103e-18
+ uc1 = -6.694918e-12
+ wmin = 9.991300540000001e-6
+ tpb = 0.001572025
+ capmod = 3
+ pvth0 = 1.18629e-15
+ tox = 4.02740781e-9
+ lkt1 = -1.5333228e-8
+ lkt2 = -3.0725886e-9
+ drout = 0.0
+ lmax = 1.0005259219000001e-5
+ tpbsw = 0.001572025
+ ute = -0.8385549
+ lmin = 1.205259219e-6
+ wln = 1.0
+ wu0 = 1.97715e-11
+ cjswg = 4.00995e-10
+ wwl = 0.0
+ wwn = 1.0
+ mjswg = 0.3683619
+ lnfactor = 3.9543e-9
+ xti = 3
+ mobmod = 1
+ nfactor = 1.0
+ wvoff = 0.0
+ hdif = 2e-7
+ lub1 = 4.802326e-26
+ luc1 = 2.0897466e-17
+ weta0 = 0
+ mjsw = 0.3683619
+ lpdiblc2 = 5.201137e-9
+ wvsat = 0.0
+ lute = 9.620972e-8
+ lpclm = 2.6005682e-7
+ wvth0 = 1.18629e-9
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0004772727
+ pdiblcb = 0.01
+ lpscbe1 = 195.04263
+ cdsc = 0.0
+ cgdo = 3.444e-10
+ binunit = 2
+ cgso = 3.444e-10
+ tcjswg = 0.0004130718
+ lketa = -2.0462676e-9
+ cjsw = 2.35695e-10
+ xpart = 1
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ pbswg = 0.895226
+ tnom = 25.0
+ lvoff = -3.274108999999997e-10
+ toxm = 4.08e-9
+ beta0 = 22.67827
+ version = 3.24
+ pbsw = 0.895226
+ pclm = 0.5738637
+ leta0 = 4.745160018966694e-10
+ lvsat = -0.013002843
+ lvth0 = -2.0859753e-8
+ ags = 0.02
+ delta = 0.01
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ cit = -0.0001
+ dlc = 2e-9
+ dvt0w = 0.0
+ dvt1w = 0.0
+ pscbe1 = 180397680.0
+ pscbe2 = 5e-7
+ dvt2w = 0.0
+ k3b = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ keta = 0.026837848
+ nqsmod = 0
+ tpbswg = 0.001572025
+ dsub = 0.0
+ noimod = 2
+ a0 = 1.0385712
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ at = 10000.0
+ cf = 0
+ cj = 0.00106495
+ la0 = 7.548124e-8
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ ef = 1.064
+ k1 = 0.5356447
+ k2 = 0.030048010000000003
+ k3 = 0.0
+ em = 30000000.0
+ js = 2.5e-7
+ jsw = 1.2e-12
+ ll = 0.0
+ )

.model pch_ff_3 pmos (
+ level = 49
+ cjswg = 4.00995e-10
+ mjswg = 0.3683619
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ wvoff = 0.0
+ tnom = 25.0
+ weta0 = 0
+ wvsat = 0.0
+ toxm = 4.08e-9
+ a0 = 1.0045335
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ lpclm = 1.4785704e-7
+ wvth0 = 1.18629e-9
+ pbsw = 0.895226
+ pclm = 0.6714287
+ at = 10000.0
+ cf = 0
+ cj = 0.00106495
+ ef = 1.064
+ k1 = 0.5405614
+ k2 = 0.02936555
+ k3 = 0.0
+ em = 30000000.0
+ js = 2.5e-7
+ version = 3.24
+ ll = 0.0
+ mj = 0.4476
+ lw = 0.0
+ u0 = 0.0102799442
+ pb = 0.895226
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ua = 5.26694e-10
+ ub = 1.1734415e-18
+ uc = -4.332115e-11
+ wl = 0.0
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -2.5259219000000002e-8
+ ww = 0.0
+ xw = 8.69946e-9
+ pnfactor = 0
+ wnfactor = 0.0
+ tcjswg = 0.0004130718
+ lketa = -8.158225e-9
+ keta = 0.03215259
+ xpart = 1
+ dsub = 0.0
+ lnfactor = 3.9543e-9
+ ags = 0.02
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ pbswg = 0.895226
+ lvoff = 6.329375000000001e-10
+ lcit = 2.2402701e-10
+ cit = -0.00029480609
+ voff = -0.1282353
+ lpdiblc2 = 3.696428e-9
+ ldif = 9e-8
+ dlc = 2e-9
+ beta0 = 22.67827
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ k3b = 0.0
+ dwb = 0.0
+ leta0 = 5.114802818966694e-10
+ dwg = 0.0
+ eta0 = 1.7857143e-5
+ letab = -3.696428e-11
+ pvag = 0.0
+ etab = -1.7857143e-5
+ lvsat = -0.007392833
+ vsat = 146428.53
+ wint = 5e-9
+ lvth0 = -2.735142e-9
+ vth0 = -0.42802199999999996
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ rdsw = 530.0
+ delta = 0.01
+ lint = 1.4999999e-8
+ wmax = 0.000900001
+ pscbe1 = 349999900.0
+ pscbe2 = 5e-7
+ la0 = 1.146246e-7
+ wmin = 9.991300540000001e-6
+ jsw = 1.2e-12
+ lkt1 = 1.5747348e-9
+ lkt2 = 9.740028e-10
+ kt1 = -0.2442909
+ lk1 = 1.3129389e-8
+ kt2 = -0.027549893
+ lk2 = -5.888625e-9
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ lmax = 1.205259219e-6
+ llc = -0.039
+ lln = -1
+ lu0 = -3.287146e-10
+ lmin = 5.052592189999999e-7
+ lua = -4.198125e-18
+ lub = -1.631654e-25
+ luc = -3.214129e-17
+ nch = 3.9e+17
+ nqsmod = 0
+ lwl = 0.0
+ lwn = 1.0
+ tpbswg = 0.001572025
+ noimod = 2
+ nlx = 0.0
+ pu0 = 0.0
+ prt = 0
+ hdif = 2e-7
+ rsh = 7.2
+ tcj = 0.0009739001
+ nfactor = 1.0
+ ua1 = 1.224e-9
+ lub1 = 3.0810812e-26
+ ub1 = -1.3827429e-18
+ luc1 = 2.9752128e-17
+ uc1 = -1.4394627e-11
+ mjsw = 0.3683619
+ tpb = 0.001572025
+ tox = 4.02740781e-9
+ tcjsw = 0.0004130718
+ lute = 3.654092e-8
+ ute = -0.786669
+ wln = 1.0
+ pvoff = 0.0
+ wu0 = 1.97715e-11
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0017857148
+ wwl = 0.0
+ wwn = 1.0
+ pdiblcb = 0.01
+ cdsc = 0.0
+ xti = 3
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 4.7451600189666944e-17
+ capmod = 3
+ cgdo = 3.444e-10
+ pvth0 = 1.18629e-15
+ cgso = 3.444e-10
+ drout = 0.0
+ binunit = 2
+ tpbsw = 0.001572025
+ cjsw = 2.35695e-10
+ mobmod = 1
+ )

.model pch_ff_4 pmos (
+ level = 49
+ wmin = 9.991300540000001e-6
+ lkt1 = -2.665e-9
+ lkt2 = -2.325577e-10
+ lmax = 5.052592189999999e-7
+ cit = -4.054396e-5
+ lmin = 1.8e-7
+ lketa = -8.307595e-10
+ dlc = 2e-9
+ k3b = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ xpart = 1
+ pbswg = 0.895226
+ hdif = 2e-7
+ lub1 = 2.883988e-26
+ luc1 = -6.846759e-18
+ lvoff = 1.5460040800000002e-9
+ la0 = 1.6196543e-8
+ mjsw = 0.3683619
+ jsw = 1.2e-12
+ kt1 = -0.2348693
+ lk1 = 1.6807924e-8
+ kt2 = -0.024868647
+ lk2 = -7.0625049999999995e-9
+ beta0 = 22.67827
+ nfactor = 1.0
+ llc = -0.039
+ lln = -1
+ lu0 = -1.9861809999999995e-11
+ lute = 1.6013461e-9
+ leta0 = 7.304535218966694e-10
+ lua = -1.5999061e-16
+ lub = 1.2197973e-25
+ luc = 1.8500639e-17
+ nch = 3.9e+17
+ letab = -5.298917e-10
+ lwl = 0.0
+ lwn = 1.0
+ lvsat = -0.0003656265
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ nlx = 0.0
+ lvth0 = -4.286252e-9
+ cdsc = 0.0
+ pscbe1 = 350000000.0
+ pscbe2 = 5e-7
+ pnfactor = 0
+ pu0 = 0.0
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.00796875
+ delta = 0.01
+ a0 = 1.2232625
+ a1 = 0.0
+ a2 = 0.4
+ prt = 0
+ b0 = 0.0
+ b1 = 0.0
+ cgdo = 3.444e-10
+ wnfactor = 0.0
+ pdiblcb = 0.01
+ at = 10000.0
+ cf = 0
+ cj = 0.00106495
+ ef = 1.064
+ k1 = 0.5323869
+ k2 = 0.031974169999999996
+ k3 = 0.0
+ em = 30000000.0
+ cgso = 3.444e-10
+ js = 2.5e-7
+ dvt0w = 0.0
+ dvt1w = 0.0
+ ll = 0.0
+ rsh = 7.2
+ mj = 0.4476
+ dvt2w = 0.0
+ lw = 0.0
+ u0 = 0.0095936042
+ tcj = 0.0009739001
+ nqsmod = 0
+ pb = 0.895226
+ ua1 = 1.224e-9
+ w0 = 0.0
+ ub1 = -1.3783631e-18
+ rd = 0
+ uc1 = 6.693623e-11
+ tpbswg = 0.001572025
+ rs = 0
+ ua = 8.728995e-10
+ ub = 5.397856e-19
+ uc = -1.5585878e-10
+ noimod = 2
+ wl = 0.0
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -2.5259219000000002e-8
+ ww = 0.0
+ xw = 8.69946e-9
+ tpb = 0.001572025
+ tox = 4.02740781e-9
+ binunit = 2
+ cjsw = 2.35695e-10
+ ute = -0.7090256
+ lnfactor = 3.9543e-9
+ wln = 1.0
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ wu0 = 1.97715e-11
+ wwl = 0.0
+ wwn = 1.0
+ xti = 3
+ tnom = 25.0
+ lcdscd = 3.65625e-11
+ lpdiblc2 = 9.140626e-10
+ toxm = 4.08e-9
+ tcjsw = 0.0004130718
+ pbsw = 0.895226
+ pclm = 0.9102259
+ pvoff = 0.0
+ capmod = 3
+ version = 3.24
+ cdscb = 0.0
+ cdscd = -8.125e-5
+ peta0 = 4.7451600189666944e-17
+ pvth0 = 1.18629e-15
+ drout = 0.0
+ tpbsw = 0.001572025
+ mobmod = 1
+ keta = 0.015869336
+ cjswg = 4.00995e-10
+ mjswg = 0.3683619
+ dsub = 0.0
+ wvoff = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ weta0 = 0
+ lcit = 1.0960905e-10
+ voff = -0.1302643
+ ldif = 9e-8
+ wvsat = 0.0
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ lpclm = 4.03983e-8
+ wvth0 = 1.18629e-9
+ eta0 = -0.0004687502
+ pvag = 0.0
+ etab = 0.0010775371
+ vsat = 130812.52
+ wint = 5e-9
+ vth0 = -0.4245751
+ rdsw = 530.0
+ tcjswg = 0.0004130718
+ lint = 1.4999999e-8
+ wmax = 0.000900001
+ ags = 0.02
+ )

.model pch_ff_5 pmos (
+ level = 49
+ wa0 = -4.787191e-8
+ pscbe1 = 199999970.0
+ pscbe2 = 5e-7
+ ute = -0.8394966
+ lvth0 = 3.9543e-9
+ wk1 = 1.2456701e-8
+ wk2 = -5.940143e-9
+ wln = 1.0
+ wu0 = -1.2297032e-9
+ delta = 0.01
+ wua = 1.7543858e-16
+ wub = -6.530953e-25
+ wuc = -7.950096e-17
+ wwl = 0.0
+ wwn = 1.0
+ nqsmod = 0
+ xti = 3
+ version = 3.24
+ tpbswg = 0.001572025
+ noimod = 2
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ keta = 0.02600144
+ dsub = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ voff = -0.1274889
+ ldif = 9e-8
+ tcjsw = 0.0004130718
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ eta0 = 5e-5
+ pvoff = 0.0
+ capmod = 3
+ pvag = 0.0
+ etab = -5e-5
+ vsat = 149999.98
+ wint = 5e-9
+ vth0 = -0.41604359999999996
+ cdscb = 0.0
+ rdsw = 530.0
+ cdscd = 0.0
+ pnfactor = 0
+ peta0 = 4.7451600189666944e-17
+ wkt1 = 8.228274e-9
+ wkt2 = 1.4868883e-9
+ lint = 1.4999999e-8
+ wnfactor = 0.0
+ wmax = 9.991300540000001e-6
+ wketa = 6.301227e-9
+ wmin = 1.19130054e-6
+ pvth0 = 1.18629e-15
+ mobmod = 1
+ drout = 0.0
+ tpbsw = 0.001572025
+ lmax = 2.0001e-5
+ lmin = 1.0005259219000001e-5
+ cjswg = 4.00995e-10
+ a0 = 1.0509492
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ at = 10000.0
+ mjswg = 0.3683619
+ cf = 0
+ cj = 0.00106495
+ lnfactor = 3.9543e-9
+ ef = 1.064
+ k1 = 0.5362856
+ k2 = 0.03009115
+ k3 = 0.0
+ em = 30000000.0
+ js = 2.5e-7
+ ll = 0.0
+ mj = 0.4476
+ lw = 0.0
+ u0 = 0.0110455512
+ pb = 0.895226
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ wvoff = -1.0305298e-9
+ ua = 8.057326e-10
+ ub = 7.508071e-19
+ uc = -7.859605e-11
+ wub1 = 6.909715e-26
+ wuc1 = 3.0354498e-17
+ wl = 0.0
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -2.5259219000000002e-8
+ ww = 0.0
+ xw = 8.69946e-9
+ hdif = 2e-7
+ weta0 = 0
+ ags = 0.02
+ wute = 1.0600407e-7
+ mjsw = 0.3683619
+ wvsat = 0.0
+ wvth0 = 1.4056747999999999e-8
+ cit = -0.0001
+ dlc = 2e-9
+ nfactor = 1.0
+ k3b = 0.0
+ tcjswg = 0.0004130718
+ dwb = 0.0
+ dwg = 0.0
+ cdsc = 0.0
+ cgdo = 3.444e-10
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0010000004
+ cgso = 3.444e-10
+ pdiblcb = 0.01
+ jsw = 1.2e-12
+ kt1 = -0.231953
+ kt2 = -0.024488758
+ lk2 = -1.18629e-9
+ llc = -0.039
+ lln = -1
+ cjsw = 2.35695e-10
+ lu0 = 7.9086e-11
+ xpart = 1
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ binunit = 2
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ nlx = 0.0
+ pbswg = 0.895226
+ pu0 = 0.0
+ prt = 0
+ tnom = 25.0
+ lvoff = 1.5817200000000002e-9
+ rsh = 7.2
+ beta0 = 22.67827
+ toxm = 4.08e-9
+ tcj = 0.0009739001
+ ua1 = 1.224e-9
+ ub1 = -1.3998005e-18
+ uc1 = -7.633158e-12
+ leta0 = 4.745160018966694e-10
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ pbsw = 0.895226
+ pclm = 0.6000001
+ tpb = 0.001572025
+ tox = 4.02740781e-9
+ )

.model pch_ff_6 pmos (
+ level = 49
+ lub1 = 5.442727e-26
+ luc1 = 1.8276951e-17
+ wute = 1.0644106e-7
+ mjsw = 0.3683619
+ tcjsw = 0.0004130718
+ capmod = 3
+ lute = 9.664497e-8
+ pvoff = -4.403278e-15
+ nfactor = 1.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 4.7451600189666944e-17
+ mobmod = 1
+ cgdo = 3.444e-10
+ wketa = 7.084359e-9
+ pvth0 = -4.150182e-15
+ cgso = 3.444e-10
+ drout = 0.0
+ tpbsw = 0.001572025
+ ags = 0.02
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0004772728
+ pdiblcb = 0.01
+ lpscbe1 = 195.04262
+ cjswg = 4.00995e-10
+ cit = -0.0001
+ cjsw = 2.35695e-10
+ mjswg = 0.3683619
+ dlc = 2e-9
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ k3b = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ wvoff = -5.879894e-10
+ binunit = 2
+ tnom = 25.0
+ weta0 = 0
+ wvsat = 0.0
+ toxm = 4.08e-9
+ lpclm = 2.6005682e-7
+ wvth0 = 1.4593076e-8
+ la0 = 6.878132e-8
+ pbsw = 0.895226
+ tcjswg = 0.0004130718
+ pclm = 0.5738637
+ jsw = 1.2e-12
+ kt1 = -0.2303147
+ lk1 = 1.8184398e-8
+ kt2 = -0.024155809
+ lk2 = -6.466925e-9
+ llc = -0.039
+ lln = -1
+ lu0 = -1.2264377e-9
+ lua = -3.935608e-16
+ lub = 4.219459e-25
+ luc = 1.8883157e-17
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ pnfactor = 0
+ pa0 = 6.693222e-14
+ nlx = 0.0
+ wnfactor = 0.0
+ pk1 = 5.986243e-15
+ pk2 = -2.063307e-15
+ pu0 = 1.1543239e-16
+ prt = 0
+ pua = 3.1465633e-23
+ pub = 2.8088595e-31
+ puc = 9.8941e-24
+ version = 3.24
+ lketa = -1.2662711e-9
+ rsh = 7.2
+ pkt1 = 9.666697e-15
+ tcj = 0.0009739001
+ pkt2 = 2.4000725e-15
+ ua1 = 1.224e-9
+ keta = 0.026128704
+ ub1 = -1.4052706e-18
+ uc1 = -9.470036e-12
+ xpart = 1
+ tpb = 0.001572025
+ lnfactor = 3.9543e-9
+ tox = 4.02740781e-9
+ dsub = 0.0
+ wa0 = -5.459876e-8
+ ute = -0.8492097
+ wk1 = 1.185507e-8
+ wk2 = -5.732776e-9
+ pbswg = 0.895226
+ wln = 1.0
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ wu0 = -1.2413044999999998e-9
+ wua = 1.7227619e-16
+ wub = -6.81325e-25
+ wuc = -8.049533e-17
+ wwl = 0.0
+ wwn = 1.0
+ a0 = 1.0440365
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ lvoff = 1.1335760000000018e-10
+ xti = 3
+ at = 10000.0
+ cf = 0
+ lpdiblc2 = 5.201137e-9
+ cj = 0.00106495
+ voff = -0.1273414
+ ef = 1.064
+ k1 = 0.534458
+ k2 = 0.03062187
+ k3 = 0.0
+ em = 30000000.0
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ ldif = 9e-8
+ beta0 = 22.67827
+ js = 2.5e-7
+ ll = 0.0
+ mj = 0.4476
+ lw = 0.0
+ u0 = 0.0111767602
+ pb = 0.895226
+ kt1l = 0.0
+ w0 = 0.0
+ prwb = 0.0
+ rd = 0
+ pub1 = -6.397619e-32
+ prwg = 0.0
+ leta0 = 4.745160018966694e-10
+ puc1 = 2.6178952e-23
+ rs = 0
+ ua = 8.452865e-10
+ ub = 7.084005e-19
+ uc = -8.049386e-11
+ pscbe1 = 180397700.0
+ pscbe2 = 5e-7
+ wl = 0.0
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -2.5259219000000002e-8
+ ww = 0.0
+ xw = 8.69946e-9
+ eta0 = 5e-5
+ lvsat = -0.013002842
+ pvag = 0.0
+ etab = -5e-5
+ vsat = 151306.8
+ lvth0 = -2.0325569e-8
+ wint = 5e-9
+ pute = -4.348101e-15
+ vth0 = -0.41360349999999996
+ nqsmod = 0
+ rdsw = 530.0
+ tpbswg = 0.001572025
+ delta = 0.01
+ wkt1 = 7.256747e-9
+ wkt2 = 1.245675e-9
+ noimod = 2
+ lint = 1.4999999e-8
+ wmax = 9.991300540000001e-6
+ wmin = 1.19130054e-6
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ lkt1 = -1.6300865e-8
+ lkt2 = -3.312836e-9
+ lmax = 1.0005259219000001e-5
+ lmin = 1.205259219e-6
+ pketa = -7.792167e-15
+ wub1 = 7.552692e-26
+ wuc1 = 2.7723443e-17
+ hdif = 2e-7
+ )

.model pch_ff_7 pmos (
+ level = 49
+ mjswg = 0.3683619
+ jsw = 1.2e-12
+ kt1 = -0.2459144
+ lk1 = 8.371453e-9
+ kt2 = -0.027846618
+ lk2 = -4.402144e-9
+ dsub = 0.0
+ llc = -0.039
+ lln = -1
+ lu0 = -2.666366e-10
+ wvoff = -7.866491e-9
+ lua = 3.0792715e-17
+ lub = -1.9665828e-25
+ luc = -3.700045e-17
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ wcit = -1.788104e-11
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ pa0 = -1.2519753e-13
+ nlx = 0.0
+ weta0 = 0
+ pk1 = 4.753178e-14
+ pk2 = -1.4849934e-14
+ lcit = 2.2196864e-10
+ voff = -0.1274479
+ pu0 = -6.201592e-16
+ wvsat = 0.0
+ ldif = 9e-8
+ tcjswg = 0.0004130718
+ prt = 0
+ pua = -3.495584e-22
+ pub = 3.345938e-31
+ puc = 4.854297e-23
+ lpclm = 1.4785702e-7
+ wvth0 = 1.1317e-8
+ kt1l = 0.0
+ prwb = 0.0
+ pub1 = -1.382964e-31
+ prwg = 0.0
+ puc1 = -5.043768e-23
+ eta0 = 1.7857139e-5
+ rsh = 7.2
+ tcj = 0.0009739001
+ ua1 = 1.224e-9
+ pvag = 0.0
+ ub1 = -1.3967723e-18
+ etab = -1.7857139e-5
+ uc1 = -2.3838735e-11
+ vsat = 146428.53
+ wint = 5e-9
+ pute = 2.0900147e-14
+ tpb = 0.001572025
+ tox = 4.02740781e-9
+ vth0 = -0.4290361
+ wa0 = 1.1247056e-7
+ rdsw = 530.0
+ ute = -0.7951261
+ wkt1 = 1.6218328e-8
+ wkt2 = 2.9642964e-9
+ wk1 = -2.4271484e-8
+ wk2 = 5.386031e-9
+ lint = 1.4999999e-8
+ wmax = 9.991300540000001e-6
+ wln = 1.0
+ wu0 = -6.016596e-10
+ wmin = 1.19130054e-6
+ wua = 5.036014e-16
+ wub = -7.280275e-25
+ wuc = -1.1410304e-16
+ lkt1 = 1.6387112e-9
+ lkt2 = 9.315946e-10
+ wwl = 0.0
+ wwn = 1.0
+ xti = 3
+ lmax = 1.205259219e-6
+ lketa = -8.380984e-9
+ lmin = 5.052592189999999e-7
+ xpart = 1
+ wub1 = 1.4015321e-25
+ pbswg = 0.895226
+ wuc1 = 9.434661e-17
+ hdif = 2e-7
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ lvoff = 2.3584050000000025e-10
+ lub1 = 4.46543e-26
+ luc1 = 3.480094e-17
+ wute = 8.448607e-8
+ mjsw = 0.3683619
+ pscbe1 = 349999900.0
+ pscbe2 = 5e-7
+ beta0 = 22.67827
+ leta0 = 5.114802918966694e-10
+ lute = 3.444881e-8
+ letab = -3.696429e-11
+ lvsat = -0.007392833
+ lvth0 = -2.5780870000000004e-9
+ nqsmod = 0
+ tpbswg = 0.001572025
+ noimod = 2
+ cdsc = 0.0
+ pnfactor = 0
+ delta = 0.01
+ wnfactor = 0.0
+ cgdo = 3.444e-10
+ nfactor = 1.0
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ cgso = 3.444e-10
+ cjsw = 2.35695e-10
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0017857144
+ lnfactor = 3.9543e-9
+ pdiblcb = 0.01
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ pketa = 2.2253538e-15
+ tnom = 25.0
+ binunit = 2
+ capmod = 3
+ lpdiblc2 = 3.696428e-9
+ tcjsw = 0.0004130718
+ toxm = 4.08e-9
+ ags = 0.02
+ pcit = 2.0563189e-17
+ pbsw = 0.895226
+ pclm = 0.6714287
+ pvoff = 3.966999e-15
+ cit = -0.0002930162
+ a0 = 0.9932752
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ at = 10000.0
+ mobmod = 1
+ cf = 0
+ dlc = 2e-9
+ cj = 0.00106495
+ ef = 1.064
+ k1 = 0.542991
+ k2 = 0.0288264
+ k3 = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ em = 30000000.0
+ peta0 = 4.7451600189666944e-17
+ k3b = 0.0
+ js = 2.5e-7
+ ll = 0.0
+ mj = 0.4476
+ lw = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ u0 = 0.0103421492
+ pb = 0.895226
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ua = 4.762835e-10
+ ub = 1.2463172e-18
+ uc = -3.189942e-11
+ wl = 0.0
+ wr = 1.0
+ xj = 1.7000001e-7
+ wketa = -1.6265284e-9
+ xl = -2.5259219000000002e-8
+ ww = 0.0
+ xw = 8.69946e-9
+ pvth0 = -3.826928e-16
+ drout = 0.0
+ tpbsw = 0.001572025
+ pkt1 = -6.391237e-16
+ pkt2 = 4.236579e-16
+ keta = 0.03231541
+ cjswg = 4.00995e-10
+ version = 3.24
+ la0 = 1.2715688e-7
+ )

.model pch_ff_8 pmos (
+ level = 49
+ cgso = 3.444e-10
+ nfactor = 1.0
+ a0 = 1.2640158
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ lketa = -5.872592e-10
+ at = 10000.0
+ cf = 0
+ cj = 0.00106495
+ ef = 1.064
+ k1 = 0.5203763
+ k2 = 0.036403239999999996
+ k3 = 0.0
+ em = 30000000.0
+ pcdscd = -7.408954e-18
+ js = 2.5e-7
+ ll = 0.0
+ mj = 0.4476
+ lw = 0.0
+ u0 = 0.0098511212
+ pb = 0.895226
+ xpart = 1
+ w0 = 0.0
+ rd = 0
+ cjsw = 2.35695e-10
+ rs = 0
+ ua = 9.357863e-10
+ ub = 5.091257e-19
+ uc = -1.5731644e-10
+ wl = 0.0
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -2.5259219000000002e-8
+ ww = 0.0
+ xw = 8.69946e-9
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.007987866
+ pbswg = 0.895226
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ pdiblcb = 0.01
+ pscbe1 = 350000000.0
+ pscbe2 = 5e-7
+ lvoff = 1.7452549500000003e-9
+ tnom = 25.0
+ pags = -6.875222e-16
+ beta0 = 22.67827
+ toxm = 4.08e-9
+ binunit = 2
+ leta0 = 7.304535218966694e-10
+ letab = -5.545772e-10
+ nqsmod = 0
+ pcit = -7.907631e-17
+ pbsw = 0.895226
+ pclm = 0.9107697
+ tpbswg = 0.001572025
+ lvsat = -0.0003656271
+ noimod = 2
+ lvth0 = -4.173726e-9
+ ppclm = 2.4445072e-15
+ delta = 0.01
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ lcdscd = 3.730414e-11
+ pkt1 = -1.8229216e-15
+ pkt2 = -1.2254391e-15
+ keta = 0.014996022
+ ags = 0.019847063
+ wags = 1.5278273e-9
+ dsub = 0.0
+ version = 3.24
+ cit = -6.09184e-5
+ pketa = -2.4325694e-15
+ dlc = 2e-9
+ lags = 6.882101e-11
+ wcit = 2.0354016e-10
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ k3b = 0.0
+ capmod = 3
+ dwb = 0.0
+ dwg = 0.0
+ wpclm = -5.432238e-9
+ lcit = 1.1752459e-10
+ voff = -0.1308021
+ tcjsw = 0.0004130718
+ ldif = 9e-8
+ kt1l = 0.0
+ prwb = 0.0
+ pub1 = 2.7781507e-32
+ prwg = 0.0
+ puc1 = 8.113434e-24
+ pvoff = -1.9905158e-15
+ eta0 = -0.0004687502
+ mobmod = 1
+ pvag = 0.0
+ etab = 0.0011323938
+ la0 = 5.323636e-9
+ vsat = 130812.52
+ wint = 5e-9
+ pute = 9.798417e-15
+ jsw = 1.2e-12
+ kt1 = -0.2367561
+ lk1 = 1.854804e-8
+ kt2 = -0.025532207
+ lk2 = -7.811716e-9
+ vth0 = -0.4254902
+ cdscb = 0.0
+ cdscd = -8.289813e-5
+ pnfactor = 0
+ peta0 = 4.7451600189666944e-17
+ llc = -0.039
+ rdsw = 530.0
+ lln = -1
+ lu0 = -4.5673330000000005e-11
+ petab = 2.4660761e-16
+ wnfactor = 0.0
+ wkt1 = 1.8848993e-8
+ wkt2 = 6.628956e-9
+ lua = -1.759835e-16
+ lub = 1.3507784e-25
+ luc = 1.9437196e-17
+ lint = 1.4999999e-8
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ wmax = 9.991300540000001e-6
+ wketa = 8.724413e-9
+ pvth0 = 6.215440000000003e-17
+ pa0 = 1.0862038e-13
+ nlx = 0.0
+ wmin = 1.19130054e-6
+ drout = 0.0
+ lkt1 = -2.4825255e-9
+ lkt2 = -1.0989117e-10
+ tpbsw = 0.001572025
+ pk1 = -1.7383759e-14
+ pk2 = 7.484627e-15
+ lmax = 5.052592189999999e-7
+ pu0 = 2.5785697e-16
+ lmin = 1.8e-7
+ ppdiblc2 = 8.594017e-17
+ prt = 0
+ pua = 1.5976873e-22
+ pub = -1.3085017e-31
+ puc = -9.356197e-24
+ cjswg = 4.00995e-10
+ wpdiblc2 = -1.9097854e-10
+ mjswg = 0.3683619
+ lnfactor = 3.9543e-9
+ rsh = 7.2
+ tcj = 0.0009739001
+ ua1 = 1.224e-9
+ ub1 = -1.3554493e-18
+ uc1 = 7.051652e-11
+ wvoff = 5.372431e-9
+ tpb = 0.001572025
+ tox = 4.02740781e-9
+ wub1 = -2.2890885e-25
+ wuc1 = -3.576699e-17
+ wa0 = -4.071248e-7
+ hdif = 2e-7
+ ute = -0.7199521
+ wk1 = 1.1998529e-7
+ wk2 = -4.424634e-8
+ weta0 = 0
+ tcjswg = 0.0004130718
+ lub1 = 2.6058948e-26
+ luc1 = -7.658915e-18
+ wln = 1.0
+ wetab = -5.480169e-10
+ lpdiblc2 = 9.0546e-10
+ wu0 = -2.5528067e-9
+ wute = 1.0915658e-7
+ mjsw = 0.3683619
+ wvsat = 0.0
+ wua = -6.282368e-16
+ wub = 3.0629255e-25
+ wuc = 1.4561782e-17
+ wwl = 0.0
+ wwn = 1.0
+ lpclm = 4.015361e-8
+ wvth0 = 1.0328453999999999e-8
+ xti = 3
+ lute = 6.205235e-10
+ cdsc = 0.0
+ wcdscd = 1.6464351e-11
+ cgdo = 3.444e-10
+ )

.model pch_ff_9 pmos (
+ level = 49
+ pvag = 0.0
+ etab = -5e-5
+ lvth0 = 3.9543e-9
+ ags = 0.02
+ vsat = 149999.98
+ wint = 5e-9
+ vth0 = -0.40491299999999997
+ delta = 0.01
+ rdsw = 530.0
+ cit = -0.0001
+ wkt1 = 6.74333e-9
+ wkt2 = 1.2948118e-10
+ lint = 1.4999999e-8
+ dlc = 2e-9
+ wmax = 1.19130054e-6
+ dvt0w = 0.0
+ k3b = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ wmin = 4.9130054e-7
+ dwb = 0.0
+ dwg = 0.0
+ lmax = 2.0001e-5
+ lmin = 1.0005259219000001e-5
+ capmod = 3
+ a0 = 0.9810578
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ jsw = 1.2e-12
+ kt1 = -0.2307052
+ kt2 = -0.02334808
+ lk2 = -1.18629e-9
+ wub1 = 3.495163e-26
+ wuc1 = 1.9335648e-17
+ at = 10000.0
+ cf = 0
+ cj = 0.00106495
+ ef = 1.064
+ k1 = 0.5449055
+ k2 = 0.02831336
+ k3 = 0.0
+ em = 30000000.0
+ llc = -0.039
+ lln = -1
+ lu0 = 7.9086e-11
+ hdif = 2e-7
+ js = 2.5e-7
+ ll = 0.0
+ mj = 0.4476
+ lw = 0.0
+ u0 = 0.0101875252
+ nch = 3.9e+17
+ pb = 0.895226
+ w0 = 0.0
+ rd = 0
+ lwl = 0.0
+ lwn = 1.0
+ rs = 0
+ ua = 1.0698959e-9
+ ub = 3.0837888e-19
+ uc = -1.1659398e-10
+ wl = 0.0
+ wute = -2.7886795e-9
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -2.5259219000000002e-8
+ ww = 0.0
+ xw = 8.69946e-9
+ mjsw = 0.3683619
+ nlx = 0.0
+ tcjsw = 0.0004130718
+ mobmod = 1
+ pu0 = 0.0
+ pvoff = 0.0
+ prt = 0
+ rsh = 7.2
+ cdscb = 0.0
+ cdscd = 0.0
+ tcj = 0.0009739001
+ peta0 = 4.7451600189666944e-17
+ cdsc = 0.0
+ ua1 = 1.224e-9
+ ub1 = -1.3711068e-18
+ uc1 = 1.6263793e-12
+ tpb = 0.001572025
+ tox = 4.02740781e-9
+ cgdo = 3.444e-10
+ wketa = -1.0458587e-9
+ wa0 = 3.529885e-8
+ pvth0 = 1.18629e-15
+ drout = 0.0
+ ute = -0.7480742
+ wk1 = 2.1990281e-9
+ cgso = 3.444e-10
+ wk2 = -3.824582e-9
+ tpbsw = 0.001572025
+ wln = 1.0
+ wu0 = -2.086521e-10
+ wua = -1.3891575e-16
+ wub = -1.2660565e-25
+ wuc = -3.428342e-17
+ wwl = 0.0
+ wwn = 1.0
+ cjswg = 4.00995e-10
+ nfactor = 1.0
+ xti = 3
+ cjsw = 2.35695e-10
+ mjswg = 0.3683619
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ wvoff = -4.105241e-10
+ tcjswg = 0.0004130718
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0009999998
+ weta0 = 0
+ tnom = 25.0
+ pdiblcb = 0.01
+ wvsat = 0.0
+ wvth0 = 8.112289000000001e-10
+ toxm = 4.08e-9
+ pbsw = 0.895226
+ pclm = 0.6
+ binunit = 2
+ pnfactor = 0
+ wnfactor = 0.0
+ keta = 0.03217546
+ xpart = 1
+ lnfactor = 3.9543e-9
+ alpha0 = 0.0
+ dsub = 0.0
+ alpha1 = 6.8730453846
+ pbswg = 0.895226
+ pscbe1 = 199999970.0
+ pscbe2 = 5e-7
+ dvt0 = 0.0
+ version = 3.24
+ dvt1 = 0.0
+ dvt2 = 0.0
+ lvoff = 1.5817200000000002e-9
+ voff = -0.12801
+ beta0 = 22.67827
+ nqsmod = 0
+ ldif = 9e-8
+ tpbswg = 0.001572025
+ noimod = 2
+ leta0 = 4.745160018966694e-10
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ eta0 = 5e-5
+ )

.model pch_ff_10 pmos (
+ level = 49
+ dsub = 0.0
+ wk1 = 1.7598129e-9
+ wk2 = -3.600003e-9
+ wln = 1.0
+ wu0 = -1.7835274000000001e-10
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ wua = -1.6455617e-16
+ wub = -7.150721e-26
+ wuc = -2.8652769e-17
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ wwl = 0.0
+ wwn = 1.0
+ xti = 3
+ pscbe1 = 180397680.0
+ pscbe2 = 5e-7
+ voff = -0.1269095
+ ldif = 9e-8
+ nfactor = 1.0
+ kt1l = 0.0
+ prwb = 0.0
+ pub1 = -8.629597e-32
+ prwg = 0.0
+ puc1 = 1.5034668e-23
+ nqsmod = 0
+ tpbswg = 0.001572025
+ lketa = -6.417587e-9
+ eta0 = 5e-5
+ noimod = 2
+ pvag = 0.0
+ etab = -5e-5
+ vsat = 151306.8
+ wint = 5e-9
+ pute = 3.909688e-14
+ xpart = 1
+ vth0 = -0.40084529999999996
+ rdsw = 530.0
+ wkt1 = 6.495125e-9
+ wkt2 = 2.3726165e-10
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0004772722
+ lint = 1.4999999e-8
+ pdiblcb = 0.01
+ lpscbe1 = 195.04263
+ wmax = 1.19130054e-6
+ pbswg = 0.895226
+ wmin = 4.9130054e-7
+ lkt1 = -1.0252924e-8
+ lkt2 = -3.947785e-10
+ lmax = 1.0005259219000001e-5
+ lvoff = -9.367244999999999e-9
+ lmin = 1.205259219e-6
+ beta0 = 22.67827
+ binunit = 2
+ leta0 = 4.745160018966694e-10
+ lvsat = -0.013002842
+ lvth0 = -3.651863e-8
+ wub1 = 4.362458e-26
+ wuc1 = 1.7824627e-17
+ capmod = 3
+ hdif = 2e-7
+ delta = 0.01
+ lub1 = 7.318341e-26
+ luc1 = 2.7641896e-17
+ pnfactor = 0
+ wute = -6.718015e-9
+ mjsw = 0.3683619
+ wnfactor = 0.0
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ lute = 6.013659e-8
+ mobmod = 1
+ cdsc = 0.0
+ version = 3.24
+ lnfactor = 3.9543e-9
+ pketa = -1.6621007e-15
+ cgdo = 3.444e-10
+ ags = 0.02
+ cgso = 3.444e-10
+ cit = -0.0001
+ tcjsw = 0.0004130718
+ dlc = 2e-9
+ lpdiblc2 = 5.201137e-9
+ cjsw = 2.35695e-10
+ k3b = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ pvoff = 6.87864e-15
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 4.7451600189666944e-17
+ tcjswg = 0.0004130718
+ tnom = 25.0
+ wketa = -8.788133e-10
+ pvth0 = 1.511956e-14
+ la0 = 1.2176828e-7
+ drout = 0.0
+ toxm = 4.08e-9
+ jsw = 1.2e-12
+ kt1 = -0.2296747
+ lk1 = 1.9542425e-8
+ kt2 = -0.023308404
+ lk2 = -6.323008999999999e-9
+ tpbsw = 0.001572025
+ pbsw = 0.895226
+ llc = -0.039
+ pclm = 0.5738636
+ lln = -1
+ lu0 = -8.760922000000001e-10
+ lua = -5.815077e-16
+ lub = 1.1186816e-24
+ luc = 7.427734e-17
+ nch = 3.9e+17
+ a0 = 0.9688198
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ lwl = 0.0
+ lwn = 1.0
+ cjswg = 4.00995e-10
+ at = 10000.0
+ cf = 0
+ cj = 0.00106495
+ pa0 = 3.87773e-15
+ nlx = 0.0
+ ef = 1.064
+ k1 = 0.5429414
+ k2 = 0.028829620000000004
+ k3 = 0.0
+ em = 30000000.0
+ mjswg = 0.3683619
+ js = 2.5e-7
+ ll = 0.0
+ mj = 0.4476
+ lw = 0.0
+ pk1 = 4.370194e-15
+ pk2 = -2.2345663e-15
+ u0 = 0.0102835232
+ pb = 0.895226
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ua = 1.1283389e-9
+ ub = 1.9594849e-19
+ uc = -1.2405904e-10
+ wvoff = -1.1018445e-9
+ wl = 0.0
+ pu0 = -3.0147877e-16
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -2.5259219000000002e-8
+ ww = 0.0
+ xw = 8.69946e-9
+ prt = 0
+ pua = 2.5512236e-22
+ pub = -5.482294e-31
+ puc = -5.602498e-23
+ weta0 = 0
+ rsh = 7.2
+ tcj = 0.0009739001
+ ua1 = 1.224e-9
+ ub1 = -1.3784619e-18
+ uc1 = -1.1517035e-12
+ wvsat = 0.0
+ pkt1 = 2.469645e-15
+ pkt2 = -1.0724159e-15
+ keta = 0.03282044
+ tpb = 0.001572025
+ tox = 4.02740781e-9
+ lpclm = 2.6005682e-7
+ wvth0 = -5.891015e-10
+ wa0 = 3.490912e-8
+ ute = -0.754118
+ )

.model pch_ff_11 pmos (
+ level = 49
+ cgso = 3.444e-10
+ a0 = 1.1936638
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ lvoff = 6.818931000000001e-9
+ at = 10000.0
+ cf = 0
+ cj = 0.00106495
+ ef = 1.064
+ k1 = 0.4715038
+ k2 = 0.05425073
+ k3 = 0.0
+ em = 30000000.0
+ js = 2.5e-7
+ ll = 0.0
+ mj = 0.4476
+ lw = 0.0
+ beta0 = 22.67827
+ u0 = 0.0107824642
+ pb = 0.895226
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ua = 1.036115e-9
+ ub = 1.0523674e-18
+ uc = -7.205117e-11
+ cjsw = 2.35695e-10
+ leta0 = 5.114802618966694e-10
+ wl = 0.0
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -2.5259219000000002e-8
+ ww = 0.0
+ xw = 8.69946e-9
+ letab = -3.696426e-11
+ lvsat = -0.007392855
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ capmod = 3
+ lvth0 = 3.9159799999999995e-10
+ delta = 0.01
+ tnom = 25.0
+ ags = 0.02
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ toxm = 4.08e-9
+ mobmod = 1
+ pcit = -1.0851648e-17
+ pbsw = 0.895226
+ pclm = 0.6714286
+ cit = -0.00031597191
+ dlc = 2e-9
+ k3b = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ pketa = 4.024799e-15
+ la0 = -1.3680231e-7
+ pkt1 = -6.051915e-15
+ pkt2 = -1.4802061e-15
+ tcjsw = 0.0004130718
+ keta = 0.03584265
+ jsw = 1.2e-12
+ kt1 = -0.2439705
+ lk1 = 1.0169572e-7
+ kt2 = -0.025852976
+ lk2 = -3.555729e-8
+ llc = -0.039
+ lln = -1
+ lu0 = -1.4498735e-9
+ dsub = 0.0
+ pvoff = -3.866879e-15
+ lua = -4.754501e-16
+ lub = 1.337998e-25
+ luc = 1.4468274e-17
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ pa0 = 1.8891395e-13
+ nlx = 0.0
+ tcjswg = 0.0004130718
+ wcit = 9.436221e-12
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ pk1 = -6.35241e-14
+ pk2 = 2.2224691e-14
+ peta0 = 4.7451600189666944e-17
+ pu0 = 7.878928e-16
+ pnfactor = 0
+ prt = 0
+ lcit = 2.4836766e-10
+ pua = 2.5287059e-22
+ pub = -5.865131e-32
+ puc = -1.2704817e-23
+ wketa = -5.823942e-9
+ voff = -0.1409845
+ pvth0 = -3.9166180000000005e-15
+ wnfactor = 0.0
+ ldif = 9e-8
+ drout = 0.0
+ kt1l = 0.0
+ tpbsw = 0.001572025
+ prwb = 0.0
+ pub1 = 4.97241e-32
+ prwg = 0.0
+ rsh = 7.2
+ puc1 = 1.7282469e-23
+ tcj = 0.0009739001
+ ua1 = 1.224e-9
+ ub1 = -1.2162624e-18
+ uc1 = 4.210797e-11
+ eta0 = 1.7857154e-5
+ nfactor = 1.0
+ pvag = 0.0
+ etab = -1.7857154e-5
+ tpb = 0.001572025
+ tox = 4.02740781e-9
+ cjswg = 4.00995e-10
+ vsat = 146428.56
+ wa0 = -1.2599192e-7
+ wint = 5e-9
+ pute = -5.928695e-14
+ mjswg = 0.3683619
+ vth0 = -0.43294119999999997
+ ute = -0.7903757
+ wk1 = 6.079834e-8
+ wk2 = -2.4868919e-8
+ rdsw = 530.0
+ wln = 1.0
+ wkt1 = 1.3905176e-8
+ wkt2 = 5.918618e-10
+ lnfactor = 3.9543e-9
+ wu0 = -1.1256324e-9
+ lint = 1.4999999e-8
+ wvoff = 8.242083e-9
+ wua = -1.625981e-16
+ wmax = 1.19130054e-6
+ wub = -4.972273e-25
+ wuc = -6.632247e-17
+ wwl = 0.0
+ wwn = 1.0
+ wmin = 4.9130054e-7
+ xti = 3
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0017857137
+ lkt1 = 6.187276e-9
+ lkt2 = 2.5314804e-9
+ pdiblcb = 0.01
+ weta0 = 0
+ lmax = 1.205259219e-6
+ lmin = 5.052592189999999e-7
+ wvsat = 0.0
+ lpclm = 1.4785714e-7
+ wvth0 = 1.5964097e-8
+ lpdiblc2 = 3.696429e-9
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ binunit = 2
+ pscbe1 = 349999900.0
+ pscbe2 = 5e-7
+ wub1 = -7.465372e-26
+ wuc1 = 1.5870021e-17
+ hdif = 2e-7
+ lub1 = -1.133461e-25
+ luc1 = -2.2106738e-17
+ wute = 7.883313e-8
+ mjsw = 0.3683619
+ nqsmod = 0
+ tpbswg = 0.001572025
+ noimod = 2
+ lute = 1.0183292e-7
+ lketa = -9.893122e-9
+ xpart = 1
+ cdsc = 0.0
+ cgdo = 3.444e-10
+ pbswg = 0.895226
+ version = 3.24
+ )

.model pch_ff_12 pmos (
+ level = 49
+ wint = 5e-9
+ llc = -0.039
+ pute = 1.3160581e-15
+ lln = -1
+ lu0 = 2.9107207000000003e-10
+ vth0 = -0.42263
+ nfactor = 1.0
+ lua = 2.3815556e-17
+ lub = -3.425063e-26
+ luc = 8.803578e-18
+ nch = 3.9e+17
+ rdsw = 530.0
+ lwl = 0.0
+ lwn = 1.0
+ pketa = -9.609158e-16
+ wkt1 = 2.7434011e-10
+ wkt2 = -6.113567e-9
+ lint = 1.4999999e-8
+ pa0 = -8.476619e-14
+ nlx = 0.0
+ wmax = 1.19130054e-6
+ pk1 = 1.5213101e-14
+ pk2 = -6.235986e-15
+ wmin = 4.9130054e-7
+ lkt1 = -4.083267e-9
+ lkt2 = -2.4314675e-9
+ wpclm = 5.671285e-8
+ pu0 = -1.4287007e-16
+ lmax = 5.052592189999999e-7
+ prt = 0
+ pua = -7.799214e-23
+ pub = 7.065072e-32
+ puc = 3.297807e-24
+ lmin = 1.8e-7
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.009150297
+ tcjsw = 0.0004130718
+ pdiblcb = 0.01
+ rsh = 7.2
+ tcj = 0.0009739001
+ ua1 = 1.224e-9
+ ub1 = -1.6175756e-18
+ uc1 = -2.2818641e-11
+ pvoff = -1.4343533e-15
+ tcjswg = 0.0004130718
+ tpb = 0.001572025
+ tox = 4.02740781e-9
+ a0 = 0.5166956
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ wa0 = 4.821862e-7
+ at = 10000.0
+ cf = 0
+ cj = 0.00106495
+ wub1 = 8.30214e-26
+ ute = -0.5812994
+ wuc1 = 7.530186e-17
+ ef = 1.064
+ k1 = 0.7171482
+ k2 = -0.033028159
+ k3 = 0.0
+ em = 30000000.0
+ wk1 = -1.1417325e-7
+ wk2 = 3.837703e-8
+ binunit = 2
+ cdscb = 0.0
+ cdscd = -5.200001e-5
+ peta0 = 4.7451600189666944e-17
+ js = 2.5e-7
+ ll = 0.0
+ mj = 0.4476
+ hdif = 2e-7
+ lw = 0.0
+ u0 = 0.0069136952
+ wln = 1.0
+ pb = 0.895226
+ w0 = 0.0
+ wu0 = 9.427299e-10
+ rd = 0
+ rs = 0
+ ua = -7.336427e-11
+ ub = 1.4258127e-18
+ uc = -5.946296e-11
+ lub1 = 6.724484e-26
+ wua = 5.726523e-16
+ wub = -7.845651e-25
+ wuc = -1.0188386e-16
+ wl = 0.0
+ luc1 = 7.110234e-18
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -2.5259219000000002e-8
+ ww = 0.0
+ xw = 8.69946e-9
+ wwl = 0.0
+ wwn = 1.0
+ wute = -5.584022e-8
+ wketa = 5.255423e-9
+ mjsw = 0.3683619
+ pvth0 = 1.5103980000000002e-16
+ xti = 3
+ drout = 0.0
+ tpbsw = 0.001572025
+ lute = 7.748556e-9
+ wcdscd = -2.0304376e-11
+ cjswg = 4.00995e-10
+ mjswg = 0.3683619
+ cdsc = 0.0
+ wvoff = 2.8364715e-9
+ cgdo = 3.444e-10
+ pcdscd = 9.13697e-18
+ cgso = 3.444e-10
+ weta0 = 0
+ version = 3.24
+ wvsat = 0.0
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ lpclm = 6.365384e-8
+ wvth0 = 6.924854999999999e-9
+ cjsw = 2.35695e-10
+ pscbe1 = 350000000.0
+ pscbe2 = 5e-7
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ nqsmod = 0
+ tpbswg = 0.001572025
+ tnom = 25.0
+ pnfactor = 0
+ noimod = 2
+ pags = -5.667374e-15
+ wnfactor = 0.0
+ toxm = 4.08e-9
+ pcit = 2.6834248e-18
+ pbsw = 0.895226
+ lketa = -1.8239428e-9
+ pclm = 0.858547
+ xpart = 1
+ ppdiblc2 = 7.08422e-16
+ wpdiblc2 = -1.5742713e-9
+ lnfactor = 3.9543e-9
+ pbswg = 0.895226
+ lcdscd = 2.3400004e-11
+ lvoff = 1.2778913700000001e-9
+ ags = 0.010547621
+ beta0 = 22.67827
+ pkt1 = 8.196091e-17
+ pkt2 = 1.5372367e-15
+ keta = 0.01791114
+ lpdiblc2 = 3.823661e-10
+ leta0 = 7.304534718966694e-10
+ capmod = 3
+ letab = -3.473438e-10
+ cit = 0.00012746976
+ wags = 1.2594167e-8
+ lvsat = -0.0003656142
+ dsub = 0.0
+ dlc = 2e-9
+ lvth0 = -4.248419000000001e-9
+ k3b = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ lags = 4.253569e-9
+ wcit = -2.0641719e-11
+ ppclm = -2.5520774e-14
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ delta = 0.01
+ mobmod = 1
+ lcit = 4.881893e-11
+ voff = -0.1286711
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ ldif = 9e-8
+ kt1l = 0.0
+ prwb = 0.0
+ pub1 = -2.1229706e-32
+ prwg = 0.0
+ puc1 = -9.461855e-24
+ la0 = 1.6783336e-7
+ eta0 = -0.00046875
+ pvag = 0.0
+ jsw = 1.2e-12
+ etab = 0.0006718753
+ kt1 = -0.2211471
+ lk1 = -8.844278e-9
+ kt2 = -0.014824204
+ lk2 = 3.718209e-9
+ vsat = 130812.46
+ )

.model pch_ff_13 pmos (
+ level = 49
+ wketa = -6.403492e-9
+ pvth0 = 1.18629e-15
+ drout = 0.0
+ toxm = 4.08e-9
+ tpbsw = 0.001572025
+ pbsw = 0.895226
+ pclm = 0.5999999
+ cjswg = 4.00995e-10
+ mjswg = 0.3683619
+ wvoff = -1.320298e-9
+ weta0 = 0
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ wvsat = 0.0
+ keta = 0.04310941
+ pscbe1 = 199999970.0
+ pscbe2 = 5e-7
+ wvth0 = 1.0526903e-8
+ dsub = 0.0
+ nqsmod = 0
+ tpbswg = 0.001572025
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ noimod = 2
+ voff = -0.1261533
+ ldif = 9e-8
+ a0 = 0.8704194
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ at = 10000.0
+ cf = 0
+ cj = 0.00106495
+ ef = 1.064
+ k1 = 0.5421249
+ k2 = 0.0301404
+ k3 = 0.0
+ em = 30000000.0
+ ags = 0.02
+ eta0 = 5e-5
+ js = 2.5e-7
+ ll = 0.0
+ mj = 0.4476
+ lw = 0.0
+ pvag = 0.0
+ etab = -5e-5
+ u0 = 0.009803694200000001
+ pb = 0.895226
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ vsat = 149999.98
+ xpart = 1
+ ua = 1.2584637e-9
+ ub = 4.999999e-20
+ uc = -1.6065008e-10
+ wint = 5e-9
+ wl = 0.0
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -2.5259219000000002e-8
+ ww = 0.0
+ xw = 8.69946e-9
+ cit = -0.0001
+ vth0 = -0.4247409
+ rdsw = 530.0
+ dlc = 2e-9
+ wkt1 = 3.830554e-9
+ wkt2 = 1.9527771e-9
+ k3b = 0.0
+ lint = 1.4999999e-8
+ pbswg = 0.895226
+ dwb = 0.0
+ wmax = 4.9130054e-7
+ dwg = 0.0
+ nfactor = 1.0
+ wmin = 2.2e-7
+ lvoff = 1.5817200000000002e-9
+ lmax = 2.0001e-5
+ lmin = 1.0005259219000001e-5
+ capmod = 3
+ beta0 = 22.67827
+ leta0 = 4.745160018966694e-10
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.001
+ pdiblcb = 0.01
+ jsw = 1.2e-12
+ kt1 = -0.2247607
+ kt2 = -0.027069092
+ lk2 = -1.18629e-9
+ lvth0 = 3.9543e-9
+ llc = -0.039
+ lln = -1
+ lu0 = 7.9086e-11
+ wub1 = 2.1644123e-27
+ wuc1 = -1.2526765e-17
+ nch = 3.9e+17
+ mobmod = 1
+ lwl = 0.0
+ lwn = 1.0
+ delta = 0.01
+ hdif = 2e-7
+ nlx = 0.0
+ pnfactor = 0
+ binunit = 2
+ wute = 6.898109e-9
+ mjsw = 0.3683619
+ wnfactor = 0.0
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ pu0 = 0.0
+ prt = 0
+ rsh = 7.2
+ tcj = 0.0009739001
+ ua1 = 1.224e-9
+ ub1 = -1.3041941e-18
+ uc1 = 6.665171e-11
+ cdsc = 0.0
+ tpb = 0.001572025
+ tox = 4.02740781e-9
+ wa0 = 8.951166e-8
+ lnfactor = 3.9543e-9
+ cgdo = 3.444e-10
+ ute = -0.7678431
+ wk1 = 3.561511e-9
+ wk2 = -4.719829e-9
+ wln = 1.0
+ cgso = 3.444e-10
+ wu0 = -2.057536e-11
+ wua = -2.3131395e-16
+ wuc = -1.2695932e-17
+ wwl = 0.0
+ wwn = 1.0
+ xti = 3
+ tcjsw = 0.0004130718
+ tcjswg = 0.0004130718
+ version = 3.24
+ cjsw = 2.35695e-10
+ pvoff = 0.0
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 4.7451600189666944e-17
+ tnom = 25.0
+ )

.model pch_ff_14 pmos (
+ level = 49
+ tpbswg = 0.001572025
+ noimod = 2
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0004772729
+ cit = -0.0001
+ wub1 = -3.0198158e-27
+ wuc1 = -1.0513175e-17
+ pdiblcb = 0.01
+ lpscbe1 = 195.04262
+ dlc = 2e-9
+ hdif = 2e-7
+ k3b = 0.0
+ lub1 = -2.0820251e-25
+ dwb = 0.0
+ dwg = 0.0
+ luc1 = 9.921307e-17
+ wute = 1.1298283e-8
+ mjsw = 0.3683619
+ binunit = 2
+ lketa = -4.562476e-8
+ lute = 2.2927659e-7
+ xpart = 1
+ la0 = 5.081137e-7
+ cdsc = 0.0
+ jsw = 1.2e-12
+ kt1 = -0.2237138
+ lk1 = -4.88067e-8
+ kt2 = -0.026908273
+ lk2 = 2.2115907999999998e-8
+ llc = -0.039
+ lln = -1
+ cgdo = 3.444e-10
+ lu0 = -2.2091919e-10
+ pbswg = 0.895226
+ lua = -3.24011e-17
+ lub = -3.941427e-28
+ luc = -6.882293e-17
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ cgso = 3.444e-10
+ pa0 = -1.854315e-13
+ lvoff = -8.068828999999997e-10
+ nlx = 0.0
+ capmod = 3
+ pk1 = 3.786126e-14
+ pk2 = -1.6169635e-14
+ beta0 = 22.67827
+ pu0 = -6.225135e-16
+ leta0 = 4.745160018966694e-10
+ prt = 0
+ pua = -1.3939852e-23
+ pub = 1.1764949e-34
+ puc = 1.4094153e-23
+ cjsw = 2.35695e-10
+ lvsat = -0.013002842
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ lvth0 = -6.54035e-10
+ version = 3.24
+ rsh = 7.2
+ tcj = 0.0009739001
+ mobmod = 1
+ ua1 = 1.224e-9
+ ub1 = -1.2832692e-18
+ uc1 = 5.668055e-11
+ tpb = 0.001572025
+ tox = 4.02740781e-9
+ delta = 0.01
+ wa0 = 1.0814799e-7
+ tnom = 25.0
+ ute = -0.790886
+ wk1 = -2.4364055e-10
+ wk2 = -3.0947396e-9
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ wln = 1.0
+ wu0 = 4.1988812999999995e-11
+ toxm = 4.08e-9
+ wua = -2.2991296e-16
+ wub = -1.1822094e-29
+ wuc = -1.4112429e-17
+ wwl = 0.0
+ wwn = 1.0
+ pbsw = 0.895226
+ xti = 3
+ pclm = 0.5738635
+ pketa = 1.7549415e-14
+ a0 = 0.8193527
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ at = 10000.0
+ cf = 0
+ cj = 0.00106495
+ ef = 1.064
+ k1 = 0.5470301
+ k2 = 0.027798470000000002
+ k3 = 0.0
+ em = 30000000.0
+ js = 2.5e-7
+ ll = 0.0
+ mj = 0.4476
+ lw = 0.0
+ u0 = 0.0098338462
+ pb = 0.895226
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ua = 1.2617201e-9
+ ub = 5.00396e-20
+ uc = -1.5373321e-10
+ wl = 0.0
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -2.5259219000000002e-8
+ ww = 0.0
+ tcjswg = 0.0004130718
+ xw = 8.69946e-9
+ tcjsw = 0.0004130718
+ pkt1 = 2.5501714e-15
+ pkt2 = -4.817884e-16
+ keta = 0.04769481
+ pvoff = 2.6840621e-15
+ dsub = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 4.7451600189666944e-17
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ pnfactor = 0
+ wketa = -8.167253e-9
+ pvth0 = -2.454092e-15
+ wnfactor = 0.0
+ voff = -0.1259132
+ drout = 0.0
+ ldif = 9e-8
+ tpbsw = 0.001572025
+ kt1l = 0.0
+ prwb = 0.0
+ pub1 = 5.158311e-32
+ prwg = 0.0
+ puc1 = -2.0035212e-23
+ eta0 = 5e-5
+ cjswg = 4.00995e-10
+ pvag = 0.0
+ etab = -5e-5
+ vsat = 151306.8
+ mjswg = 0.3683619
+ wint = 5e-9
+ pute = -4.378173e-14
+ vth0 = -0.4242777
+ rdsw = 530.0
+ lnfactor = 3.9543e-9
+ wvoff = -1.590053e-9
+ wkt1 = 3.574256e-9
+ wkt2 = 2.0011981e-9
+ lint = 1.4999999e-8
+ wmax = 4.9130054e-7
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ wmin = 2.2e-7
+ lkt1 = -1.0417262e-8
+ lkt2 = -1.6001408e-9
+ weta0 = 0
+ nfactor = 1.0
+ lmax = 1.0005259219000001e-5
+ pscbe1 = 180397700.0
+ pscbe2 = 5e-7
+ wvsat = 0.0
+ lmin = 1.205259219e-6
+ lpclm = 2.6005691e-7
+ wvth0 = 1.089277e-8
+ lpdiblc2 = 5.201136e-9
+ ags = 0.02
+ nqsmod = 0
+ )

.model pch_ff_15 pmos (
+ level = 49
+ ute = -0.5904401
+ wk1 = 4.182789e-8
+ wk2 = -2.2085489e-8
+ beta0 = 22.67827
+ wln = 1.0
+ wu0 = -3.789626e-10
+ pkt1 = -8.599671e-15
+ pkt2 = 1.9347028e-16
+ lpdiblc2 = 3.696429e-9
+ keta = 0.0004484208
+ wua = -1.9008923e-16
+ leta0 = 5.114802818966694e-10
+ wub = 8.369847e-27
+ wuc = 5.370726e-18
+ wwl = 0.0
+ wwn = 1.0
+ letab = -3.696428e-11
+ xti = 3
+ mobmod = 1
+ lvsat = -0.007392816
+ dsub = 0.0
+ lvth0 = -1.1578233000000001e-8
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ delta = 0.01
+ lcit = 2.2622144e-10
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ voff = -0.1186655
+ ldif = 9e-8
+ kt1l = 0.0
+ prwb = 0.0
+ pub1 = -1.2589071e-33
+ prwg = 0.0
+ puc1 = 4.27717e-24
+ eta0 = 1.7857146e-5
+ pvag = 0.0
+ etab = -1.7857146e-5
+ vsat = 146428.52
+ wint = 5e-9
+ pute = -8.783067e-15
+ vth0 = -0.4147784
+ rdsw = 530.0
+ pketa = -5.090041e-15
+ wkt1 = 1.3269771e-8
+ wkt2 = 1.4140165e-9
+ lint = 1.4999999e-8
+ wmax = 4.9130054e-7
+ tcjswg = 0.0004130718
+ wmin = 2.2e-7
+ lkt1 = 1.1386779e-8
+ lkt2 = -8.841858e-10
+ lmax = 1.205259219e-6
+ lmin = 5.052592189999999e-7
+ tcjsw = 0.0004130718
+ nfactor = 1.0
+ pvoff = 3.95383e-15
+ wub1 = 4.292976e-26
+ cdscb = 0.0
+ wuc1 = -3.165437e-17
+ cdscd = 0.0
+ peta0 = 4.7451600189666944e-17
+ hdif = 2e-7
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0017857139
+ pdiblcb = 0.01
+ lub1 = -9.299159e-27
+ wketa = 1.1519229e-8
+ luc1 = 4.434689e-18
+ pvth0 = 1.9485986e-15
+ wute = -1.9135335e-8
+ mjsw = 0.3683619
+ drout = 0.0
+ tpbsw = 0.001572025
+ lute = -1.2362289e-9
+ cjswg = 4.00995e-10
+ binunit = 2
+ mjswg = 0.3683619
+ ags = 0.02
+ cdsc = 0.0
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ wvoff = -2.6941984e-9
+ cit = -0.00029671428
+ cgdo = 3.444e-10
+ pscbe1 = 349999900.0
+ pscbe2 = 5e-7
+ dlc = 2e-9
+ cgso = 3.444e-10
+ k3b = 0.0
+ weta0 = 0
+ dwb = 0.0
+ dwg = 0.0
+ wvsat = 0.0
+ lpclm = 1.4785714e-7
+ wvth0 = 7.064344e-9
+ nqsmod = 0
+ a0 = 1.1508681
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ tpbswg = 0.001572025
+ cjsw = 2.35695e-10
+ noimod = 2
+ at = 10000.0
+ cf = 0
+ cj = 0.00106495
+ ef = 1.064
+ k1 = 0.510219
+ k2 = 0.04857026
+ k3 = 0.0
+ em = 30000000.0
+ js = 2.5e-7
+ ll = 0.0
+ noia = 9.5e+18
+ mj = 0.4476
+ noib = 100000.0
+ noic = 1.4e-12
+ lw = 0.0
+ u0 = 0.0092586472
+ pb = 0.895226
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ua = 1.0922192e-9
+ ub = 2.0536515e-20
+ uc = -2.183638e-10
+ la0 = 1.2687106e-7
+ wl = 0.0
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -2.5259219000000002e-8
+ ww = 0.0
+ xw = 8.69946e-9
+ jsw = 1.2e-12
+ version = 3.24
+ kt1 = -0.2426738
+ lk1 = -6.473878e-9
+ kt2 = -0.027530843
+ lk2 = -1.7716528e-9
+ llc = -0.039
+ lln = -1
+ pnfactor = 0
+ lu0 = 4.405597e-10
+ tnom = 25.0
+ lua = 1.6252487e-16
+ lub = 3.353441e-26
+ luc = 5.502275e-18
+ nch = 3.9e+17
+ wnfactor = 0.0
+ lwl = 0.0
+ lwn = 1.0
+ pa0 = 5.971399e-14
+ nlx = 0.0
+ toxm = 4.08e-9
+ lketa = 8.708591e-9
+ pk1 = -1.0521005e-14
+ pk2 = 5.669729e-15
+ pbsw = 0.895226
+ pclm = 0.6714286
+ pu0 = -1.384194e-16
+ xpart = 1
+ prt = 0
+ pua = -5.973716e-23
+ pub = -9.521269e-33
+ puc = -8.311478e-24
+ rsh = 7.2
+ lnfactor = 3.9543e-9
+ tcj = 0.0009739001
+ ua1 = 1.224e-9
+ ub1 = -1.4562286e-18
+ uc1 = 1.3909653e-10
+ pbswg = 0.895226
+ capmod = 3
+ tpb = 0.001572025
+ tox = 4.02740781e-9
+ wa0 = -1.0502199e-7
+ lvoff = -9.141699e-9
+ )

.model pch_ff_16 pmos (
+ level = 49
+ cdsc = 0.0
+ binunit = 2
+ pketa = 7.45672e-16
+ lnfactor = 3.9543e-9
+ tcjswg = 0.0004130718
+ cgdo = 3.444e-10
+ wpclm = 4.634222e-9
+ cgso = 3.444e-10
+ tcjsw = 0.0004130718
+ lpdiblc2 = 1.8281252e-9
+ cjsw = 2.35695e-10
+ pvoff = 1.4541431e-15
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ wcdscd = -1.4183201e-11
+ ags = 0.03625
+ cdscb = 0.0
+ cdscd = -6.449223e-5
+ peta0 = 4.7451600189666944e-17
+ cit = 8.534377e-5
+ tnom = 25.0
+ wketa = -1.4490222e-9
+ pvth0 = 9.0214192e-16
+ version = 3.24
+ dlc = 2e-9
+ drout = 0.0
+ pcdscd = 6.382441e-18
+ tpbsw = 0.001572025
+ k3b = 0.0
+ toxm = 4.08e-9
+ dwb = 0.0
+ dwg = 0.0
+ pbsw = 0.895226
+ pclm = 0.9648299
+ cjswg = 4.00995e-10
+ mjswg = 0.3683619
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ wvoff = 2.8606606e-9
+ pscbe1 = 350000000.0
+ pscbe2 = 5e-7
+ la0 = 7.233052e-9
+ jsw = 1.2e-12
+ kt1 = -0.2130934
+ lk1 = 1.3789155e-8
+ kt2 = -0.03589084
+ lk2 = -4.293236e-9
+ llc = -0.039
+ weta0 = 0
+ lln = -1
+ lu0 = -2.775402e-10
+ nqsmod = 0
+ lua = -2.6402067e-16
+ lub = 2.6345733e-25
+ luc = 3.340897e-17
+ nch = 3.9e+17
+ wvsat = 0.0
+ tpbswg = 0.001572025
+ lwl = 0.0
+ lwn = 1.0
+ noimod = 2
+ lpclm = 1.5826547e-8
+ pa0 = -6.072043e-15
+ wvth0 = 9.389803e-9
+ nlx = 0.0
+ pkt1 = -9.758805e-16
+ pkt2 = -1.0643102e-15
+ keta = 0.03159368
+ pk1 = 4.122718e-15
+ pk2 = -2.3103772e-15
+ dsub = 0.0
+ pu0 = 1.3574996e-16
+ prt = 0
+ pua = 6.304761e-23
+ pub = -7.522618e-32
+ puc = -8.758834e-24
+ lags = -7.312499e-9
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ rsh = 7.2
+ tcj = 0.0009739001
+ ua1 = 1.224e-9
+ ub1 = -1.4433942e-18
+ uc1 = 2.0396977e-10
+ tpb = 0.001572025
+ tox = 4.02740781e-9
+ lcit = 5.429531e-11
+ voff = -0.1287204
+ wa0 = 4.116919e-8
+ lcdscd = 2.9021494e-11
+ ldif = 9e-8
+ ute = -0.5893072
+ wk1 = 9.286284e-9
+ kt1l = 0.0
+ wk2 = -4.351921e-9
+ prwb = 0.0
+ pub1 = 1.9106841e-32
+ prwg = 0.0
+ lketa = -5.306775e-9
+ puc1 = 6.153712e-24
+ wln = 1.0
+ wu0 = -9.882279e-10
+ eta0 = -0.0004687502
+ wua = -4.629443e-16
+ pvag = 0.0
+ wub = 1.5438073e-25
+ wuc = 6.364847e-18
+ etab = 0.0006718753
+ xpart = 1
+ wwl = 0.0
+ wwn = 1.0
+ vsat = 130812.55
+ xti = 3
+ wint = 5e-9
+ pute = 5.968411e-15
+ vth0 = -0.4276605
+ capmod = 3
+ rdsw = 530.0
+ wkt1 = -3.671987e-9
+ wkt2 = 4.209085e-9
+ pbswg = 0.895226
+ lint = 1.4999999e-8
+ wmax = 4.9130054e-7
+ wmin = 2.2e-7
+ lvoff = -4.616999000000001e-9
+ lkt1 = -1.9244071e-9
+ lkt2 = 2.877812e-9
+ lmax = 5.052592189999999e-7
+ beta0 = 22.67827
+ lmin = 1.8e-7
+ mobmod = 1
+ leta0 = 7.304535818966694e-10
+ letab = -3.473438e-10
+ lvsat = -0.0003656336
+ nfactor = 1.0
+ lvth0 = -5.781281000000001e-9
+ ppclm = -2.0853998e-15
+ wub1 = -2.3274574e-27
+ wuc1 = -3.582447e-17
+ delta = 0.01
+ hdif = 2e-7
+ a0 = 1.4167303
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ pnfactor = 0
+ lub1 = -1.5074642e-26
+ luc1 = -2.4758267e-17
+ at = 10000.0
+ cf = 0
+ cj = 0.00106495
+ ef = 1.064
+ k1 = 0.46519
+ dvt0w = 0.0
+ k2 = 0.05417378
+ k3 = 0.0
+ em = 30000000.0
+ wnfactor = 0.0
+ wute = -5.191639e-8
+ dvt1w = 0.0
+ dvt2w = 0.0
+ mjsw = 0.3683619
+ js = 2.5e-7
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.005937499
+ ll = 0.0
+ mj = 0.4476
+ lw = 0.0
+ u0 = 0.0108544242
+ pb = 0.895226
+ w0 = 0.0
+ rd = 0
+ pdiblcb = 0.01
+ rs = 0
+ ua = 2.0400983e-9
+ ub = -4.904033e-19
+ uc = -2.8037866e-10
+ wl = 0.0
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -2.5259219000000002e-8
+ ww = 0.0
+ lute = -1.7460413e-9
+ xw = 8.69946e-9
+ )

.model pch_tt_1 pmos (
+ level = 49
+ lvth0 = 0.0
+ cdsc = 0.0
+ binunit = 2
+ pnfactor = 0
+ cgdo = 3.28e-10
+ delta = 0.01
+ wnfactor = 0.0
+ cgso = 3.28e-10
+ dvt0w = 0.0
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ dvt1w = 0.0
+ dvt2w = 0.0
+ pscbe1 = 199999970.0
+ pscbe2 = 5e-7
+ cjsw = 2.481e-10
+ ags = 0.02
+ lnfactor = 0.0
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ nqsmod = 0
+ tpbswg = 0.001572025
+ noimod = 2
+ cit = -0.0001
+ dlc = 2e-9
+ tnom = 25.0
+ version = 3.24
+ k3b = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ toxm = 4.08e-9
+ tcjsw = 0.0004130718
+ pbsw = 0.895226
+ pclm = 0.6000001
+ pvoff = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ jsw = 1.2e-12
+ peta0 = 3.0000000000000003e-21
+ kt1 = -0.2311294
+ lk2 = 0.0
+ kt2 = -0.02433992
+ llc = -0.039
+ lln = -1
+ lu0 = 0.0
+ nch = 3.9e+17
+ pvth0 = 0.0
+ lwl = 0.0
+ lwn = 1.0
+ drout = 0.0
+ nlx = 0.0
+ tpbsw = 0.001572025
+ capmod = 3
+ keta = 0.026632193
+ pu0 = 0.0
+ cjswg = 4.221e-10
+ prt = 0
+ dsub = 0.0
+ mjswg = 0.3683619
+ rsh = 7.2
+ tcj = 0.0009739001
+ ua1 = 1.224e-9
+ ub1 = -1.3928839e-18
+ uc1 = -4.59467e-12
+ wvoff = 0.0
+ mobmod = 1
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ tpb = 0.001572025
+ tox = 4.08e-9
+ ute = -0.8288856
+ voff = -0.1275921
+ weta0 = 0
+ ldif = 9e-8
+ wvsat = 0.0
+ wln = 1.0
+ kt1l = 0.0
+ prwb = 0.0
+ wu0 = 0.0
+ prwg = 0.0
+ wvth0 = 0.0
+ wwl = 0.0
+ wwn = 1.0
+ eta0 = 5e-5
+ xti = 3
+ pvag = 0.0
+ etab = -5e-5
+ vsat = 149999.98
+ wint = 5e-9
+ vth0 = -0.4384811
+ rdsw = 530.0
+ lint = 1.4999999e-8
+ wmax = 0.000900001
+ wmin = 1e-5
+ a0 = 1.0461572
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ lmax = 2.0001e-5
+ at = 10000.0
+ cf = 0
+ cj = 0.001121
+ lmin = 1e-5
+ ef = 1.064
+ k1 = 0.5375325
+ k2 = 0.03503256
+ k3 = 0.0
+ em = 30000000.0
+ tcjswg = 0.0004130718
+ js = 2.5e-7
+ ll = 0.0
+ mj = 0.4476
+ lw = 0.0
+ u0 = 0.010865118
+ pb = 0.895226
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ua = 8.23294e-10
+ ub = 6.854322e-19
+ uc = -8.655411e-11
+ wl = 0.0
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ xpart = 1
+ nfactor = 1.0
+ pbswg = 0.895226
+ hdif = 2e-7
+ lvoff = 0.0
+ mjsw = 0.3683619
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0010000003
+ pdiblcb = 0.01
+ beta0 = 22.67827
+ leta0 = 3e-14
+ )

.model pch_tt_2 pmos (
+ level = 49
+ mj = 0.4476
+ lw = 0.0
+ kt1 = -0.2295883
+ lk1 = 1.8783622e-8
+ kt2 = -0.024031118
+ lk2 = -5.487172e-9
+ u0 = 0.010995165
+ pb = 0.895226
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ua = 8.625313e-10
+ ub = 6.401998e-19
+ uc = -8.855145e-11
+ llc = -0.039
+ lln = -1
+ wl = 0.0
+ lu0 = -1.2939689e-9
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ voff = -0.1274002
+ lua = -3.904111e-16
+ lub = 4.500626e-25
+ luc = 1.9873557e-17
+ ldif = 9e-8
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ kt1l = 0.0
+ tcjsw = 0.0004130718
+ prwb = 0.0
+ prwg = 0.0
+ nlx = 0.0
+ eta0 = 5e-5
+ pvag = 0.0
+ etab = -5e-5
+ pvoff = 0.0
+ vsat = 151306.8
+ pu0 = 0.0
+ wint = 5e-9
+ prt = 0
+ vth0 = -0.4359872
+ rdsw = 530.0
+ pnfactor = 0
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 3.0000000000000003e-21
+ lint = 1.4999999e-8
+ rsh = 7.2
+ tcj = 0.0009739001
+ ua1 = 1.224e-9
+ wnfactor = 0.0
+ wmax = 0.000900001
+ ub1 = -1.3977103e-18
+ uc1 = -6.694918e-12
+ wmin = 1e-5
+ tpb = 0.001572025
+ capmod = 3
+ pvth0 = 0.0
+ tox = 4.08e-9
+ lkt1 = -1.5333228e-8
+ lkt2 = -3.0725886e-9
+ drout = 0.0
+ lmax = 1e-5
+ tpbsw = 0.001572025
+ ute = -0.8385549
+ lmin = 1.2e-6
+ wln = 1.0
+ wu0 = 0.0
+ cjswg = 4.221e-10
+ wwl = 0.0
+ wwn = 1.0
+ mjswg = 0.3683619
+ lnfactor = 0.0
+ xti = 3
+ mobmod = 1
+ nfactor = 1.0
+ wvoff = 0.0
+ hdif = 2e-7
+ lub1 = 4.802326e-26
+ luc1 = 2.0897466e-17
+ weta0 = 0
+ mjsw = 0.3683619
+ lpdiblc2 = 5.201137e-9
+ wvsat = 0.0
+ lute = 9.620972e-8
+ lpclm = 2.6005682e-7
+ wvth0 = 0.0
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0004772727
+ pdiblcb = 0.01
+ lpscbe1 = 195.04263
+ cdsc = 0.0
+ cgdo = 3.28e-10
+ binunit = 2
+ cgso = 3.28e-10
+ tcjswg = 0.0004130718
+ lketa = -2.0462676e-9
+ cjsw = 2.481e-10
+ xpart = 1
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ pbswg = 0.895226
+ tnom = 25.0
+ lvoff = -1.9091309e-9
+ toxm = 4.08e-9
+ beta0 = 22.67827
+ version = 3.24
+ pbsw = 0.895226
+ pclm = 0.5738637
+ leta0 = 3e-14
+ lvsat = -0.013002843
+ lvth0 = -2.4814053e-8
+ ags = 0.02
+ delta = 0.01
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ cit = -0.0001
+ dlc = 2e-9
+ dvt0w = 0.0
+ dvt1w = 0.0
+ pscbe1 = 180397680.0
+ pscbe2 = 5e-7
+ dvt2w = 0.0
+ k3b = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ keta = 0.026837848
+ nqsmod = 0
+ tpbswg = 0.001572025
+ dsub = 0.0
+ noimod = 2
+ a0 = 1.0385712
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ at = 10000.0
+ cf = 0
+ cj = 0.001121
+ la0 = 7.548124e-8
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ ef = 1.064
+ k1 = 0.5356447
+ k2 = 0.03558403
+ k3 = 0.0
+ em = 30000000.0
+ js = 2.5e-7
+ jsw = 1.2e-12
+ ll = 0.0
+ )

.model pch_tt_3 pmos (
+ level = 49
+ cjswg = 4.221e-10
+ mjswg = 0.3683619
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ wvoff = 0.0
+ tnom = 25.0
+ weta0 = 0
+ wvsat = 0.0
+ toxm = 4.08e-9
+ a0 = 1.0045335
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ lpclm = 1.4785704e-7
+ wvth0 = 0.0
+ pbsw = 0.895226
+ pclm = 0.6714287
+ at = 10000.0
+ cf = 0
+ cj = 0.001121
+ ef = 1.064
+ k1 = 0.5405614
+ k2 = 0.03490157
+ k3 = 0.0
+ em = 30000000.0
+ js = 2.5e-7
+ version = 3.24
+ ll = 0.0
+ mj = 0.4476
+ lw = 0.0
+ u0 = 0.010224584
+ pb = 0.895226
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ua = 5.26694e-10
+ ub = 1.1734415e-18
+ uc = -4.332115e-11
+ wl = 0.0
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ pnfactor = 0
+ wnfactor = 0.0
+ tcjswg = 0.0004130718
+ lketa = -8.158225e-9
+ keta = 0.03215259
+ xpart = 1
+ dsub = 0.0
+ lnfactor = 0.0
+ ags = 0.02
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ pbswg = 0.895226
+ lvoff = -9.487825e-10
+ lcit = 2.2402701e-10
+ cit = -0.00029480609
+ voff = -0.1282353
+ lpdiblc2 = 3.696428e-9
+ ldif = 9e-8
+ dlc = 2e-9
+ beta0 = 22.67827
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ k3b = 0.0
+ dwb = 0.0
+ leta0 = 3.699428e-11
+ dwg = 0.0
+ eta0 = 1.7857143e-5
+ letab = -3.696428e-11
+ pvag = 0.0
+ etab = -1.7857143e-5
+ lvsat = -0.007392833
+ vsat = 146428.53
+ wint = 5e-9
+ lvth0 = -6.689442e-9
+ vth0 = -0.4517478
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ rdsw = 530.0
+ delta = 0.01
+ lint = 1.4999999e-8
+ wmax = 0.000900001
+ pscbe1 = 349999900.0
+ pscbe2 = 5e-7
+ la0 = 1.146246e-7
+ wmin = 1e-5
+ jsw = 1.2e-12
+ lkt1 = 1.5747348e-9
+ lkt2 = 9.740028e-10
+ kt1 = -0.2442909
+ lk1 = 1.3129389e-8
+ kt2 = -0.027549893
+ lk2 = -4.702335e-9
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ lmax = 1.2e-6
+ llc = -0.039
+ lln = -1
+ lu0 = -4.078006e-10
+ lmin = 5e-7
+ lua = -4.198125e-18
+ lub = -1.631654e-25
+ luc = -3.214129e-17
+ nch = 3.9e+17
+ nqsmod = 0
+ lwl = 0.0
+ lwn = 1.0
+ tpbswg = 0.001572025
+ noimod = 2
+ nlx = 0.0
+ pu0 = 0.0
+ prt = 0
+ hdif = 2e-7
+ rsh = 7.2
+ tcj = 0.0009739001
+ nfactor = 1.0
+ ua1 = 1.224e-9
+ lub1 = 3.0810812e-26
+ ub1 = -1.3827429e-18
+ luc1 = 2.9752128e-17
+ uc1 = -1.4394627e-11
+ mjsw = 0.3683619
+ tpb = 0.001572025
+ tox = 4.08e-9
+ tcjsw = 0.0004130718
+ lute = 3.654092e-8
+ ute = -0.786669
+ wln = 1.0
+ pvoff = 0.0
+ wu0 = 0.0
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0017857148
+ wwl = 0.0
+ wwn = 1.0
+ pdiblcb = 0.01
+ cdsc = 0.0
+ xti = 3
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 3.0000000000000003e-21
+ capmod = 3
+ cgdo = 3.28e-10
+ pvth0 = 0.0
+ cgso = 3.28e-10
+ drout = 0.0
+ binunit = 2
+ tpbsw = 0.001572025
+ cjsw = 2.481e-10
+ mobmod = 1
+ )

.model pch_tt_4 pmos (
+ level = 49
+ wmin = 1e-5
+ lkt1 = -2.665e-9
+ lkt2 = -2.325577e-10
+ lmax = 5e-7
+ cit = -4.054396e-5
+ lmin = 1.8e-7
+ lketa = -8.307595e-10
+ dlc = 2e-9
+ k3b = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ xpart = 1
+ pbswg = 0.895226
+ hdif = 2e-7
+ lub1 = 2.883988e-26
+ luc1 = -6.846759e-18
+ lvoff = -3.571592e-11
+ la0 = 1.6196543e-8
+ mjsw = 0.3683619
+ jsw = 1.2e-12
+ kt1 = -0.2348693
+ lk1 = 1.6807924e-8
+ kt2 = -0.024868647
+ lk2 = -5.876215e-9
+ beta0 = 22.67827
+ nfactor = 1.0
+ llc = -0.039
+ lln = -1
+ lu0 = -9.894781e-11
+ lute = 1.6013461e-9
+ leta0 = 2.5596752e-10
+ lua = -1.5999061e-16
+ lub = 1.2197973e-25
+ luc = 1.8500639e-17
+ nch = 3.9e+17
+ letab = -5.298917e-10
+ lwl = 0.0
+ lwn = 1.0
+ lvsat = -0.0003656265
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ nlx = 0.0
+ lvth0 = -8.240552e-9
+ cdsc = 0.0
+ pscbe1 = 350000000.0
+ pscbe2 = 5e-7
+ pnfactor = 0
+ pu0 = 0.0
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.00796875
+ delta = 0.01
+ a0 = 1.2232625
+ a1 = 0.0
+ a2 = 0.4
+ prt = 0
+ b0 = 0.0
+ b1 = 0.0
+ cgdo = 3.28e-10
+ wnfactor = 0.0
+ pdiblcb = 0.01
+ at = 10000.0
+ cf = 0
+ cj = 0.001121
+ ef = 1.064
+ k1 = 0.5323869
+ k2 = 0.03751019
+ k3 = 0.0
+ em = 30000000.0
+ cgso = 3.28e-10
+ js = 2.5e-7
+ dvt0w = 0.0
+ dvt1w = 0.0
+ ll = 0.0
+ rsh = 7.2
+ mj = 0.4476
+ dvt2w = 0.0
+ lw = 0.0
+ u0 = 0.009538244
+ tcj = 0.0009739001
+ nqsmod = 0
+ pb = 0.895226
+ ua1 = 1.224e-9
+ w0 = 0.0
+ ub1 = -1.3783631e-18
+ rd = 0
+ uc1 = 6.693623e-11
+ tpbswg = 0.001572025
+ rs = 0
+ ua = 8.728995e-10
+ ub = 5.397856e-19
+ uc = -1.5585878e-10
+ noimod = 2
+ wl = 0.0
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ tpb = 0.001572025
+ tox = 4.08e-9
+ binunit = 2
+ cjsw = 2.481e-10
+ ute = -0.7090256
+ lnfactor = 0.0
+ wln = 1.0
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ wu0 = 0.0
+ wwl = 0.0
+ wwn = 1.0
+ xti = 3
+ tnom = 25.0
+ lcdscd = 3.65625e-11
+ lpdiblc2 = 9.140626e-10
+ toxm = 4.08e-9
+ tcjsw = 0.0004130718
+ pbsw = 0.895226
+ pclm = 0.9102259
+ pvoff = 0.0
+ capmod = 3
+ version = 3.24
+ cdscb = 0.0
+ cdscd = -8.125e-5
+ peta0 = 3.0000000000000003e-21
+ pvth0 = 0.0
+ drout = 0.0
+ tpbsw = 0.001572025
+ mobmod = 1
+ keta = 0.015869336
+ cjswg = 4.221e-10
+ mjswg = 0.3683619
+ dsub = 0.0
+ wvoff = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ weta0 = 0
+ lcit = 1.0960905e-10
+ voff = -0.1302643
+ ldif = 9e-8
+ wvsat = 0.0
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ lpclm = 4.03983e-8
+ wvth0 = 0.0
+ eta0 = -0.0004687502
+ pvag = 0.0
+ etab = 0.0010775371
+ vsat = 130812.52
+ wint = 5e-9
+ vth0 = -0.4483009
+ rdsw = 530.0
+ tcjswg = 0.0004130718
+ lint = 1.4999999e-8
+ wmax = 0.000900001
+ ags = 0.02
+ )

.model pch_tt_5 pmos (
+ level = 49
+ wa0 = -4.787191e-8
+ pscbe1 = 199999970.0
+ pscbe2 = 5e-7
+ ute = -0.8394966
+ lvth0 = 0.0
+ wk1 = 1.2456701e-8
+ wk2 = -5.940143e-9
+ wln = 1.0
+ wu0 = -1.2494747e-9
+ delta = 0.01
+ wua = 1.7543858e-16
+ wub = -6.530953e-25
+ wuc = -7.950096e-17
+ wwl = 0.0
+ wwn = 1.0
+ nqsmod = 0
+ xti = 3
+ version = 3.24
+ tpbswg = 0.001572025
+ noimod = 2
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ keta = 0.02600144
+ dsub = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ voff = -0.1274889
+ ldif = 9e-8
+ tcjsw = 0.0004130718
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ eta0 = 5e-5
+ pvoff = 0.0
+ capmod = 3
+ pvag = 0.0
+ etab = -5e-5
+ vsat = 149999.98
+ wint = 5e-9
+ vth0 = -0.4397694
+ cdscb = 0.0
+ rdsw = 530.0
+ cdscd = 0.0
+ pnfactor = 0
+ peta0 = 3.0000000000000003e-21
+ wkt1 = 8.228274e-9
+ wkt2 = 1.4868883e-9
+ lint = 1.4999999e-8
+ wnfactor = 0.0
+ wmax = 1e-5
+ wketa = 6.301227e-9
+ wmin = 1.2e-6
+ pvth0 = 0.0
+ mobmod = 1
+ drout = 0.0
+ tpbsw = 0.001572025
+ lmax = 2.0001e-5
+ lmin = 1e-5
+ cjswg = 4.221e-10
+ a0 = 1.0509492
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ at = 10000.0
+ mjswg = 0.3683619
+ cf = 0
+ cj = 0.001121
+ lnfactor = 0.0
+ ef = 1.064
+ k1 = 0.5362856
+ k2 = 0.03562717
+ k3 = 0.0
+ em = 30000000.0
+ js = 2.5e-7
+ ll = 0.0
+ mj = 0.4476
+ lw = 0.0
+ u0 = 0.010990191
+ pb = 0.895226
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ wvoff = -1.0305298e-9
+ ua = 8.057326e-10
+ ub = 7.508071e-19
+ uc = -7.859605e-11
+ wub1 = 6.909715e-26
+ wuc1 = 3.0354498e-17
+ wl = 0.0
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ hdif = 2e-7
+ weta0 = 0
+ ags = 0.02
+ wute = 1.0600407e-7
+ mjsw = 0.3683619
+ wvsat = 0.0
+ wvth0 = 1.2870458e-8
+ cit = -0.0001
+ dlc = 2e-9
+ nfactor = 1.0
+ k3b = 0.0
+ tcjswg = 0.0004130718
+ dwb = 0.0
+ dwg = 0.0
+ cdsc = 0.0
+ cgdo = 3.28e-10
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0010000004
+ cgso = 3.28e-10
+ pdiblcb = 0.01
+ jsw = 1.2e-12
+ kt1 = -0.231953
+ kt2 = -0.024488758
+ lk2 = 0.0
+ llc = -0.039
+ lln = -1
+ cjsw = 2.481e-10
+ lu0 = 0.0
+ xpart = 1
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ binunit = 2
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ nlx = 0.0
+ pbswg = 0.895226
+ pu0 = 0.0
+ prt = 0
+ tnom = 25.0
+ lvoff = 0.0
+ rsh = 7.2
+ beta0 = 22.67827
+ toxm = 4.08e-9
+ tcj = 0.0009739001
+ ua1 = 1.224e-9
+ ub1 = -1.3998005e-18
+ uc1 = -7.633158e-12
+ leta0 = 3e-14
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ pbsw = 0.895226
+ pclm = 0.6000001
+ tpb = 0.001572025
+ tox = 4.08e-9
+ )

.model pch_tt_6 pmos (
+ level = 49
+ lub1 = 5.442727e-26
+ luc1 = 1.8276951e-17
+ wute = 1.0644106e-7
+ mjsw = 0.3683619
+ tcjsw = 0.0004130718
+ capmod = 3
+ lute = 9.664497e-8
+ pvoff = -4.403278e-15
+ nfactor = 1.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 3.0000000000000003e-21
+ mobmod = 1
+ cgdo = 3.28e-10
+ wketa = 7.084359e-9
+ pvth0 = -5.336472e-15
+ cgso = 3.28e-10
+ drout = 0.0
+ tpbsw = 0.001572025
+ ags = 0.02
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0004772728
+ pdiblcb = 0.01
+ lpscbe1 = 195.04262
+ cjswg = 4.221e-10
+ cit = -0.0001
+ cjsw = 2.481e-10
+ mjswg = 0.3683619
+ dlc = 2e-9
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ k3b = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ wvoff = -5.879894e-10
+ binunit = 2
+ tnom = 25.0
+ weta0 = 0
+ wvsat = 0.0
+ toxm = 4.08e-9
+ lpclm = 2.6005682e-7
+ wvth0 = 1.3406786e-8
+ la0 = 6.878132e-8
+ pbsw = 0.895226
+ tcjswg = 0.0004130718
+ pclm = 0.5738637
+ jsw = 1.2e-12
+ kt1 = -0.2303147
+ lk1 = 1.8184398e-8
+ kt2 = -0.024155809
+ lk2 = -5.280635e-9
+ llc = -0.039
+ lln = -1
+ lu0 = -1.3055237e-9
+ lua = -3.935608e-16
+ lub = 4.219459e-25
+ luc = 1.8883157e-17
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ pnfactor = 0
+ pa0 = 6.693222e-14
+ nlx = 0.0
+ wnfactor = 0.0
+ pk1 = 5.986243e-15
+ pk2 = -2.063307e-15
+ pu0 = 1.1543239e-16
+ prt = 0
+ pua = 3.1465633e-23
+ pub = 2.8088595e-31
+ puc = 9.8941e-24
+ version = 3.24
+ lketa = -1.2662711e-9
+ rsh = 7.2
+ pkt1 = 9.666697e-15
+ tcj = 0.0009739001
+ pkt2 = 2.4000725e-15
+ ua1 = 1.224e-9
+ keta = 0.026128704
+ ub1 = -1.4052706e-18
+ uc1 = -9.470036e-12
+ xpart = 1
+ tpb = 0.001572025
+ lnfactor = 0.0
+ tox = 4.08e-9
+ dsub = 0.0
+ wa0 = -5.459876e-8
+ ute = -0.8492097
+ wk1 = 1.185507e-8
+ wk2 = -5.732776e-9
+ pbswg = 0.895226
+ wln = 1.0
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ wu0 = -1.261076e-9
+ wua = 1.7227619e-16
+ wub = -6.81325e-25
+ wuc = -8.049533e-17
+ wwl = 0.0
+ wwn = 1.0
+ a0 = 1.0440365
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ lvoff = -1.4683624e-9
+ xti = 3
+ at = 10000.0
+ cf = 0
+ lpdiblc2 = 5.201137e-9
+ cj = 0.001121
+ voff = -0.1273414
+ ef = 1.064
+ k1 = 0.534458
+ k2 = 0.03615789
+ k3 = 0.0
+ em = 30000000.0
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ ldif = 9e-8
+ beta0 = 22.67827
+ js = 2.5e-7
+ ll = 0.0
+ mj = 0.4476
+ lw = 0.0
+ u0 = 0.0111214
+ pb = 0.895226
+ kt1l = 0.0
+ w0 = 0.0
+ prwb = 0.0
+ rd = 0
+ pub1 = -6.397619e-32
+ prwg = 0.0
+ leta0 = 3e-14
+ puc1 = 2.6178952e-23
+ rs = 0
+ ua = 8.452865e-10
+ ub = 7.084005e-19
+ uc = -8.049386e-11
+ pscbe1 = 180397700.0
+ pscbe2 = 5e-7
+ wl = 0.0
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ eta0 = 5e-5
+ lvsat = -0.013002842
+ pvag = 0.0
+ etab = -5e-5
+ vsat = 151306.8
+ lvth0 = -2.4279869e-8
+ wint = 5e-9
+ pute = -4.348101e-15
+ vth0 = -0.4373293
+ nqsmod = 0
+ rdsw = 530.0
+ tpbswg = 0.001572025
+ delta = 0.01
+ wkt1 = 7.256747e-9
+ wkt2 = 1.245675e-9
+ noimod = 2
+ lint = 1.4999999e-8
+ wmax = 1e-5
+ wmin = 1.2e-6
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ lkt1 = -1.6300865e-8
+ lkt2 = -3.312836e-9
+ lmax = 1e-5
+ lmin = 1.2e-6
+ pketa = -7.792167e-15
+ wub1 = 7.552692e-26
+ wuc1 = 2.7723443e-17
+ hdif = 2e-7
+ )

.model pch_tt_7 pmos (
+ level = 49
+ mjswg = 0.3683619
+ jsw = 1.2e-12
+ kt1 = -0.2459144
+ lk1 = 8.371453e-9
+ kt2 = -0.027846618
+ lk2 = -3.215854e-9
+ dsub = 0.0
+ llc = -0.039
+ lln = -1
+ lu0 = -3.457226e-10
+ wvoff = -7.866491e-9
+ lua = 3.0792715e-17
+ lub = -1.9665828e-25
+ luc = -3.700045e-17
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ wcit = -1.788104e-11
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ pa0 = -1.2519753e-13
+ nlx = 0.0
+ weta0 = 0
+ pk1 = 4.753178e-14
+ pk2 = -1.4849934e-14
+ lcit = 2.2196864e-10
+ voff = -0.1274479
+ pu0 = -6.201592e-16
+ wvsat = 0.0
+ ldif = 9e-8
+ tcjswg = 0.0004130718
+ prt = 0
+ pua = -3.495584e-22
+ pub = 3.345938e-31
+ puc = 4.854297e-23
+ lpclm = 1.4785702e-7
+ wvth0 = 1.013071e-8
+ kt1l = 0.0
+ prwb = 0.0
+ pub1 = -1.382964e-31
+ prwg = 0.0
+ puc1 = -5.043768e-23
+ eta0 = 1.7857139e-5
+ rsh = 7.2
+ tcj = 0.0009739001
+ ua1 = 1.224e-9
+ pvag = 0.0
+ ub1 = -1.3967723e-18
+ etab = -1.7857139e-5
+ uc1 = -2.3838735e-11
+ vsat = 146428.53
+ wint = 5e-9
+ pute = 2.0900147e-14
+ tpb = 0.001572025
+ tox = 4.08e-9
+ vth0 = -0.4527619
+ wa0 = 1.1247056e-7
+ rdsw = 530.0
+ ute = -0.7951261
+ wkt1 = 1.6218328e-8
+ wkt2 = 2.9642964e-9
+ wk1 = -2.4271484e-8
+ wk2 = 5.386031e-9
+ lint = 1.4999999e-8
+ wmax = 1e-5
+ wln = 1.0
+ wu0 = -6.214311e-10
+ wmin = 1.2e-6
+ wua = 5.036014e-16
+ wub = -7.280275e-25
+ wuc = -1.1410304e-16
+ lkt1 = 1.6387112e-9
+ lkt2 = 9.315946e-10
+ wwl = 0.0
+ wwn = 1.0
+ xti = 3
+ lmax = 1.2e-6
+ lketa = -8.380984e-9
+ lmin = 5e-7
+ xpart = 1
+ wub1 = 1.4015321e-25
+ pbswg = 0.895226
+ wuc1 = 9.434661e-17
+ hdif = 2e-7
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ lvoff = -1.3458795e-9
+ lub1 = 4.46543e-26
+ luc1 = 3.480094e-17
+ wute = 8.448607e-8
+ mjsw = 0.3683619
+ pscbe1 = 349999900.0
+ pscbe2 = 5e-7
+ beta0 = 22.67827
+ leta0 = 3.699429e-11
+ lute = 3.444881e-8
+ letab = -3.696429e-11
+ lvsat = -0.007392833
+ lvth0 = -6.532387e-9
+ nqsmod = 0
+ tpbswg = 0.001572025
+ noimod = 2
+ cdsc = 0.0
+ pnfactor = 0
+ delta = 0.01
+ wnfactor = 0.0
+ cgdo = 3.28e-10
+ nfactor = 1.0
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ cgso = 3.28e-10
+ cjsw = 2.481e-10
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0017857144
+ lnfactor = 0.0
+ pdiblcb = 0.01
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ pketa = 2.2253538e-15
+ tnom = 25.0
+ binunit = 2
+ capmod = 3
+ lpdiblc2 = 3.696428e-9
+ tcjsw = 0.0004130718
+ toxm = 4.08e-9
+ ags = 0.02
+ pcit = 2.0563189e-17
+ pbsw = 0.895226
+ pclm = 0.6714287
+ pvoff = 3.966999e-15
+ cit = -0.0002930162
+ a0 = 0.9932752
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ at = 10000.0
+ mobmod = 1
+ cf = 0
+ dlc = 2e-9
+ cj = 0.001121
+ ef = 1.064
+ k1 = 0.542991
+ k2 = 0.03436242
+ k3 = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ em = 30000000.0
+ peta0 = 3.0000000000000003e-21
+ k3b = 0.0
+ js = 2.5e-7
+ ll = 0.0
+ mj = 0.4476
+ lw = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ u0 = 0.010286789
+ pb = 0.895226
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ua = 4.762835e-10
+ ub = 1.2463172e-18
+ uc = -3.189942e-11
+ wl = 0.0
+ wr = 1.0
+ xj = 1.7000001e-7
+ wketa = -1.6265284e-9
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ pvth0 = -1.5689828e-15
+ drout = 0.0
+ tpbsw = 0.001572025
+ pkt1 = -6.391237e-16
+ pkt2 = 4.236579e-16
+ keta = 0.03231541
+ cjswg = 4.221e-10
+ version = 3.24
+ la0 = 1.2715688e-7
+ )

.model pch_tt_8 pmos (
+ level = 49
+ cgso = 3.28e-10
+ nfactor = 1.0
+ a0 = 1.2640158
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ lketa = -5.872592e-10
+ at = 10000.0
+ cf = 0
+ cj = 0.001121
+ ef = 1.064
+ k1 = 0.5203763
+ k2 = 0.04193926
+ k3 = 0.0
+ em = 30000000.0
+ pcdscd = -7.408954e-18
+ js = 2.5e-7
+ ll = 0.0
+ mj = 0.4476
+ lw = 0.0
+ u0 = 0.009795761
+ pb = 0.895226
+ xpart = 1
+ w0 = 0.0
+ rd = 0
+ cjsw = 2.481e-10
+ rs = 0
+ ua = 9.357863e-10
+ ub = 5.091257e-19
+ uc = -1.5731644e-10
+ wl = 0.0
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.007987866
+ pbswg = 0.895226
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ pdiblcb = 0.01
+ pscbe1 = 350000000.0
+ pscbe2 = 5e-7
+ lvoff = 1.6353495e-10
+ tnom = 25.0
+ pags = -6.875222e-16
+ beta0 = 22.67827
+ toxm = 4.08e-9
+ binunit = 2
+ leta0 = 2.5596752e-10
+ letab = -5.545772e-10
+ nqsmod = 0
+ pcit = -7.907631e-17
+ pbsw = 0.895226
+ pclm = 0.9107697
+ tpbswg = 0.001572025
+ lvsat = -0.0003656271
+ noimod = 2
+ lvth0 = -8.128026e-9
+ ppclm = 2.4445072e-15
+ delta = 0.01
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ lcdscd = 3.730414e-11
+ pkt1 = -1.8229216e-15
+ pkt2 = -1.2254391e-15
+ keta = 0.014996022
+ ags = 0.019847063
+ wags = 1.5278273e-9
+ dsub = 0.0
+ version = 3.24
+ cit = -6.09184e-5
+ pketa = -2.4325694e-15
+ dlc = 2e-9
+ lags = 6.882101e-11
+ wcit = 2.0354016e-10
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ k3b = 0.0
+ capmod = 3
+ dwb = 0.0
+ dwg = 0.0
+ wpclm = -5.432238e-9
+ lcit = 1.1752459e-10
+ voff = -0.1308021
+ tcjsw = 0.0004130718
+ ldif = 9e-8
+ kt1l = 0.0
+ prwb = 0.0
+ pub1 = 2.7781507e-32
+ prwg = 0.0
+ puc1 = 8.113434e-24
+ pvoff = -1.9905158e-15
+ eta0 = -0.0004687502
+ mobmod = 1
+ pvag = 0.0
+ etab = 0.0011323938
+ la0 = 5.323636e-9
+ vsat = 130812.52
+ wint = 5e-9
+ pute = 9.798417e-15
+ jsw = 1.2e-12
+ kt1 = -0.2367561
+ lk1 = 1.854804e-8
+ kt2 = -0.025532207
+ lk2 = -6.625426e-9
+ vth0 = -0.449216
+ cdscb = 0.0
+ cdscd = -8.289813e-5
+ pnfactor = 0
+ peta0 = 3.0000000000000003e-21
+ llc = -0.039
+ rdsw = 530.0
+ lln = -1
+ lu0 = -1.2475933e-10
+ petab = 2.4660761e-16
+ wnfactor = 0.0
+ wkt1 = 1.8848993e-8
+ wkt2 = 6.628956e-9
+ lua = -1.759835e-16
+ lub = 1.3507784e-25
+ luc = 1.9437196e-17
+ lint = 1.4999999e-8
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ wmax = 1e-5
+ wketa = 8.724413e-9
+ pvth0 = -1.1241356e-15
+ pa0 = 1.0862038e-13
+ nlx = 0.0
+ wmin = 1.2e-6
+ drout = 0.0
+ lkt1 = -2.4825255e-9
+ lkt2 = -1.0989117e-10
+ tpbsw = 0.001572025
+ pk1 = -1.7383759e-14
+ pk2 = 7.484627e-15
+ lmax = 5e-7
+ pu0 = 2.5785697e-16
+ lmin = 1.8e-7
+ ppdiblc2 = 8.594017e-17
+ prt = 0
+ pua = 1.5976873e-22
+ pub = -1.3085017e-31
+ puc = -9.356197e-24
+ cjswg = 4.221e-10
+ wpdiblc2 = -1.9097854e-10
+ mjswg = 0.3683619
+ lnfactor = 0.0
+ rsh = 7.2
+ tcj = 0.0009739001
+ ua1 = 1.224e-9
+ ub1 = -1.3554493e-18
+ uc1 = 7.051652e-11
+ wvoff = 5.372431e-9
+ tpb = 0.001572025
+ tox = 4.08e-9
+ wub1 = -2.2890885e-25
+ wuc1 = -3.576699e-17
+ wa0 = -4.071248e-7
+ hdif = 2e-7
+ ute = -0.7199521
+ wk1 = 1.1998529e-7
+ wk2 = -4.424634e-8
+ weta0 = 0
+ tcjswg = 0.0004130718
+ lub1 = 2.6058948e-26
+ luc1 = -7.658915e-18
+ wln = 1.0
+ wetab = -5.480169e-10
+ lpdiblc2 = 9.0546e-10
+ wu0 = -2.5725782e-9
+ wute = 1.0915658e-7
+ mjsw = 0.3683619
+ wvsat = 0.0
+ wua = -6.282368e-16
+ wub = 3.0629255e-25
+ wuc = 1.4561782e-17
+ wwl = 0.0
+ wwn = 1.0
+ lpclm = 4.015361e-8
+ wvth0 = 9.142164e-9
+ xti = 3
+ lute = 6.205235e-10
+ cdsc = 0.0
+ wcdscd = 1.6464351e-11
+ cgdo = 3.28e-10
+ )

.model pch_tt_9 pmos (
+ level = 49
+ pvag = 0.0
+ etab = -5e-5
+ lvth0 = 0.0
+ ags = 0.02
+ vsat = 149999.98
+ wint = 5e-9
+ vth0 = -0.4286388
+ delta = 0.01
+ rdsw = 530.0
+ cit = -0.0001
+ wkt1 = 6.74333e-9
+ wkt2 = 1.2948118e-10
+ lint = 1.4999999e-8
+ dlc = 2e-9
+ wmax = 1.2e-6
+ dvt0w = 0.0
+ k3b = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ wmin = 5e-7
+ dwb = 0.0
+ dwg = 0.0
+ lmax = 2.0001e-5
+ lmin = 1e-5
+ capmod = 3
+ a0 = 0.9810578
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ jsw = 1.2e-12
+ kt1 = -0.2307052
+ kt2 = -0.02334808
+ lk2 = 0.0
+ wub1 = 3.495163e-26
+ wuc1 = 1.9335648e-17
+ at = 10000.0
+ cf = 0
+ cj = 0.001121
+ ef = 1.064
+ k1 = 0.5449055
+ k2 = 0.03384938
+ k3 = 0.0
+ em = 30000000.0
+ llc = -0.039
+ lln = -1
+ lu0 = 0.0
+ hdif = 2e-7
+ js = 2.5e-7
+ ll = 0.0
+ mj = 0.4476
+ lw = 0.0
+ u0 = 0.010132165
+ nch = 3.9e+17
+ pb = 0.895226
+ w0 = 0.0
+ rd = 0
+ lwl = 0.0
+ lwn = 1.0
+ rs = 0
+ ua = 1.0698959e-9
+ ub = 3.0837888e-19
+ uc = -1.1659398e-10
+ wl = 0.0
+ wute = -2.7886795e-9
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ mjsw = 0.3683619
+ nlx = 0.0
+ tcjsw = 0.0004130718
+ mobmod = 1
+ pu0 = 0.0
+ pvoff = 0.0
+ prt = 0
+ rsh = 7.2
+ cdscb = 0.0
+ cdscd = 0.0
+ tcj = 0.0009739001
+ peta0 = 3.0000000000000003e-21
+ cdsc = 0.0
+ ua1 = 1.224e-9
+ ub1 = -1.3711068e-18
+ uc1 = 1.6263793e-12
+ tpb = 0.001572025
+ tox = 4.08e-9
+ cgdo = 3.28e-10
+ wketa = -1.0458587e-9
+ wa0 = 3.529885e-8
+ pvth0 = 0.0
+ drout = 0.0
+ ute = -0.7480742
+ wk1 = 2.1990281e-9
+ cgso = 3.28e-10
+ wk2 = -3.824582e-9
+ tpbsw = 0.001572025
+ wln = 1.0
+ wu0 = -2.284236e-10
+ wua = -1.3891575e-16
+ wub = -1.2660565e-25
+ wuc = -3.428342e-17
+ wwl = 0.0
+ wwn = 1.0
+ cjswg = 4.221e-10
+ nfactor = 1.0
+ xti = 3
+ cjsw = 2.481e-10
+ mjswg = 0.3683619
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ wvoff = -4.105241e-10
+ tcjswg = 0.0004130718
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0009999998
+ weta0 = 0
+ tnom = 25.0
+ pdiblcb = 0.01
+ wvsat = 0.0
+ wvth0 = -3.750611e-10
+ toxm = 4.08e-9
+ pbsw = 0.895226
+ pclm = 0.6
+ binunit = 2
+ pnfactor = 0
+ wnfactor = 0.0
+ keta = 0.03217546
+ xpart = 1
+ lnfactor = 0.0
+ alpha0 = 0.0
+ dsub = 0.0
+ alpha1 = 6.8730453846
+ pbswg = 0.895226
+ pscbe1 = 199999970.0
+ pscbe2 = 5e-7
+ dvt0 = 0.0
+ version = 3.24
+ dvt1 = 0.0
+ dvt2 = 0.0
+ lvoff = 0.0
+ voff = -0.12801
+ beta0 = 22.67827
+ nqsmod = 0
+ ldif = 9e-8
+ tpbswg = 0.001572025
+ noimod = 2
+ leta0 = 3e-14
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ eta0 = 5e-5
+ )

.model pch_tt_10 pmos (
+ level = 49
+ dsub = 0.0
+ wk1 = 1.7598129e-9
+ wk2 = -3.600003e-9
+ wln = 1.0
+ wu0 = -1.9812424e-10
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ wua = -1.6455617e-16
+ wub = -7.150721e-26
+ wuc = -2.8652769e-17
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ wwl = 0.0
+ wwn = 1.0
+ xti = 3
+ pscbe1 = 180397680.0
+ pscbe2 = 5e-7
+ voff = -0.1269095
+ ldif = 9e-8
+ nfactor = 1.0
+ kt1l = 0.0
+ prwb = 0.0
+ pub1 = -8.629597e-32
+ prwg = 0.0
+ puc1 = 1.5034668e-23
+ nqsmod = 0
+ tpbswg = 0.001572025
+ lketa = -6.417587e-9
+ eta0 = 5e-5
+ noimod = 2
+ pvag = 0.0
+ etab = -5e-5
+ vsat = 151306.8
+ wint = 5e-9
+ pute = 3.909688e-14
+ xpart = 1
+ vth0 = -0.4245711
+ rdsw = 530.0
+ wkt1 = 6.495125e-9
+ wkt2 = 2.3726165e-10
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0004772722
+ lint = 1.4999999e-8
+ pdiblcb = 0.01
+ lpscbe1 = 195.04263
+ wmax = 1.2e-6
+ pbswg = 0.895226
+ wmin = 5e-7
+ lkt1 = -1.0252924e-8
+ lkt2 = -3.947785e-10
+ lmax = 1e-5
+ lvoff = -1.0948965e-8
+ lmin = 1.2e-6
+ beta0 = 22.67827
+ binunit = 2
+ leta0 = 3e-14
+ lvsat = -0.013002842
+ lvth0 = -4.047293e-8
+ wub1 = 4.362458e-26
+ wuc1 = 1.7824627e-17
+ capmod = 3
+ hdif = 2e-7
+ delta = 0.01
+ lub1 = 7.318341e-26
+ luc1 = 2.7641896e-17
+ pnfactor = 0
+ wute = -6.718015e-9
+ mjsw = 0.3683619
+ wnfactor = 0.0
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ lute = 6.013659e-8
+ mobmod = 1
+ cdsc = 0.0
+ version = 3.24
+ lnfactor = 0.0
+ pketa = -1.6621007e-15
+ cgdo = 3.28e-10
+ ags = 0.02
+ cgso = 3.28e-10
+ cit = -0.0001
+ tcjsw = 0.0004130718
+ dlc = 2e-9
+ lpdiblc2 = 5.201137e-9
+ cjsw = 2.481e-10
+ k3b = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ pvoff = 6.87864e-15
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 3.0000000000000003e-21
+ tcjswg = 0.0004130718
+ tnom = 25.0
+ wketa = -8.788133e-10
+ pvth0 = 1.393327e-14
+ la0 = 1.2176828e-7
+ drout = 0.0
+ toxm = 4.08e-9
+ jsw = 1.2e-12
+ kt1 = -0.2296747
+ lk1 = 1.9542425e-8
+ kt2 = -0.023308404
+ lk2 = -5.136719e-9
+ tpbsw = 0.001572025
+ pbsw = 0.895226
+ llc = -0.039
+ pclm = 0.5738636
+ lln = -1
+ lu0 = -9.551782e-10
+ lua = -5.815077e-16
+ lub = 1.1186816e-24
+ luc = 7.427734e-17
+ nch = 3.9e+17
+ a0 = 0.9688198
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ lwl = 0.0
+ lwn = 1.0
+ cjswg = 4.221e-10
+ at = 10000.0
+ cf = 0
+ cj = 0.001121
+ pa0 = 3.87773e-15
+ nlx = 0.0
+ ef = 1.064
+ k1 = 0.5429414
+ k2 = 0.03436564
+ k3 = 0.0
+ em = 30000000.0
+ mjswg = 0.3683619
+ js = 2.5e-7
+ ll = 0.0
+ mj = 0.4476
+ lw = 0.0
+ pk1 = 4.370194e-15
+ pk2 = -2.2345663e-15
+ u0 = 0.010228163
+ pb = 0.895226
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ua = 1.1283389e-9
+ ub = 1.9594849e-19
+ uc = -1.2405904e-10
+ wvoff = -1.1018445e-9
+ wl = 0.0
+ pu0 = -3.0147877e-16
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ prt = 0
+ pua = 2.5512236e-22
+ pub = -5.482294e-31
+ puc = -5.602498e-23
+ weta0 = 0
+ rsh = 7.2
+ tcj = 0.0009739001
+ ua1 = 1.224e-9
+ ub1 = -1.3784619e-18
+ uc1 = -1.1517035e-12
+ wvsat = 0.0
+ pkt1 = 2.469645e-15
+ pkt2 = -1.0724159e-15
+ keta = 0.03282044
+ tpb = 0.001572025
+ tox = 4.08e-9
+ lpclm = 2.6005682e-7
+ wvth0 = -1.7753915e-9
+ wa0 = 3.490912e-8
+ ute = -0.754118
+ )

.model pch_tt_11 pmos (
+ level = 49
+ cgso = 3.28e-10
+ a0 = 1.1936638
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ lvoff = 5.237211e-9
+ at = 10000.0
+ cf = 0
+ cj = 0.001121
+ ef = 1.064
+ k1 = 0.4715038
+ k2 = 0.05978675
+ k3 = 0.0
+ em = 30000000.0
+ js = 2.5e-7
+ ll = 0.0
+ mj = 0.4476
+ lw = 0.0
+ beta0 = 22.67827
+ u0 = 0.010727104
+ pb = 0.895226
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ua = 1.036115e-9
+ ub = 1.0523674e-18
+ uc = -7.205117e-11
+ cjsw = 2.481e-10
+ leta0 = 3.6994259999999997e-11
+ wl = 0.0
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ letab = -3.696426e-11
+ lvsat = -0.007392855
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ capmod = 3
+ lvth0 = -3.562702e-9
+ delta = 0.01
+ tnom = 25.0
+ ags = 0.02
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ toxm = 4.08e-9
+ mobmod = 1
+ pcit = -1.0851648e-17
+ pbsw = 0.895226
+ pclm = 0.6714286
+ cit = -0.00031597191
+ dlc = 2e-9
+ k3b = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ pketa = 4.024799e-15
+ la0 = -1.3680231e-7
+ pkt1 = -6.051915e-15
+ pkt2 = -1.4802061e-15
+ tcjsw = 0.0004130718
+ keta = 0.03584265
+ jsw = 1.2e-12
+ kt1 = -0.2439705
+ lk1 = 1.0169572e-7
+ kt2 = -0.025852976
+ lk2 = -3.4371e-8
+ llc = -0.039
+ lln = -1
+ lu0 = -1.5289595e-9
+ dsub = 0.0
+ pvoff = -3.866879e-15
+ lua = -4.754501e-16
+ lub = 1.337998e-25
+ luc = 1.4468274e-17
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ pa0 = 1.8891395e-13
+ nlx = 0.0
+ tcjswg = 0.0004130718
+ wcit = 9.436221e-12
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ pk1 = -6.35241e-14
+ pk2 = 2.2224691e-14
+ peta0 = 3.0000000000000003e-21
+ pu0 = 7.878928e-16
+ pnfactor = 0
+ prt = 0
+ lcit = 2.4836766e-10
+ pua = 2.5287059e-22
+ pub = -5.865131e-32
+ puc = -1.2704817e-23
+ wketa = -5.823942e-9
+ voff = -0.1409845
+ pvth0 = -5.102908e-15
+ wnfactor = 0.0
+ ldif = 9e-8
+ drout = 0.0
+ kt1l = 0.0
+ tpbsw = 0.001572025
+ prwb = 0.0
+ pub1 = 4.97241e-32
+ prwg = 0.0
+ rsh = 7.2
+ puc1 = 1.7282469e-23
+ tcj = 0.0009739001
+ ua1 = 1.224e-9
+ ub1 = -1.2162624e-18
+ uc1 = 4.210797e-11
+ eta0 = 1.7857154e-5
+ nfactor = 1.0
+ pvag = 0.0
+ etab = -1.7857154e-5
+ tpb = 0.001572025
+ tox = 4.08e-9
+ cjswg = 4.221e-10
+ vsat = 146428.56
+ wa0 = -1.2599192e-7
+ wint = 5e-9
+ pute = -5.928695e-14
+ mjswg = 0.3683619
+ vth0 = -0.456667
+ ute = -0.7903757
+ wk1 = 6.079834e-8
+ wk2 = -2.4868919e-8
+ rdsw = 530.0
+ wln = 1.0
+ wkt1 = 1.3905176e-8
+ wkt2 = 5.918618e-10
+ lnfactor = 0.0
+ wu0 = -1.1454039e-9
+ lint = 1.4999999e-8
+ wvoff = 8.242083e-9
+ wua = -1.625981e-16
+ wmax = 1.2e-6
+ wub = -4.972273e-25
+ wuc = -6.632247e-17
+ wwl = 0.0
+ wwn = 1.0
+ wmin = 5e-7
+ xti = 3
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0017857137
+ lkt1 = 6.187276e-9
+ lkt2 = 2.5314804e-9
+ pdiblcb = 0.01
+ weta0 = 0
+ lmax = 1.2e-6
+ lmin = 5e-7
+ wvsat = 0.0
+ lpclm = 1.4785714e-7
+ wvth0 = 1.4777807e-8
+ lpdiblc2 = 3.696429e-9
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ binunit = 2
+ pscbe1 = 349999900.0
+ pscbe2 = 5e-7
+ wub1 = -7.465372e-26
+ wuc1 = 1.5870021e-17
+ hdif = 2e-7
+ lub1 = -1.133461e-25
+ luc1 = -2.2106738e-17
+ wute = 7.883313e-8
+ mjsw = 0.3683619
+ nqsmod = 0
+ tpbswg = 0.001572025
+ noimod = 2
+ lute = 1.0183292e-7
+ lketa = -9.893122e-9
+ xpart = 1
+ cdsc = 0.0
+ cgdo = 3.28e-10
+ pbswg = 0.895226
+ version = 3.24
+ )

.model pch_tt_12 pmos (
+ level = 49
+ wint = 5e-9
+ llc = -0.039
+ pute = 1.3160581e-15
+ lln = -1
+ lu0 = 2.1198607e-10
+ vth0 = -0.4463558
+ nfactor = 1.0
+ lua = 2.3815556e-17
+ lub = -3.425063e-26
+ luc = 8.803578e-18
+ nch = 3.9e+17
+ rdsw = 530.0
+ lwl = 0.0
+ lwn = 1.0
+ pketa = -9.609158e-16
+ wkt1 = 2.7434011e-10
+ wkt2 = -6.113567e-9
+ lint = 1.4999999e-8
+ pa0 = -8.476619e-14
+ nlx = 0.0
+ wmax = 1.2e-6
+ pk1 = 1.5213101e-14
+ pk2 = -6.235986e-15
+ wmin = 5e-7
+ lkt1 = -4.083267e-9
+ lkt2 = -2.4314675e-9
+ wpclm = 5.671285e-8
+ pu0 = -1.4287007e-16
+ lmax = 5e-7
+ prt = 0
+ pua = -7.799214e-23
+ pub = 7.065072e-32
+ puc = 3.297807e-24
+ lmin = 1.8e-7
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.009150297
+ tcjsw = 0.0004130718
+ pdiblcb = 0.01
+ rsh = 7.2
+ tcj = 0.0009739001
+ ua1 = 1.224e-9
+ ub1 = -1.6175756e-18
+ uc1 = -2.2818641e-11
+ pvoff = -1.4343533e-15
+ tcjswg = 0.0004130718
+ tpb = 0.001572025
+ tox = 4.08e-9
+ a0 = 0.5166956
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ wa0 = 4.821862e-7
+ at = 10000.0
+ cf = 0
+ cj = 0.001121
+ wub1 = 8.30214e-26
+ ute = -0.5812994
+ wuc1 = 7.530186e-17
+ ef = 1.064
+ k1 = 0.7171482
+ k2 = -0.027492139
+ k3 = 0.0
+ em = 30000000.0
+ wk1 = -1.1417325e-7
+ wk2 = 3.837703e-8
+ binunit = 2
+ cdscb = 0.0
+ cdscd = -5.200001e-5
+ peta0 = 3.0000000000000003e-21
+ js = 2.5e-7
+ ll = 0.0
+ mj = 0.4476
+ hdif = 2e-7
+ lw = 0.0
+ u0 = 0.006858335
+ wln = 1.0
+ pb = 0.895226
+ w0 = 0.0
+ wu0 = 9.229584e-10
+ rd = 0
+ rs = 0
+ ua = -7.336427e-11
+ ub = 1.4258127e-18
+ uc = -5.946296e-11
+ lub1 = 6.724484e-26
+ wua = 5.726523e-16
+ wub = -7.845651e-25
+ wuc = -1.0188386e-16
+ wl = 0.0
+ luc1 = 7.110234e-18
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ wwl = 0.0
+ wwn = 1.0
+ wute = -5.584022e-8
+ wketa = 5.255423e-9
+ mjsw = 0.3683619
+ pvth0 = -1.0352502e-15
+ xti = 3
+ drout = 0.0
+ tpbsw = 0.001572025
+ lute = 7.748556e-9
+ wcdscd = -2.0304376e-11
+ cjswg = 4.221e-10
+ mjswg = 0.3683619
+ cdsc = 0.0
+ wvoff = 2.8364715e-9
+ cgdo = 3.28e-10
+ pcdscd = 9.13697e-18
+ cgso = 3.28e-10
+ weta0 = 0
+ version = 3.24
+ wvsat = 0.0
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ lpclm = 6.365384e-8
+ wvth0 = 5.738565e-9
+ cjsw = 2.481e-10
+ pscbe1 = 350000000.0
+ pscbe2 = 5e-7
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ nqsmod = 0
+ tpbswg = 0.001572025
+ tnom = 25.0
+ pnfactor = 0
+ noimod = 2
+ pags = -5.667374e-15
+ wnfactor = 0.0
+ toxm = 4.08e-9
+ pcit = 2.6834248e-18
+ pbsw = 0.895226
+ lketa = -1.8239428e-9
+ pclm = 0.858547
+ xpart = 1
+ ppdiblc2 = 7.08422e-16
+ wpdiblc2 = -1.5742713e-9
+ lnfactor = 0.0
+ pbswg = 0.895226
+ lcdscd = 2.3400004e-11
+ lvoff = -3.0382863e-10
+ ags = 0.010547621
+ beta0 = 22.67827
+ pkt1 = 8.196091e-17
+ pkt2 = 1.5372367e-15
+ keta = 0.01791114
+ lpdiblc2 = 3.823661e-10
+ leta0 = 2.5596747e-10
+ capmod = 3
+ letab = -3.473438e-10
+ cit = 0.00012746976
+ wags = 1.2594167e-8
+ lvsat = -0.0003656142
+ dsub = 0.0
+ dlc = 2e-9
+ lvth0 = -8.202719e-9
+ k3b = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ lags = 4.253569e-9
+ wcit = -2.0641719e-11
+ ppclm = -2.5520774e-14
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ delta = 0.01
+ mobmod = 1
+ lcit = 4.881893e-11
+ voff = -0.1286711
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ ldif = 9e-8
+ kt1l = 0.0
+ prwb = 0.0
+ pub1 = -2.1229706e-32
+ prwg = 0.0
+ puc1 = -9.461855e-24
+ la0 = 1.6783336e-7
+ eta0 = -0.00046875
+ pvag = 0.0
+ jsw = 1.2e-12
+ etab = 0.0006718753
+ kt1 = -0.2211471
+ lk1 = -8.844278e-9
+ kt2 = -0.014824204
+ lk2 = 4.904499e-9
+ vsat = 130812.46
+ )

.model pch_tt_13 pmos (
+ level = 49
+ wketa = -6.403492e-9
+ pvth0 = 0.0
+ drout = 0.0
+ toxm = 4.08e-9
+ tpbsw = 0.001572025
+ pbsw = 0.895226
+ pclm = 0.5999999
+ cjswg = 4.221e-10
+ mjswg = 0.3683619
+ wvoff = -1.320298e-9
+ weta0 = 0
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ wvsat = 0.0
+ keta = 0.04310941
+ pscbe1 = 199999970.0
+ pscbe2 = 5e-7
+ wvth0 = 9.340613e-9
+ dsub = 0.0
+ nqsmod = 0
+ tpbswg = 0.001572025
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ noimod = 2
+ voff = -0.1261533
+ ldif = 9e-8
+ a0 = 0.8704194
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ at = 10000.0
+ cf = 0
+ cj = 0.001121
+ ef = 1.064
+ k1 = 0.5421249
+ k2 = 0.03567642
+ k3 = 0.0
+ em = 30000000.0
+ ags = 0.02
+ eta0 = 5e-5
+ js = 2.5e-7
+ ll = 0.0
+ mj = 0.4476
+ lw = 0.0
+ pvag = 0.0
+ etab = -5e-5
+ u0 = 0.009748334
+ pb = 0.895226
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ vsat = 149999.98
+ xpart = 1
+ ua = 1.2584637e-9
+ ub = 4.999999e-20
+ uc = -1.6065008e-10
+ wint = 5e-9
+ wl = 0.0
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ cit = -0.0001
+ vth0 = -0.4484667
+ rdsw = 530.0
+ dlc = 2e-9
+ wkt1 = 3.830554e-9
+ wkt2 = 1.9527771e-9
+ k3b = 0.0
+ lint = 1.4999999e-8
+ pbswg = 0.895226
+ dwb = 0.0
+ wmax = 5e-7
+ dwg = 0.0
+ nfactor = 1.0
+ wmin = 2.2e-7
+ lvoff = 0.0
+ lmax = 2.0001e-5
+ lmin = 1e-5
+ capmod = 3
+ beta0 = 22.67827
+ leta0 = 3e-14
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.001
+ pdiblcb = 0.01
+ jsw = 1.2e-12
+ kt1 = -0.2247607
+ kt2 = -0.027069092
+ lk2 = 0.0
+ lvth0 = 0.0
+ llc = -0.039
+ lln = -1
+ lu0 = 0.0
+ wub1 = 2.1644123e-27
+ wuc1 = -1.2526765e-17
+ nch = 3.9e+17
+ mobmod = 1
+ lwl = 0.0
+ lwn = 1.0
+ delta = 0.01
+ hdif = 2e-7
+ nlx = 0.0
+ pnfactor = 0
+ binunit = 2
+ wute = 6.898109e-9
+ mjsw = 0.3683619
+ wnfactor = 0.0
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ pu0 = 0.0
+ prt = 0
+ rsh = 7.2
+ tcj = 0.0009739001
+ ua1 = 1.224e-9
+ ub1 = -1.3041941e-18
+ uc1 = 6.665171e-11
+ cdsc = 0.0
+ tpb = 0.001572025
+ tox = 4.08e-9
+ wa0 = 8.951166e-8
+ lnfactor = 0.0
+ cgdo = 3.28e-10
+ ute = -0.7678431
+ wk1 = 3.561511e-9
+ wk2 = -4.719829e-9
+ wln = 1.0
+ cgso = 3.28e-10
+ wu0 = -4.034686e-11
+ wua = -2.3131395e-16
+ wuc = -1.2695932e-17
+ wwl = 0.0
+ wwn = 1.0
+ xti = 3
+ tcjsw = 0.0004130718
+ tcjswg = 0.0004130718
+ version = 3.24
+ cjsw = 2.481e-10
+ pvoff = 0.0
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 3.0000000000000003e-21
+ tnom = 25.0
+ )

.model pch_tt_14 pmos (
+ level = 49
+ tpbswg = 0.001572025
+ noimod = 2
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0004772729
+ cit = -0.0001
+ wub1 = -3.0198158e-27
+ wuc1 = -1.0513175e-17
+ pdiblcb = 0.01
+ lpscbe1 = 195.04262
+ dlc = 2e-9
+ hdif = 2e-7
+ k3b = 0.0
+ lub1 = -2.0820251e-25
+ dwb = 0.0
+ dwg = 0.0
+ luc1 = 9.921307e-17
+ wute = 1.1298283e-8
+ mjsw = 0.3683619
+ binunit = 2
+ lketa = -4.562476e-8
+ lute = 2.2927659e-7
+ xpart = 1
+ la0 = 5.081137e-7
+ cdsc = 0.0
+ jsw = 1.2e-12
+ kt1 = -0.2237138
+ lk1 = -4.88067e-8
+ kt2 = -0.026908273
+ lk2 = 2.3302198e-8
+ llc = -0.039
+ lln = -1
+ cgdo = 3.28e-10
+ lu0 = -3.0000519e-10
+ pbswg = 0.895226
+ lua = -3.24011e-17
+ lub = -3.941427e-28
+ luc = -6.882293e-17
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ cgso = 3.28e-10
+ pa0 = -1.854315e-13
+ lvoff = -2.3886029e-9
+ nlx = 0.0
+ capmod = 3
+ pk1 = 3.786126e-14
+ pk2 = -1.6169635e-14
+ beta0 = 22.67827
+ pu0 = -6.225135e-16
+ leta0 = 3e-14
+ prt = 0
+ pua = -1.3939852e-23
+ pub = 1.1764949e-34
+ puc = 1.4094153e-23
+ cjsw = 2.481e-10
+ lvsat = -0.013002842
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ lvth0 = -4.608335e-9
+ version = 3.24
+ rsh = 7.2
+ tcj = 0.0009739001
+ mobmod = 1
+ ua1 = 1.224e-9
+ ub1 = -1.2832692e-18
+ uc1 = 5.668055e-11
+ tpb = 0.001572025
+ tox = 4.08e-9
+ delta = 0.01
+ wa0 = 1.0814799e-7
+ tnom = 25.0
+ ute = -0.790886
+ wk1 = -2.4364055e-10
+ wk2 = -3.0947396e-9
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ wln = 1.0
+ wu0 = 2.2217313e-11
+ toxm = 4.08e-9
+ wua = -2.2991296e-16
+ wub = -1.1822094e-29
+ wuc = -1.4112429e-17
+ wwl = 0.0
+ wwn = 1.0
+ pbsw = 0.895226
+ xti = 3
+ pclm = 0.5738635
+ pketa = 1.7549415e-14
+ a0 = 0.8193527
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ at = 10000.0
+ cf = 0
+ cj = 0.001121
+ ef = 1.064
+ k1 = 0.5470301
+ k2 = 0.03333449
+ k3 = 0.0
+ em = 30000000.0
+ js = 2.5e-7
+ ll = 0.0
+ mj = 0.4476
+ lw = 0.0
+ u0 = 0.009778486
+ pb = 0.895226
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ua = 1.2617201e-9
+ ub = 5.00396e-20
+ uc = -1.5373321e-10
+ wl = 0.0
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -2e-8
+ ww = 0.0
+ tcjswg = 0.0004130718
+ xw = 0.0
+ tcjsw = 0.0004130718
+ pkt1 = 2.5501714e-15
+ pkt2 = -4.817884e-16
+ keta = 0.04769481
+ pvoff = 2.6840621e-15
+ dsub = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 3.0000000000000003e-21
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ pnfactor = 0
+ wketa = -8.167253e-9
+ pvth0 = -3.640382e-15
+ wnfactor = 0.0
+ voff = -0.1259132
+ drout = 0.0
+ ldif = 9e-8
+ tpbsw = 0.001572025
+ kt1l = 0.0
+ prwb = 0.0
+ pub1 = 5.158311e-32
+ prwg = 0.0
+ puc1 = -2.0035212e-23
+ eta0 = 5e-5
+ cjswg = 4.221e-10
+ pvag = 0.0
+ etab = -5e-5
+ vsat = 151306.8
+ mjswg = 0.3683619
+ wint = 5e-9
+ pute = -4.378173e-14
+ vth0 = -0.4480035
+ rdsw = 530.0
+ lnfactor = 0.0
+ wvoff = -1.590053e-9
+ wkt1 = 3.574256e-9
+ wkt2 = 2.0011981e-9
+ lint = 1.4999999e-8
+ wmax = 5e-7
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ wmin = 2.2e-7
+ lkt1 = -1.0417262e-8
+ lkt2 = -1.6001408e-9
+ weta0 = 0
+ nfactor = 1.0
+ lmax = 1e-5
+ pscbe1 = 180397700.0
+ pscbe2 = 5e-7
+ wvsat = 0.0
+ lmin = 1.2e-6
+ lpclm = 2.6005691e-7
+ wvth0 = 9.70648e-9
+ lpdiblc2 = 5.201136e-9
+ ags = 0.02
+ nqsmod = 0
+ )

.model pch_tt_15 pmos (
+ level = 49
+ ute = -0.5904401
+ wk1 = 4.182789e-8
+ wk2 = -2.2085489e-8
+ beta0 = 22.67827
+ wln = 1.0
+ wu0 = -3.987341e-10
+ pkt1 = -8.599671e-15
+ pkt2 = 1.9347028e-16
+ lpdiblc2 = 3.696429e-9
+ keta = 0.0004484208
+ wua = -1.9008923e-16
+ leta0 = 3.699428e-11
+ wub = 8.369847e-27
+ wuc = 5.370726e-18
+ wwl = 0.0
+ wwn = 1.0
+ letab = -3.696428e-11
+ xti = 3
+ mobmod = 1
+ lvsat = -0.007392816
+ dsub = 0.0
+ lvth0 = -1.5532533e-8
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ delta = 0.01
+ lcit = 2.2622144e-10
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ voff = -0.1186655
+ ldif = 9e-8
+ kt1l = 0.0
+ prwb = 0.0
+ pub1 = -1.2589071e-33
+ prwg = 0.0
+ puc1 = 4.27717e-24
+ eta0 = 1.7857146e-5
+ pvag = 0.0
+ etab = -1.7857146e-5
+ vsat = 146428.52
+ wint = 5e-9
+ pute = -8.783067e-15
+ vth0 = -0.4385042
+ rdsw = 530.0
+ pketa = -5.090041e-15
+ wkt1 = 1.3269771e-8
+ wkt2 = 1.4140165e-9
+ lint = 1.4999999e-8
+ wmax = 5e-7
+ tcjswg = 0.0004130718
+ wmin = 2.2e-7
+ lkt1 = 1.1386779e-8
+ lkt2 = -8.841858e-10
+ lmax = 1.2e-6
+ lmin = 5e-7
+ tcjsw = 0.0004130718
+ nfactor = 1.0
+ pvoff = 3.95383e-15
+ wub1 = 4.292976e-26
+ cdscb = 0.0
+ wuc1 = -3.165437e-17
+ cdscd = 0.0
+ peta0 = 3.0000000000000003e-21
+ hdif = 2e-7
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0017857139
+ pdiblcb = 0.01
+ lub1 = -9.299159e-27
+ wketa = 1.1519229e-8
+ luc1 = 4.434689e-18
+ pvth0 = 7.623086e-16
+ wute = -1.9135335e-8
+ mjsw = 0.3683619
+ drout = 0.0
+ tpbsw = 0.001572025
+ lute = -1.2362289e-9
+ cjswg = 4.221e-10
+ binunit = 2
+ mjswg = 0.3683619
+ ags = 0.02
+ cdsc = 0.0
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ wvoff = -2.6941984e-9
+ cit = -0.00029671428
+ cgdo = 3.28e-10
+ pscbe1 = 349999900.0
+ pscbe2 = 5e-7
+ dlc = 2e-9
+ cgso = 3.28e-10
+ k3b = 0.0
+ weta0 = 0
+ dwb = 0.0
+ dwg = 0.0
+ wvsat = 0.0
+ lpclm = 1.4785714e-7
+ wvth0 = 5.878054e-9
+ nqsmod = 0
+ a0 = 1.1508681
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ tpbswg = 0.001572025
+ cjsw = 2.481e-10
+ noimod = 2
+ at = 10000.0
+ cf = 0
+ cj = 0.001121
+ ef = 1.064
+ k1 = 0.510219
+ k2 = 0.05410628
+ k3 = 0.0
+ em = 30000000.0
+ js = 2.5e-7
+ ll = 0.0
+ noia = 9.5e+18
+ mj = 0.4476
+ noib = 100000.0
+ noic = 1.4e-12
+ lw = 0.0
+ u0 = 0.009203287
+ pb = 0.895226
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ua = 1.0922192e-9
+ ub = 2.0536515e-20
+ uc = -2.183638e-10
+ la0 = 1.2687106e-7
+ wl = 0.0
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ jsw = 1.2e-12
+ version = 3.24
+ kt1 = -0.2426738
+ lk1 = -6.473878e-9
+ kt2 = -0.027530843
+ lk2 = -5.853628e-10
+ llc = -0.039
+ lln = -1
+ pnfactor = 0
+ lu0 = 3.614737e-10
+ tnom = 25.0
+ lua = 1.6252487e-16
+ lub = 3.353441e-26
+ luc = 5.502275e-18
+ nch = 3.9e+17
+ wnfactor = 0.0
+ lwl = 0.0
+ lwn = 1.0
+ pa0 = 5.971399e-14
+ nlx = 0.0
+ toxm = 4.08e-9
+ lketa = 8.708591e-9
+ pk1 = -1.0521005e-14
+ pk2 = 5.669729e-15
+ pbsw = 0.895226
+ pclm = 0.6714286
+ pu0 = -1.384194e-16
+ xpart = 1
+ prt = 0
+ pua = -5.973716e-23
+ pub = -9.521269e-33
+ puc = -8.311478e-24
+ rsh = 7.2
+ lnfactor = 0.0
+ tcj = 0.0009739001
+ ua1 = 1.224e-9
+ ub1 = -1.4562286e-18
+ uc1 = 1.3909653e-10
+ pbswg = 0.895226
+ capmod = 3
+ tpb = 0.001572025
+ tox = 4.08e-9
+ wa0 = -1.0502199e-7
+ lvoff = -1.0723419e-8
+ )

.model pch_tt_16 pmos (
+ level = 49
+ cdsc = 0.0
+ binunit = 2
+ pketa = 7.45672e-16
+ lnfactor = 0.0
+ tcjswg = 0.0004130718
+ cgdo = 3.28e-10
+ wpclm = 4.634222e-9
+ cgso = 3.28e-10
+ tcjsw = 0.0004130718
+ lpdiblc2 = 1.8281252e-9
+ cjsw = 2.481e-10
+ pvoff = 1.4541431e-15
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ wcdscd = -1.4183201e-11
+ ags = 0.03625
+ cdscb = 0.0
+ cdscd = -6.449223e-5
+ peta0 = 3.0000000000000003e-21
+ cit = 8.534377e-5
+ tnom = 25.0
+ wketa = -1.4490222e-9
+ pvth0 = -2.8414808e-16
+ version = 3.24
+ dlc = 2e-9
+ drout = 0.0
+ pcdscd = 6.382441e-18
+ tpbsw = 0.001572025
+ k3b = 0.0
+ toxm = 4.08e-9
+ dwb = 0.0
+ dwg = 0.0
+ pbsw = 0.895226
+ pclm = 0.9648299
+ cjswg = 4.221e-10
+ mjswg = 0.3683619
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ wvoff = 2.8606606e-9
+ pscbe1 = 350000000.0
+ pscbe2 = 5e-7
+ la0 = 7.233052e-9
+ jsw = 1.2e-12
+ kt1 = -0.2130934
+ lk1 = 1.3789155e-8
+ kt2 = -0.03589084
+ lk2 = -3.106946e-9
+ llc = -0.039
+ weta0 = 0
+ lln = -1
+ lu0 = -3.566262e-10
+ nqsmod = 0
+ lua = -2.6402067e-16
+ lub = 2.6345733e-25
+ luc = 3.340897e-17
+ nch = 3.9e+17
+ wvsat = 0.0
+ tpbswg = 0.001572025
+ lwl = 0.0
+ lwn = 1.0
+ noimod = 2
+ lpclm = 1.5826547e-8
+ pa0 = -6.072043e-15
+ wvth0 = 8.203513e-9
+ nlx = 0.0
+ pkt1 = -9.758805e-16
+ pkt2 = -1.0643102e-15
+ keta = 0.03159368
+ pk1 = 4.122718e-15
+ pk2 = -2.3103772e-15
+ dsub = 0.0
+ pu0 = 1.3574996e-16
+ prt = 0
+ pua = 6.304761e-23
+ pub = -7.522618e-32
+ puc = -8.758834e-24
+ lags = -7.312499e-9
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ rsh = 7.2
+ tcj = 0.0009739001
+ ua1 = 1.224e-9
+ ub1 = -1.4433942e-18
+ uc1 = 2.0396977e-10
+ tpb = 0.001572025
+ tox = 4.08e-9
+ lcit = 5.429531e-11
+ voff = -0.1287204
+ wa0 = 4.116919e-8
+ lcdscd = 2.9021494e-11
+ ldif = 9e-8
+ ute = -0.5893072
+ wk1 = 9.286284e-9
+ kt1l = 0.0
+ wk2 = -4.351921e-9
+ prwb = 0.0
+ pub1 = 1.9106841e-32
+ prwg = 0.0
+ lketa = -5.306775e-9
+ puc1 = 6.153712e-24
+ wln = 1.0
+ wu0 = -1.0079994e-9
+ eta0 = -0.0004687502
+ wua = -4.629443e-16
+ pvag = 0.0
+ wub = 1.5438073e-25
+ wuc = 6.364847e-18
+ etab = 0.0006718753
+ xpart = 1
+ wwl = 0.0
+ wwn = 1.0
+ vsat = 130812.55
+ xti = 3
+ wint = 5e-9
+ pute = 5.968411e-15
+ vth0 = -0.4513863
+ capmod = 3
+ rdsw = 530.0
+ wkt1 = -3.671987e-9
+ wkt2 = 4.209085e-9
+ pbswg = 0.895226
+ lint = 1.4999999e-8
+ wmax = 5e-7
+ wmin = 2.2e-7
+ lvoff = -6.198719e-9
+ lkt1 = -1.9244071e-9
+ lkt2 = 2.877812e-9
+ lmax = 5e-7
+ beta0 = 22.67827
+ lmin = 1.8e-7
+ mobmod = 1
+ leta0 = 2.5596758e-10
+ letab = -3.473438e-10
+ lvsat = -0.0003656336
+ nfactor = 1.0
+ lvth0 = -9.735581e-9
+ ppclm = -2.0853998e-15
+ wub1 = -2.3274574e-27
+ wuc1 = -3.582447e-17
+ delta = 0.01
+ hdif = 2e-7
+ a0 = 1.4167303
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ pnfactor = 0
+ lub1 = -1.5074642e-26
+ luc1 = -2.4758267e-17
+ at = 10000.0
+ cf = 0
+ cj = 0.001121
+ ef = 1.064
+ k1 = 0.46519
+ dvt0w = 0.0
+ k2 = 0.0597098
+ k3 = 0.0
+ em = 30000000.0
+ wnfactor = 0.0
+ wute = -5.191639e-8
+ dvt1w = 0.0
+ dvt2w = 0.0
+ mjsw = 0.3683619
+ js = 2.5e-7
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.005937499
+ ll = 0.0
+ mj = 0.4476
+ lw = 0.0
+ u0 = 0.010799064
+ pb = 0.895226
+ w0 = 0.0
+ rd = 0
+ pdiblcb = 0.01
+ rs = 0
+ ua = 2.0400983e-9
+ ub = -4.904033e-19
+ uc = -2.8037866e-10
+ wl = 0.0
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -2e-8
+ ww = 0.0
+ lute = -1.7460413e-9
+ xw = 0.0
+ )

.model pch_fs_1 pmos (
+ level = 49
+ lvth0 = -3.9543e-9
+ cdsc = 0.0
+ binunit = 2
+ pnfactor = 0
+ cgdo = 3.28e-10
+ delta = 0.01
+ wnfactor = 0.0
+ cgso = 3.28e-10
+ dvt0w = 0.0
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ dvt1w = 0.0
+ dvt2w = 0.0
+ pscbe1 = 199999970.0
+ pscbe2 = 5e-7
+ cjsw = 2.60505e-10
+ ags = 0.02
+ lnfactor = -3.9543e-9
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ nqsmod = 0
+ tpbswg = 0.001572025
+ noimod = 2
+ cit = -0.0001
+ dlc = 2e-9
+ tnom = 25.0
+ version = 3.24
+ k3b = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ toxm = 4.08e-9
+ tcjsw = 0.0004130718
+ pbsw = 0.895226
+ pclm = 0.6000001
+ pvoff = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ jsw = 1.2e-12
+ peta0 = 1.8966694548261387e-25
+ kt1 = -0.2311294
+ lk2 = 1.18629e-9
+ kt2 = -0.02433992
+ llc = -0.039
+ lln = -1
+ lu0 = -7.9086e-11
+ nch = 3.9e+17
+ pvth0 = -1.18629e-15
+ lwl = 0.0
+ lwn = 1.0
+ drout = 0.0
+ nlx = 0.0
+ tpbsw = 0.001572025
+ capmod = 3
+ keta = 0.026632193
+ pu0 = 0.0
+ cjswg = 4.43205e-10
+ prt = 0
+ dsub = 0.0
+ mjswg = 0.3683619
+ rsh = 7.2
+ tcj = 0.0009739001
+ ua1 = 1.224e-9
+ ub1 = -1.3928839e-18
+ uc1 = -4.59467e-12
+ wvoff = 0.0
+ mobmod = 1
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ tpb = 0.001572025
+ tox = 4.08e-9
+ ute = -0.8288856
+ voff = -0.1275921
+ weta0 = 0
+ ldif = 9e-8
+ wvsat = 0.0
+ wln = 1.0
+ kt1l = 0.0
+ prwb = 0.0
+ wu0 = -1.97715e-11
+ prwg = 0.0
+ wvth0 = -1.18629e-9
+ wwl = 0.0
+ wwn = 1.0
+ eta0 = 5e-5
+ xti = 3
+ pvag = 0.0
+ etab = -5e-5
+ vsat = 149999.98
+ wint = 5e-9
+ vth0 = -0.46220690000000003
+ rdsw = 530.0
+ lint = 1.4999999e-8
+ wmax = 0.000900001
+ wmin = 1e-5
+ a0 = 1.0461572
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ lmax = 2.0001e-5
+ at = 10000.0
+ cf = 0
+ cj = 0.00117705
+ lmin = 1e-5
+ ef = 1.064
+ k1 = 0.5375325
+ k2 = 0.04056858
+ k3 = 0.0
+ em = 30000000.0
+ tcjswg = 0.0004130718
+ js = 2.5e-7
+ ll = 0.0
+ mj = 0.4476
+ lw = 0.0
+ u0 = 0.0108097578
+ pb = 0.895226
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ua = 8.23294e-10
+ ub = 6.854322e-19
+ uc = -8.655411e-11
+ wl = 0.0
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ xpart = 1
+ nfactor = 1.0
+ pbswg = 0.895226
+ hdif = 2e-7
+ lvoff = -1.5817200000000002e-9
+ mjsw = 0.3683619
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0010000003
+ pdiblcb = 0.01
+ beta0 = 22.67827
+ leta0 = 1.8966694548261387e-18
+ )

.model pch_fs_2 pmos (
+ level = 49
+ mj = 0.4476
+ lw = 0.0
+ kt1 = -0.2295883
+ lk1 = 1.8783622e-8
+ kt2 = -0.024031118
+ lk2 = -4.300882e-9
+ u0 = 0.0109398048
+ pb = 0.895226
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ua = 8.625313e-10
+ ub = 6.401998e-19
+ uc = -8.855145e-11
+ llc = -0.039
+ lln = -1
+ wl = 0.0
+ lu0 = -1.3730549e-9
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ voff = -0.1274002
+ lua = -3.904111e-16
+ lub = 4.500626e-25
+ luc = 1.9873557e-17
+ ldif = 9e-8
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ kt1l = 0.0
+ tcjsw = 0.0004130718
+ prwb = 0.0
+ prwg = 0.0
+ nlx = 0.0
+ eta0 = 5e-5
+ pvag = 0.0
+ etab = -5e-5
+ pvoff = 0.0
+ vsat = 151306.8
+ pu0 = 0.0
+ wint = 5e-9
+ prt = 0
+ vth0 = -0.45971300000000004
+ rdsw = 530.0
+ pnfactor = 0
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 1.8966694548261387e-25
+ lint = 1.4999999e-8
+ rsh = 7.2
+ tcj = 0.0009739001
+ ua1 = 1.224e-9
+ wnfactor = 0.0
+ wmax = 0.000900001
+ ub1 = -1.3977103e-18
+ uc1 = -6.694918e-12
+ wmin = 1e-5
+ tpb = 0.001572025
+ capmod = 3
+ pvth0 = -1.18629e-15
+ tox = 4.08e-9
+ lkt1 = -1.5333228e-8
+ lkt2 = -3.0725886e-9
+ drout = 0.0
+ lmax = 1e-5
+ tpbsw = 0.001572025
+ ute = -0.8385549
+ lmin = 1.2e-6
+ wln = 1.0
+ wu0 = -1.97715e-11
+ cjswg = 4.43205e-10
+ wwl = 0.0
+ wwn = 1.0
+ mjswg = 0.3683619
+ lnfactor = -3.9543e-9
+ xti = 3
+ mobmod = 1
+ nfactor = 1.0
+ wvoff = 0.0
+ hdif = 2e-7
+ lub1 = 4.802326e-26
+ luc1 = 2.0897466e-17
+ weta0 = 0
+ mjsw = 0.3683619
+ lpdiblc2 = 5.201137e-9
+ wvsat = 0.0
+ lute = 9.620972e-8
+ lpclm = 2.6005682e-7
+ wvth0 = -1.18629e-9
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0004772727
+ pdiblcb = 0.01
+ lpscbe1 = 195.04263
+ cdsc = 0.0
+ cgdo = 3.28e-10
+ binunit = 2
+ cgso = 3.28e-10
+ tcjswg = 0.0004130718
+ lketa = -2.0462676e-9
+ cjsw = 2.60505e-10
+ xpart = 1
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ pbswg = 0.895226
+ tnom = 25.0
+ lvoff = -3.4908509e-9
+ toxm = 4.08e-9
+ beta0 = 22.67827
+ version = 3.24
+ pbsw = 0.895226
+ pclm = 0.5738637
+ leta0 = 1.8966694548261387e-18
+ lvsat = -0.013002843
+ lvth0 = -2.8768353e-8
+ ags = 0.02
+ delta = 0.01
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ cit = -0.0001
+ dlc = 2e-9
+ dvt0w = 0.0
+ dvt1w = 0.0
+ pscbe1 = 180397680.0
+ pscbe2 = 5e-7
+ dvt2w = 0.0
+ k3b = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ keta = 0.026837848
+ nqsmod = 0
+ tpbswg = 0.001572025
+ dsub = 0.0
+ noimod = 2
+ a0 = 1.0385712
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ at = 10000.0
+ cf = 0
+ cj = 0.00117705
+ la0 = 7.548124e-8
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ ef = 1.064
+ k1 = 0.5356447
+ k2 = 0.041120050000000005
+ k3 = 0.0
+ em = 30000000.0
+ js = 2.5e-7
+ jsw = 1.2e-12
+ ll = 0.0
+ )

.model pch_fs_3 pmos (
+ level = 49
+ cjswg = 4.43205e-10
+ mjswg = 0.3683619
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ wvoff = 0.0
+ tnom = 25.0
+ weta0 = 0
+ wvsat = 0.0
+ toxm = 4.08e-9
+ a0 = 1.0045335
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ lpclm = 1.4785704e-7
+ wvth0 = -1.18629e-9
+ pbsw = 0.895226
+ pclm = 0.6714287
+ at = 10000.0
+ cf = 0
+ cj = 0.00117705
+ ef = 1.064
+ k1 = 0.5405614
+ k2 = 0.04043759
+ k3 = 0.0
+ em = 30000000.0
+ js = 2.5e-7
+ version = 3.24
+ ll = 0.0
+ mj = 0.4476
+ lw = 0.0
+ u0 = 0.0101692238
+ pb = 0.895226
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ua = 5.26694e-10
+ ub = 1.1734415e-18
+ uc = -4.332115e-11
+ wl = 0.0
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ pnfactor = 0
+ wnfactor = 0.0
+ tcjswg = 0.0004130718
+ lketa = -8.158225e-9
+ keta = 0.03215259
+ xpart = 1
+ dsub = 0.0
+ lnfactor = -3.9543e-9
+ ags = 0.02
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ pbswg = 0.895226
+ lvoff = -2.5305025000000003e-9
+ lcit = 2.2402701e-10
+ cit = -0.00029480609
+ voff = -0.1282353
+ lpdiblc2 = 3.696428e-9
+ ldif = 9e-8
+ dlc = 2e-9
+ beta0 = 22.67827
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ k3b = 0.0
+ dwb = 0.0
+ leta0 = 3.6964281896669455e-11
+ dwg = 0.0
+ eta0 = 1.7857143e-5
+ letab = -3.696428e-11
+ pvag = 0.0
+ etab = -1.7857143e-5
+ lvsat = -0.007392833
+ vsat = 146428.53
+ wint = 5e-9
+ lvth0 = -1.0643742e-8
+ vth0 = -0.4754736
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ rdsw = 530.0
+ delta = 0.01
+ lint = 1.4999999e-8
+ wmax = 0.000900001
+ pscbe1 = 349999900.0
+ pscbe2 = 5e-7
+ la0 = 1.146246e-7
+ wmin = 1e-5
+ jsw = 1.2e-12
+ lkt1 = 1.5747348e-9
+ lkt2 = 9.740028e-10
+ kt1 = -0.2442909
+ lk1 = 1.3129389e-8
+ kt2 = -0.027549893
+ lk2 = -3.5160449999999997e-9
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ lmax = 1.2e-6
+ llc = -0.039
+ lln = -1
+ lu0 = -4.868866e-10
+ lmin = 5e-7
+ lua = -4.198125e-18
+ lub = -1.631654e-25
+ luc = -3.214129e-17
+ nch = 3.9e+17
+ nqsmod = 0
+ lwl = 0.0
+ lwn = 1.0
+ tpbswg = 0.001572025
+ noimod = 2
+ nlx = 0.0
+ pu0 = 0.0
+ prt = 0
+ hdif = 2e-7
+ rsh = 7.2
+ tcj = 0.0009739001
+ nfactor = 1.0
+ ua1 = 1.224e-9
+ lub1 = 3.0810812e-26
+ ub1 = -1.3827429e-18
+ luc1 = 2.9752128e-17
+ uc1 = -1.4394627e-11
+ mjsw = 0.3683619
+ tpb = 0.001572025
+ tox = 4.08e-9
+ tcjsw = 0.0004130718
+ lute = 3.654092e-8
+ ute = -0.786669
+ wln = 1.0
+ pvoff = 0.0
+ wu0 = -1.97715e-11
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0017857148
+ wwl = 0.0
+ wwn = 1.0
+ pdiblcb = 0.01
+ cdsc = 0.0
+ xti = 3
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 1.8966694548261387e-25
+ capmod = 3
+ cgdo = 3.28e-10
+ pvth0 = -1.18629e-15
+ cgso = 3.28e-10
+ drout = 0.0
+ binunit = 2
+ tpbsw = 0.001572025
+ cjsw = 2.60505e-10
+ mobmod = 1
+ )

.model pch_fs_4 pmos (
+ level = 49
+ wmin = 1e-5
+ lkt1 = -2.665e-9
+ lkt2 = -2.325577e-10
+ lmax = 5e-7
+ cit = -4.054396e-5
+ lmin = 1.8e-7
+ lketa = -8.307595e-10
+ dlc = 2e-9
+ k3b = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ xpart = 1
+ pbswg = 0.895226
+ hdif = 2e-7
+ lub1 = 2.883988e-26
+ luc1 = -6.846759e-18
+ lvoff = -1.6174359200000002e-9
+ la0 = 1.6196543e-8
+ mjsw = 0.3683619
+ jsw = 1.2e-12
+ kt1 = -0.2348693
+ lk1 = 1.6807924e-8
+ kt2 = -0.024868647
+ lk2 = -4.689925e-9
+ beta0 = 22.67827
+ nfactor = 1.0
+ llc = -0.039
+ lln = -1
+ lu0 = -1.7803381e-10
+ lute = 1.6013461e-9
+ leta0 = 2.559375218966695e-10
+ lua = -1.5999061e-16
+ lub = 1.2197973e-25
+ luc = 1.8500639e-17
+ nch = 3.9e+17
+ letab = -5.298917e-10
+ lwl = 0.0
+ lwn = 1.0
+ lvsat = -0.0003656265
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ nlx = 0.0
+ lvth0 = -1.2194852e-8
+ cdsc = 0.0
+ pscbe1 = 350000000.0
+ pscbe2 = 5e-7
+ pnfactor = 0
+ pu0 = 0.0
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.00796875
+ delta = 0.01
+ a0 = 1.2232625
+ a1 = 0.0
+ a2 = 0.4
+ prt = 0
+ b0 = 0.0
+ b1 = 0.0
+ cgdo = 3.28e-10
+ wnfactor = 0.0
+ pdiblcb = 0.01
+ at = 10000.0
+ cf = 0
+ cj = 0.00117705
+ ef = 1.064
+ k1 = 0.5323869
+ k2 = 0.04304621
+ k3 = 0.0
+ em = 30000000.0
+ cgso = 3.28e-10
+ js = 2.5e-7
+ dvt0w = 0.0
+ dvt1w = 0.0
+ ll = 0.0
+ rsh = 7.2
+ mj = 0.4476
+ dvt2w = 0.0
+ lw = 0.0
+ u0 = 0.0094828838
+ tcj = 0.0009739001
+ nqsmod = 0
+ pb = 0.895226
+ ua1 = 1.224e-9
+ w0 = 0.0
+ ub1 = -1.3783631e-18
+ rd = 0
+ uc1 = 6.693623e-11
+ tpbswg = 0.001572025
+ rs = 0
+ ua = 8.728995e-10
+ ub = 5.397856e-19
+ uc = -1.5585878e-10
+ noimod = 2
+ wl = 0.0
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ tpb = 0.001572025
+ tox = 4.08e-9
+ binunit = 2
+ cjsw = 2.60505e-10
+ ute = -0.7090256
+ lnfactor = -3.9543e-9
+ wln = 1.0
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ wu0 = -1.97715e-11
+ wwl = 0.0
+ wwn = 1.0
+ xti = 3
+ tnom = 25.0
+ lcdscd = 3.65625e-11
+ lpdiblc2 = 9.140626e-10
+ toxm = 4.08e-9
+ tcjsw = 0.0004130718
+ pbsw = 0.895226
+ pclm = 0.9102259
+ pvoff = 0.0
+ capmod = 3
+ version = 3.24
+ cdscb = 0.0
+ cdscd = -8.125e-5
+ peta0 = 1.8966694548261387e-25
+ pvth0 = -1.18629e-15
+ drout = 0.0
+ tpbsw = 0.001572025
+ mobmod = 1
+ keta = 0.015869336
+ cjswg = 4.43205e-10
+ mjswg = 0.3683619
+ dsub = 0.0
+ wvoff = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ weta0 = 0
+ lcit = 1.0960905e-10
+ voff = -0.1302643
+ ldif = 9e-8
+ wvsat = 0.0
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ lpclm = 4.03983e-8
+ wvth0 = -1.18629e-9
+ eta0 = -0.0004687502
+ pvag = 0.0
+ etab = 0.0010775371
+ vsat = 130812.52
+ wint = 5e-9
+ vth0 = -0.4720267
+ rdsw = 530.0
+ tcjswg = 0.0004130718
+ lint = 1.4999999e-8
+ wmax = 0.000900001
+ ags = 0.02
+ )

.model pch_fs_5 pmos (
+ level = 49
+ wa0 = -4.787191e-8
+ pscbe1 = 199999970.0
+ pscbe2 = 5e-7
+ ute = -0.8394966
+ lvth0 = -3.9543e-9
+ wk1 = 1.2456701e-8
+ wk2 = -5.940143e-9
+ wln = 1.0
+ wu0 = -1.2692462000000002e-9
+ delta = 0.01
+ wua = 1.7543858e-16
+ wub = -6.530953e-25
+ wuc = -7.950096e-17
+ wwl = 0.0
+ wwn = 1.0
+ nqsmod = 0
+ xti = 3
+ version = 3.24
+ tpbswg = 0.001572025
+ noimod = 2
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ keta = 0.02600144
+ dsub = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ voff = -0.1274889
+ ldif = 9e-8
+ tcjsw = 0.0004130718
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ eta0 = 5e-5
+ pvoff = 0.0
+ capmod = 3
+ pvag = 0.0
+ etab = -5e-5
+ vsat = 149999.98
+ wint = 5e-9
+ vth0 = -0.4634952
+ cdscb = 0.0
+ rdsw = 530.0
+ cdscd = 0.0
+ pnfactor = 0
+ peta0 = 1.8966694548261387e-25
+ wkt1 = 8.228274e-9
+ wkt2 = 1.4868883e-9
+ lint = 1.4999999e-8
+ wnfactor = 0.0
+ wmax = 1e-5
+ wketa = 6.301227e-9
+ wmin = 1.2e-6
+ pvth0 = -1.18629e-15
+ mobmod = 1
+ drout = 0.0
+ tpbsw = 0.001572025
+ lmax = 2.0001e-5
+ lmin = 1e-5
+ cjswg = 4.43205e-10
+ a0 = 1.0509492
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ at = 10000.0
+ mjswg = 0.3683619
+ cf = 0
+ cj = 0.00117705
+ lnfactor = -3.9543e-9
+ ef = 1.064
+ k1 = 0.5362856
+ k2 = 0.04116319
+ k3 = 0.0
+ em = 30000000.0
+ js = 2.5e-7
+ ll = 0.0
+ mj = 0.4476
+ lw = 0.0
+ u0 = 0.0109348308
+ pb = 0.895226
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ wvoff = -1.0305298e-9
+ ua = 8.057326e-10
+ ub = 7.508071e-19
+ uc = -7.859605e-11
+ wub1 = 6.909715e-26
+ wuc1 = 3.0354498e-17
+ wl = 0.0
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ hdif = 2e-7
+ weta0 = 0
+ ags = 0.02
+ wute = 1.0600407e-7
+ mjsw = 0.3683619
+ wvsat = 0.0
+ wvth0 = 1.1684168e-8
+ cit = -0.0001
+ dlc = 2e-9
+ nfactor = 1.0
+ k3b = 0.0
+ tcjswg = 0.0004130718
+ dwb = 0.0
+ dwg = 0.0
+ cdsc = 0.0
+ cgdo = 3.28e-10
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0010000004
+ cgso = 3.28e-10
+ pdiblcb = 0.01
+ jsw = 1.2e-12
+ kt1 = -0.231953
+ kt2 = -0.024488758
+ lk2 = 1.18629e-9
+ llc = -0.039
+ lln = -1
+ cjsw = 2.60505e-10
+ lu0 = -7.9086e-11
+ xpart = 1
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ binunit = 2
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ nlx = 0.0
+ pbswg = 0.895226
+ pu0 = 0.0
+ prt = 0
+ tnom = 25.0
+ lvoff = -1.5817200000000002e-9
+ rsh = 7.2
+ beta0 = 22.67827
+ toxm = 4.08e-9
+ tcj = 0.0009739001
+ ua1 = 1.224e-9
+ ub1 = -1.3998005e-18
+ uc1 = -7.633158e-12
+ leta0 = 1.8966694548261387e-18
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ pbsw = 0.895226
+ pclm = 0.6000001
+ tpb = 0.001572025
+ tox = 4.08e-9
+ )

.model pch_fs_6 pmos (
+ level = 49
+ lub1 = 5.442727e-26
+ luc1 = 1.8276951e-17
+ wute = 1.0644106e-7
+ mjsw = 0.3683619
+ tcjsw = 0.0004130718
+ capmod = 3
+ lute = 9.664497e-8
+ pvoff = -4.403278e-15
+ nfactor = 1.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 1.8966694548261387e-25
+ mobmod = 1
+ cgdo = 3.28e-10
+ wketa = 7.084359e-9
+ pvth0 = -6.522762e-15
+ cgso = 3.28e-10
+ drout = 0.0
+ tpbsw = 0.001572025
+ ags = 0.02
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0004772728
+ pdiblcb = 0.01
+ lpscbe1 = 195.04262
+ cjswg = 4.43205e-10
+ cit = -0.0001
+ cjsw = 2.60505e-10
+ mjswg = 0.3683619
+ dlc = 2e-9
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ k3b = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ wvoff = -5.879894e-10
+ binunit = 2
+ tnom = 25.0
+ weta0 = 0
+ wvsat = 0.0
+ toxm = 4.08e-9
+ lpclm = 2.6005682e-7
+ wvth0 = 1.2220496e-8
+ la0 = 6.878132e-8
+ pbsw = 0.895226
+ tcjswg = 0.0004130718
+ pclm = 0.5738637
+ jsw = 1.2e-12
+ kt1 = -0.2303147
+ lk1 = 1.8184398e-8
+ kt2 = -0.024155809
+ lk2 = -4.094344999999999e-9
+ llc = -0.039
+ lln = -1
+ lu0 = -1.3846097e-9
+ lua = -3.935608e-16
+ lub = 4.219459e-25
+ luc = 1.8883157e-17
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ pnfactor = 0
+ pa0 = 6.693222e-14
+ nlx = 0.0
+ wnfactor = 0.0
+ pk1 = 5.986243e-15
+ pk2 = -2.063307e-15
+ pu0 = 1.1543239e-16
+ prt = 0
+ pua = 3.1465633e-23
+ pub = 2.8088595e-31
+ puc = 9.8941e-24
+ version = 3.24
+ lketa = -1.2662711e-9
+ rsh = 7.2
+ pkt1 = 9.666697e-15
+ tcj = 0.0009739001
+ pkt2 = 2.4000725e-15
+ ua1 = 1.224e-9
+ keta = 0.026128704
+ ub1 = -1.4052706e-18
+ uc1 = -9.470036e-12
+ xpart = 1
+ tpb = 0.001572025
+ lnfactor = -3.9543e-9
+ tox = 4.08e-9
+ dsub = 0.0
+ wa0 = -5.459876e-8
+ ute = -0.8492097
+ wk1 = 1.185507e-8
+ wk2 = -5.732776e-9
+ pbswg = 0.895226
+ wln = 1.0
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ wu0 = -1.2808475e-9
+ wua = 1.7227619e-16
+ wub = -6.81325e-25
+ wuc = -8.049533e-17
+ wwl = 0.0
+ wwn = 1.0
+ a0 = 1.0440365
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ lvoff = -3.0500824000000002e-9
+ xti = 3
+ at = 10000.0
+ cf = 0
+ lpdiblc2 = 5.201137e-9
+ cj = 0.00117705
+ voff = -0.1273414
+ ef = 1.064
+ k1 = 0.534458
+ k2 = 0.04169391
+ k3 = 0.0
+ em = 30000000.0
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ ldif = 9e-8
+ beta0 = 22.67827
+ js = 2.5e-7
+ ll = 0.0
+ mj = 0.4476
+ lw = 0.0
+ u0 = 0.0110660398
+ pb = 0.895226
+ kt1l = 0.0
+ w0 = 0.0
+ prwb = 0.0
+ rd = 0
+ pub1 = -6.397619e-32
+ prwg = 0.0
+ leta0 = 1.8966694548261387e-18
+ puc1 = 2.6178952e-23
+ rs = 0
+ ua = 8.452865e-10
+ ub = 7.084005e-19
+ uc = -8.049386e-11
+ pscbe1 = 180397700.0
+ pscbe2 = 5e-7
+ wl = 0.0
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ eta0 = 5e-5
+ lvsat = -0.013002842
+ pvag = 0.0
+ etab = -5e-5
+ vsat = 151306.8
+ lvth0 = -2.8234169e-8
+ wint = 5e-9
+ pute = -4.348101e-15
+ vth0 = -0.4610551
+ nqsmod = 0
+ rdsw = 530.0
+ tpbswg = 0.001572025
+ delta = 0.01
+ wkt1 = 7.256747e-9
+ wkt2 = 1.245675e-9
+ noimod = 2
+ lint = 1.4999999e-8
+ wmax = 1e-5
+ wmin = 1.2e-6
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ lkt1 = -1.6300865e-8
+ lkt2 = -3.312836e-9
+ lmax = 1e-5
+ lmin = 1.2e-6
+ pketa = -7.792167e-15
+ wub1 = 7.552692e-26
+ wuc1 = 2.7723443e-17
+ hdif = 2e-7
+ )

.model pch_fs_7 pmos (
+ level = 49
+ mjswg = 0.3683619
+ jsw = 1.2e-12
+ kt1 = -0.2459144
+ lk1 = 8.371453e-9
+ kt2 = -0.027846618
+ lk2 = -2.029564e-9
+ dsub = 0.0
+ llc = -0.039
+ lln = -1
+ lu0 = -4.248086e-10
+ wvoff = -7.866491e-9
+ lua = 3.0792715e-17
+ lub = -1.9665828e-25
+ luc = -3.700045e-17
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ wcit = -1.788104e-11
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ pa0 = -1.2519753e-13
+ nlx = 0.0
+ weta0 = 0
+ pk1 = 4.753178e-14
+ pk2 = -1.4849934e-14
+ lcit = 2.2196864e-10
+ voff = -0.1274479
+ pu0 = -6.201592e-16
+ wvsat = 0.0
+ ldif = 9e-8
+ tcjswg = 0.0004130718
+ prt = 0
+ pua = -3.495584e-22
+ pub = 3.345938e-31
+ puc = 4.854297e-23
+ lpclm = 1.4785702e-7
+ wvth0 = 8.94442e-9
+ kt1l = 0.0
+ prwb = 0.0
+ pub1 = -1.382964e-31
+ prwg = 0.0
+ puc1 = -5.043768e-23
+ eta0 = 1.7857139e-5
+ rsh = 7.2
+ tcj = 0.0009739001
+ ua1 = 1.224e-9
+ pvag = 0.0
+ ub1 = -1.3967723e-18
+ etab = -1.7857139e-5
+ uc1 = -2.3838735e-11
+ vsat = 146428.53
+ wint = 5e-9
+ pute = 2.0900147e-14
+ tpb = 0.001572025
+ tox = 4.08e-9
+ vth0 = -0.4764877
+ wa0 = 1.1247056e-7
+ rdsw = 530.0
+ ute = -0.7951261
+ wkt1 = 1.6218328e-8
+ wkt2 = 2.9642964e-9
+ wk1 = -2.4271484e-8
+ wk2 = 5.386031e-9
+ lint = 1.4999999e-8
+ wmax = 1e-5
+ wln = 1.0
+ wu0 = -6.412026e-10
+ wmin = 1.2e-6
+ wua = 5.036014e-16
+ wub = -7.280275e-25
+ wuc = -1.1410304e-16
+ lkt1 = 1.6387112e-9
+ lkt2 = 9.315946e-10
+ wwl = 0.0
+ wwn = 1.0
+ xti = 3
+ lmax = 1.2e-6
+ lketa = -8.380984e-9
+ lmin = 5e-7
+ xpart = 1
+ wub1 = 1.4015321e-25
+ pbswg = 0.895226
+ wuc1 = 9.434661e-17
+ hdif = 2e-7
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ lvoff = -2.9275995000000004e-9
+ lub1 = 4.46543e-26
+ luc1 = 3.480094e-17
+ wute = 8.448607e-8
+ mjsw = 0.3683619
+ pscbe1 = 349999900.0
+ pscbe2 = 5e-7
+ beta0 = 22.67827
+ leta0 = 3.6964291896669454e-11
+ lute = 3.444881e-8
+ letab = -3.696429e-11
+ lvsat = -0.007392833
+ lvth0 = -1.0486687e-8
+ nqsmod = 0
+ tpbswg = 0.001572025
+ noimod = 2
+ cdsc = 0.0
+ pnfactor = 0
+ delta = 0.01
+ wnfactor = 0.0
+ cgdo = 3.28e-10
+ nfactor = 1.0
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ cgso = 3.28e-10
+ cjsw = 2.60505e-10
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0017857144
+ lnfactor = -3.9543e-9
+ pdiblcb = 0.01
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ pketa = 2.2253538e-15
+ tnom = 25.0
+ binunit = 2
+ capmod = 3
+ lpdiblc2 = 3.696428e-9
+ tcjsw = 0.0004130718
+ toxm = 4.08e-9
+ ags = 0.02
+ pcit = 2.0563189e-17
+ pbsw = 0.895226
+ pclm = 0.6714287
+ pvoff = 3.966999e-15
+ cit = -0.0002930162
+ a0 = 0.9932752
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ at = 10000.0
+ mobmod = 1
+ cf = 0
+ dlc = 2e-9
+ cj = 0.00117705
+ ef = 1.064
+ k1 = 0.542991
+ k2 = 0.03989844
+ k3 = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ em = 30000000.0
+ peta0 = 1.8966694548261387e-25
+ k3b = 0.0
+ js = 2.5e-7
+ ll = 0.0
+ mj = 0.4476
+ lw = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ u0 = 0.0102314288
+ pb = 0.895226
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ua = 4.762835e-10
+ ub = 1.2463172e-18
+ uc = -3.189942e-11
+ wl = 0.0
+ wr = 1.0
+ xj = 1.7000001e-7
+ wketa = -1.6265284e-9
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ pvth0 = -2.7552727999999998e-15
+ drout = 0.0
+ tpbsw = 0.001572025
+ pkt1 = -6.391237e-16
+ pkt2 = 4.236579e-16
+ keta = 0.03231541
+ cjswg = 4.43205e-10
+ version = 3.24
+ la0 = 1.2715688e-7
+ )

.model pch_fs_8 pmos (
+ level = 49
+ cgso = 3.28e-10
+ nfactor = 1.0
+ a0 = 1.2640158
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ lketa = -5.872592e-10
+ at = 10000.0
+ cf = 0
+ cj = 0.00117705
+ ef = 1.064
+ k1 = 0.5203763
+ k2 = 0.04747528
+ k3 = 0.0
+ em = 30000000.0
+ pcdscd = -7.408954e-18
+ js = 2.5e-7
+ ll = 0.0
+ mj = 0.4476
+ lw = 0.0
+ u0 = 0.0097404008
+ pb = 0.895226
+ xpart = 1
+ w0 = 0.0
+ rd = 0
+ cjsw = 2.60505e-10
+ rs = 0
+ ua = 9.357863e-10
+ ub = 5.091257e-19
+ uc = -1.5731644e-10
+ wl = 0.0
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.007987866
+ pbswg = 0.895226
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ pdiblcb = 0.01
+ pscbe1 = 350000000.0
+ pscbe2 = 5e-7
+ lvoff = -1.4181850500000001e-9
+ tnom = 25.0
+ pags = -6.875222e-16
+ beta0 = 22.67827
+ toxm = 4.08e-9
+ binunit = 2
+ leta0 = 2.559375218966695e-10
+ letab = -5.545772e-10
+ nqsmod = 0
+ pcit = -7.907631e-17
+ pbsw = 0.895226
+ pclm = 0.9107697
+ tpbswg = 0.001572025
+ lvsat = -0.0003656271
+ noimod = 2
+ lvth0 = -1.2082326e-8
+ ppclm = 2.4445072e-15
+ delta = 0.01
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ lcdscd = 3.730414e-11
+ pkt1 = -1.8229216e-15
+ pkt2 = -1.2254391e-15
+ keta = 0.014996022
+ ags = 0.019847063
+ wags = 1.5278273e-9
+ dsub = 0.0
+ version = 3.24
+ cit = -6.09184e-5
+ pketa = -2.4325694e-15
+ dlc = 2e-9
+ lags = 6.882101e-11
+ wcit = 2.0354016e-10
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ k3b = 0.0
+ capmod = 3
+ dwb = 0.0
+ dwg = 0.0
+ wpclm = -5.432238e-9
+ lcit = 1.1752459e-10
+ voff = -0.1308021
+ tcjsw = 0.0004130718
+ ldif = 9e-8
+ kt1l = 0.0
+ prwb = 0.0
+ pub1 = 2.7781507e-32
+ prwg = 0.0
+ puc1 = 8.113434e-24
+ pvoff = -1.9905158e-15
+ eta0 = -0.0004687502
+ mobmod = 1
+ pvag = 0.0
+ etab = 0.0011323938
+ la0 = 5.323636e-9
+ vsat = 130812.52
+ wint = 5e-9
+ pute = 9.798417e-15
+ jsw = 1.2e-12
+ kt1 = -0.2367561
+ lk1 = 1.854804e-8
+ kt2 = -0.025532207
+ lk2 = -5.439136e-9
+ vth0 = -0.4729418
+ cdscb = 0.0
+ cdscd = -8.289813e-5
+ pnfactor = 0
+ peta0 = 1.8966694548261387e-25
+ llc = -0.039
+ rdsw = 530.0
+ lln = -1
+ lu0 = -2.0384533e-10
+ petab = 2.4660761e-16
+ wnfactor = 0.0
+ wkt1 = 1.8848993e-8
+ wkt2 = 6.628956e-9
+ lua = -1.759835e-16
+ lub = 1.3507784e-25
+ luc = 1.9437196e-17
+ lint = 1.4999999e-8
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ wmax = 1e-5
+ wketa = 8.724413e-9
+ pvth0 = -2.3104256e-15
+ pa0 = 1.0862038e-13
+ nlx = 0.0
+ wmin = 1.2e-6
+ drout = 0.0
+ lkt1 = -2.4825255e-9
+ lkt2 = -1.0989117e-10
+ tpbsw = 0.001572025
+ pk1 = -1.7383759e-14
+ pk2 = 7.484627e-15
+ lmax = 5e-7
+ pu0 = 2.5785697e-16
+ lmin = 1.8e-7
+ ppdiblc2 = 8.594017e-17
+ prt = 0
+ pua = 1.5976873e-22
+ pub = -1.3085017e-31
+ puc = -9.356197e-24
+ cjswg = 4.43205e-10
+ wpdiblc2 = -1.9097854e-10
+ mjswg = 0.3683619
+ lnfactor = -3.9543e-9
+ rsh = 7.2
+ tcj = 0.0009739001
+ ua1 = 1.224e-9
+ ub1 = -1.3554493e-18
+ uc1 = 7.051652e-11
+ wvoff = 5.372431e-9
+ tpb = 0.001572025
+ tox = 4.08e-9
+ wub1 = -2.2890885e-25
+ wuc1 = -3.576699e-17
+ wa0 = -4.071248e-7
+ hdif = 2e-7
+ ute = -0.7199521
+ wk1 = 1.1998529e-7
+ wk2 = -4.424634e-8
+ weta0 = 0
+ tcjswg = 0.0004130718
+ lub1 = 2.6058948e-26
+ luc1 = -7.658915e-18
+ wln = 1.0
+ wetab = -5.480169e-10
+ lpdiblc2 = 9.0546e-10
+ wu0 = -2.5923497e-9
+ wute = 1.0915658e-7
+ mjsw = 0.3683619
+ wvsat = 0.0
+ wua = -6.282368e-16
+ wub = 3.0629255e-25
+ wuc = 1.4561782e-17
+ wwl = 0.0
+ wwn = 1.0
+ lpclm = 4.015361e-8
+ wvth0 = 7.955874e-9
+ xti = 3
+ lute = 6.205235e-10
+ cdsc = 0.0
+ wcdscd = 1.6464351e-11
+ cgdo = 3.28e-10
+ )

.model pch_fs_9 pmos (
+ level = 49
+ pvag = 0.0
+ etab = -5e-5
+ lvth0 = -3.9543e-9
+ ags = 0.02
+ vsat = 149999.98
+ wint = 5e-9
+ vth0 = -0.4523646
+ delta = 0.01
+ rdsw = 530.0
+ cit = -0.0001
+ wkt1 = 6.74333e-9
+ wkt2 = 1.2948118e-10
+ lint = 1.4999999e-8
+ dlc = 2e-9
+ wmax = 1.2e-6
+ dvt0w = 0.0
+ k3b = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ wmin = 5e-7
+ dwb = 0.0
+ dwg = 0.0
+ lmax = 2.0001e-5
+ lmin = 1e-5
+ capmod = 3
+ a0 = 0.9810578
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ jsw = 1.2e-12
+ kt1 = -0.2307052
+ kt2 = -0.02334808
+ lk2 = 1.18629e-9
+ wub1 = 3.495163e-26
+ wuc1 = 1.9335648e-17
+ at = 10000.0
+ cf = 0
+ cj = 0.00117705
+ ef = 1.064
+ k1 = 0.5449055
+ k2 = 0.0393854
+ k3 = 0.0
+ em = 30000000.0
+ llc = -0.039
+ lln = -1
+ lu0 = -7.9086e-11
+ hdif = 2e-7
+ js = 2.5e-7
+ ll = 0.0
+ mj = 0.4476
+ lw = 0.0
+ u0 = 0.0100768048
+ nch = 3.9e+17
+ pb = 0.895226
+ w0 = 0.0
+ rd = 0
+ lwl = 0.0
+ lwn = 1.0
+ rs = 0
+ ua = 1.0698959e-9
+ ub = 3.0837888e-19
+ uc = -1.1659398e-10
+ wl = 0.0
+ wute = -2.7886795e-9
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ mjsw = 0.3683619
+ nlx = 0.0
+ tcjsw = 0.0004130718
+ mobmod = 1
+ pu0 = 0.0
+ pvoff = 0.0
+ prt = 0
+ rsh = 7.2
+ cdscb = 0.0
+ cdscd = 0.0
+ tcj = 0.0009739001
+ peta0 = 1.8966694548261387e-25
+ cdsc = 0.0
+ ua1 = 1.224e-9
+ ub1 = -1.3711068e-18
+ uc1 = 1.6263793e-12
+ tpb = 0.001572025
+ tox = 4.08e-9
+ cgdo = 3.28e-10
+ wketa = -1.0458587e-9
+ wa0 = 3.529885e-8
+ pvth0 = -1.18629e-15
+ drout = 0.0
+ ute = -0.7480742
+ wk1 = 2.1990281e-9
+ cgso = 3.28e-10
+ wk2 = -3.824582e-9
+ tpbsw = 0.001572025
+ wln = 1.0
+ wu0 = -2.481951e-10
+ wua = -1.3891575e-16
+ wub = -1.2660565e-25
+ wuc = -3.428342e-17
+ wwl = 0.0
+ wwn = 1.0
+ cjswg = 4.43205e-10
+ nfactor = 1.0
+ xti = 3
+ cjsw = 2.60505e-10
+ mjswg = 0.3683619
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ wvoff = -4.105241e-10
+ tcjswg = 0.0004130718
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0009999998
+ weta0 = 0
+ tnom = 25.0
+ pdiblcb = 0.01
+ wvsat = 0.0
+ wvth0 = -1.5613511000000001e-9
+ toxm = 4.08e-9
+ pbsw = 0.895226
+ pclm = 0.6
+ binunit = 2
+ pnfactor = 0
+ wnfactor = 0.0
+ keta = 0.03217546
+ xpart = 1
+ lnfactor = -3.9543e-9
+ alpha0 = 0.0
+ dsub = 0.0
+ alpha1 = 6.8730453846
+ pbswg = 0.895226
+ pscbe1 = 199999970.0
+ pscbe2 = 5e-7
+ dvt0 = 0.0
+ version = 3.24
+ dvt1 = 0.0
+ dvt2 = 0.0
+ lvoff = -1.5817200000000002e-9
+ voff = -0.12801
+ beta0 = 22.67827
+ nqsmod = 0
+ ldif = 9e-8
+ tpbswg = 0.001572025
+ noimod = 2
+ leta0 = 1.8966694548261387e-18
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ eta0 = 5e-5
+ )

.model pch_fs_10 pmos (
+ level = 49
+ dsub = 0.0
+ wk1 = 1.7598129e-9
+ wk2 = -3.600003e-9
+ wln = 1.0
+ wu0 = -2.1789574e-10
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ wua = -1.6455617e-16
+ wub = -7.150721e-26
+ wuc = -2.8652769e-17
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ wwl = 0.0
+ wwn = 1.0
+ xti = 3
+ pscbe1 = 180397680.0
+ pscbe2 = 5e-7
+ voff = -0.1269095
+ ldif = 9e-8
+ nfactor = 1.0
+ kt1l = 0.0
+ prwb = 0.0
+ pub1 = -8.629597e-32
+ prwg = 0.0
+ puc1 = 1.5034668e-23
+ nqsmod = 0
+ tpbswg = 0.001572025
+ lketa = -6.417587e-9
+ eta0 = 5e-5
+ noimod = 2
+ pvag = 0.0
+ etab = -5e-5
+ vsat = 151306.8
+ wint = 5e-9
+ pute = 3.909688e-14
+ xpart = 1
+ vth0 = -0.4482969
+ rdsw = 530.0
+ wkt1 = 6.495125e-9
+ wkt2 = 2.3726165e-10
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0004772722
+ lint = 1.4999999e-8
+ pdiblcb = 0.01
+ lpscbe1 = 195.04263
+ wmax = 1.2e-6
+ pbswg = 0.895226
+ wmin = 5e-7
+ lkt1 = -1.0252924e-8
+ lkt2 = -3.947785e-10
+ lmax = 1e-5
+ lvoff = -1.2530685e-8
+ lmin = 1.2e-6
+ beta0 = 22.67827
+ binunit = 2
+ leta0 = 1.8966694548261387e-18
+ lvsat = -0.013002842
+ lvth0 = -4.442723e-8
+ wub1 = 4.362458e-26
+ wuc1 = 1.7824627e-17
+ capmod = 3
+ hdif = 2e-7
+ delta = 0.01
+ lub1 = 7.318341e-26
+ luc1 = 2.7641896e-17
+ pnfactor = 0
+ wute = -6.718015e-9
+ mjsw = 0.3683619
+ wnfactor = 0.0
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ lute = 6.013659e-8
+ mobmod = 1
+ cdsc = 0.0
+ version = 3.24
+ lnfactor = -3.9543e-9
+ pketa = -1.6621007e-15
+ cgdo = 3.28e-10
+ ags = 0.02
+ cgso = 3.28e-10
+ cit = -0.0001
+ tcjsw = 0.0004130718
+ dlc = 2e-9
+ lpdiblc2 = 5.201137e-9
+ cjsw = 2.60505e-10
+ k3b = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ pvoff = 6.87864e-15
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 1.8966694548261387e-25
+ tcjswg = 0.0004130718
+ tnom = 25.0
+ wketa = -8.788133e-10
+ pvth0 = 1.274698e-14
+ la0 = 1.2176828e-7
+ drout = 0.0
+ toxm = 4.08e-9
+ jsw = 1.2e-12
+ kt1 = -0.2296747
+ lk1 = 1.9542425e-8
+ kt2 = -0.023308404
+ lk2 = -3.950429e-9
+ tpbsw = 0.001572025
+ pbsw = 0.895226
+ llc = -0.039
+ pclm = 0.5738636
+ lln = -1
+ lu0 = -1.0342642e-9
+ lua = -5.815077e-16
+ lub = 1.1186816e-24
+ luc = 7.427734e-17
+ nch = 3.9e+17
+ a0 = 0.9688198
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ lwl = 0.0
+ lwn = 1.0
+ cjswg = 4.43205e-10
+ at = 10000.0
+ cf = 0
+ cj = 0.00117705
+ pa0 = 3.87773e-15
+ nlx = 0.0
+ ef = 1.064
+ k1 = 0.5429414
+ k2 = 0.039901660000000005
+ k3 = 0.0
+ em = 30000000.0
+ mjswg = 0.3683619
+ js = 2.5e-7
+ ll = 0.0
+ mj = 0.4476
+ lw = 0.0
+ pk1 = 4.370194e-15
+ pk2 = -2.2345663e-15
+ u0 = 0.0101728028
+ pb = 0.895226
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ua = 1.1283389e-9
+ ub = 1.9594849e-19
+ uc = -1.2405904e-10
+ wvoff = -1.1018445e-9
+ wl = 0.0
+ pu0 = -3.0147877e-16
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ prt = 0
+ pua = 2.5512236e-22
+ pub = -5.482294e-31
+ puc = -5.602498e-23
+ weta0 = 0
+ rsh = 7.2
+ tcj = 0.0009739001
+ ua1 = 1.224e-9
+ ub1 = -1.3784619e-18
+ uc1 = -1.1517035e-12
+ wvsat = 0.0
+ pkt1 = 2.469645e-15
+ pkt2 = -1.0724159e-15
+ keta = 0.03282044
+ tpb = 0.001572025
+ tox = 4.08e-9
+ lpclm = 2.6005682e-7
+ wvth0 = -2.9616815e-9
+ wa0 = 3.490912e-8
+ ute = -0.754118
+ )

.model pch_fs_11 pmos (
+ level = 49
+ cgso = 3.28e-10
+ a0 = 1.1936638
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ lvoff = 3.655491e-9
+ at = 10000.0
+ cf = 0
+ cj = 0.00117705
+ ef = 1.064
+ k1 = 0.4715038
+ k2 = 0.06532277
+ k3 = 0.0
+ em = 30000000.0
+ js = 2.5e-7
+ ll = 0.0
+ mj = 0.4476
+ lw = 0.0
+ beta0 = 22.67827
+ u0 = 0.0106717438
+ pb = 0.895226
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ua = 1.036115e-9
+ ub = 1.0523674e-18
+ uc = -7.205117e-11
+ cjsw = 2.60505e-10
+ leta0 = 3.696426189666945e-11
+ wl = 0.0
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ letab = -3.696426e-11
+ lvsat = -0.007392855
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ capmod = 3
+ lvth0 = -7.517002e-9
+ delta = 0.01
+ tnom = 25.0
+ ags = 0.02
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ toxm = 4.08e-9
+ mobmod = 1
+ pcit = -1.0851648e-17
+ pbsw = 0.895226
+ pclm = 0.6714286
+ cit = -0.00031597191
+ dlc = 2e-9
+ k3b = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ pketa = 4.024799e-15
+ la0 = -1.3680231e-7
+ pkt1 = -6.051915e-15
+ pkt2 = -1.4802061e-15
+ tcjsw = 0.0004130718
+ keta = 0.03584265
+ jsw = 1.2e-12
+ kt1 = -0.2439705
+ lk1 = 1.0169572e-7
+ kt2 = -0.025852976
+ lk2 = -3.3184709999999996e-8
+ llc = -0.039
+ lln = -1
+ lu0 = -1.6080454999999999e-9
+ dsub = 0.0
+ pvoff = -3.866879e-15
+ lua = -4.754501e-16
+ lub = 1.337998e-25
+ luc = 1.4468274e-17
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ pa0 = 1.8891395e-13
+ nlx = 0.0
+ tcjswg = 0.0004130718
+ wcit = 9.436221e-12
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ pk1 = -6.35241e-14
+ pk2 = 2.2224691e-14
+ peta0 = 1.8966694548261387e-25
+ pu0 = 7.878928e-16
+ pnfactor = 0
+ prt = 0
+ lcit = 2.4836766e-10
+ pua = 2.5287059e-22
+ pub = -5.865131e-32
+ puc = -1.2704817e-23
+ wketa = -5.823942e-9
+ voff = -0.1409845
+ pvth0 = -6.289198e-15
+ wnfactor = 0.0
+ ldif = 9e-8
+ drout = 0.0
+ kt1l = 0.0
+ tpbsw = 0.001572025
+ prwb = 0.0
+ pub1 = 4.97241e-32
+ prwg = 0.0
+ rsh = 7.2
+ puc1 = 1.7282469e-23
+ tcj = 0.0009739001
+ ua1 = 1.224e-9
+ ub1 = -1.2162624e-18
+ uc1 = 4.210797e-11
+ eta0 = 1.7857154e-5
+ nfactor = 1.0
+ pvag = 0.0
+ etab = -1.7857154e-5
+ tpb = 0.001572025
+ tox = 4.08e-9
+ cjswg = 4.43205e-10
+ vsat = 146428.56
+ wa0 = -1.2599192e-7
+ wint = 5e-9
+ pute = -5.928695e-14
+ mjswg = 0.3683619
+ vth0 = -0.4803928
+ ute = -0.7903757
+ wk1 = 6.079834e-8
+ wk2 = -2.4868919e-8
+ rdsw = 530.0
+ wln = 1.0
+ wkt1 = 1.3905176e-8
+ wkt2 = 5.918618e-10
+ lnfactor = -3.9543e-9
+ wu0 = -1.1651754e-9
+ lint = 1.4999999e-8
+ wvoff = 8.242083e-9
+ wua = -1.625981e-16
+ wmax = 1.2e-6
+ wub = -4.972273e-25
+ wuc = -6.632247e-17
+ wwl = 0.0
+ wwn = 1.0
+ wmin = 5e-7
+ xti = 3
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0017857137
+ lkt1 = 6.187276e-9
+ lkt2 = 2.5314804e-9
+ pdiblcb = 0.01
+ weta0 = 0
+ lmax = 1.2e-6
+ lmin = 5e-7
+ wvsat = 0.0
+ lpclm = 1.4785714e-7
+ wvth0 = 1.3591517e-8
+ lpdiblc2 = 3.696429e-9
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ binunit = 2
+ pscbe1 = 349999900.0
+ pscbe2 = 5e-7
+ wub1 = -7.465372e-26
+ wuc1 = 1.5870021e-17
+ hdif = 2e-7
+ lub1 = -1.133461e-25
+ luc1 = -2.2106738e-17
+ wute = 7.883313e-8
+ mjsw = 0.3683619
+ nqsmod = 0
+ tpbswg = 0.001572025
+ noimod = 2
+ lute = 1.0183292e-7
+ lketa = -9.893122e-9
+ xpart = 1
+ cdsc = 0.0
+ cgdo = 3.28e-10
+ pbswg = 0.895226
+ version = 3.24
+ )

.model pch_fs_12 pmos (
+ level = 49
+ wint = 5e-9
+ llc = -0.039
+ pute = 1.3160581e-15
+ lln = -1
+ lu0 = 1.3290007e-10
+ vth0 = -0.47008160000000004
+ nfactor = 1.0
+ lua = 2.3815556e-17
+ lub = -3.425063e-26
+ luc = 8.803578e-18
+ nch = 3.9e+17
+ rdsw = 530.0
+ lwl = 0.0
+ lwn = 1.0
+ pketa = -9.609158e-16
+ wkt1 = 2.7434011e-10
+ wkt2 = -6.113567e-9
+ lint = 1.4999999e-8
+ pa0 = -8.476619e-14
+ nlx = 0.0
+ wmax = 1.2e-6
+ pk1 = 1.5213101e-14
+ pk2 = -6.235986e-15
+ wmin = 5e-7
+ lkt1 = -4.083267e-9
+ lkt2 = -2.4314675e-9
+ wpclm = 5.671285e-8
+ pu0 = -1.4287007e-16
+ lmax = 5e-7
+ prt = 0
+ pua = -7.799214e-23
+ pub = 7.065072e-32
+ puc = 3.297807e-24
+ lmin = 1.8e-7
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.009150297
+ tcjsw = 0.0004130718
+ pdiblcb = 0.01
+ rsh = 7.2
+ tcj = 0.0009739001
+ ua1 = 1.224e-9
+ ub1 = -1.6175756e-18
+ uc1 = -2.2818641e-11
+ pvoff = -1.4343533e-15
+ tcjswg = 0.0004130718
+ tpb = 0.001572025
+ tox = 4.08e-9
+ a0 = 0.5166956
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ wa0 = 4.821862e-7
+ at = 10000.0
+ cf = 0
+ cj = 0.00117705
+ wub1 = 8.30214e-26
+ ute = -0.5812994
+ wuc1 = 7.530186e-17
+ ef = 1.064
+ k1 = 0.7171482
+ k2 = -0.021956119
+ k3 = 0.0
+ em = 30000000.0
+ wk1 = -1.1417325e-7
+ wk2 = 3.837703e-8
+ binunit = 2
+ cdscb = 0.0
+ cdscd = -5.200001e-5
+ peta0 = 1.8966694548261387e-25
+ js = 2.5e-7
+ ll = 0.0
+ mj = 0.4476
+ hdif = 2e-7
+ lw = 0.0
+ u0 = 0.0068029748
+ wln = 1.0
+ pb = 0.895226
+ w0 = 0.0
+ wu0 = 9.031869e-10
+ rd = 0
+ rs = 0
+ ua = -7.336427e-11
+ ub = 1.4258127e-18
+ uc = -5.946296e-11
+ lub1 = 6.724484e-26
+ wua = 5.726523e-16
+ wub = -7.845651e-25
+ wuc = -1.0188386e-16
+ wl = 0.0
+ luc1 = 7.110234e-18
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ wwl = 0.0
+ wwn = 1.0
+ wute = -5.584022e-8
+ wketa = 5.255423e-9
+ mjsw = 0.3683619
+ pvth0 = -2.2215402e-15
+ xti = 3
+ drout = 0.0
+ tpbsw = 0.001572025
+ lute = 7.748556e-9
+ wcdscd = -2.0304376e-11
+ cjswg = 4.43205e-10
+ mjswg = 0.3683619
+ cdsc = 0.0
+ wvoff = 2.8364715e-9
+ cgdo = 3.28e-10
+ pcdscd = 9.13697e-18
+ cgso = 3.28e-10
+ weta0 = 0
+ version = 3.24
+ wvsat = 0.0
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ lpclm = 6.365384e-8
+ wvth0 = 4.552275e-9
+ cjsw = 2.60505e-10
+ pscbe1 = 350000000.0
+ pscbe2 = 5e-7
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ nqsmod = 0
+ tpbswg = 0.001572025
+ tnom = 25.0
+ pnfactor = 0
+ noimod = 2
+ pags = -5.667374e-15
+ wnfactor = 0.0
+ toxm = 4.08e-9
+ pcit = 2.6834248e-18
+ pbsw = 0.895226
+ lketa = -1.8239428e-9
+ pclm = 0.858547
+ xpart = 1
+ ppdiblc2 = 7.08422e-16
+ wpdiblc2 = -1.5742713e-9
+ lnfactor = -3.9543e-9
+ pbswg = 0.895226
+ lcdscd = 2.3400004e-11
+ lvoff = -1.8855486300000003e-9
+ ags = 0.010547621
+ beta0 = 22.67827
+ pkt1 = 8.196091e-17
+ pkt2 = 1.5372367e-15
+ keta = 0.01791114
+ lpdiblc2 = 3.823661e-10
+ leta0 = 2.5593747189666946e-10
+ capmod = 3
+ letab = -3.473438e-10
+ cit = 0.00012746976
+ wags = 1.2594167e-8
+ lvsat = -0.0003656142
+ dsub = 0.0
+ dlc = 2e-9
+ lvth0 = -1.2157019e-8
+ k3b = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ lags = 4.253569e-9
+ wcit = -2.0641719e-11
+ ppclm = -2.5520774e-14
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ delta = 0.01
+ mobmod = 1
+ lcit = 4.881893e-11
+ voff = -0.1286711
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ ldif = 9e-8
+ kt1l = 0.0
+ prwb = 0.0
+ pub1 = -2.1229706e-32
+ prwg = 0.0
+ puc1 = -9.461855e-24
+ la0 = 1.6783336e-7
+ eta0 = -0.00046875
+ pvag = 0.0
+ jsw = 1.2e-12
+ etab = 0.0006718753
+ kt1 = -0.2211471
+ lk1 = -8.844278e-9
+ kt2 = -0.014824204
+ lk2 = 6.090789e-9
+ vsat = 130812.46
+ )

.model pch_fs_13 pmos (
+ level = 49
+ wketa = -6.403492e-9
+ pvth0 = -1.18629e-15
+ drout = 0.0
+ toxm = 4.08e-9
+ tpbsw = 0.001572025
+ pbsw = 0.895226
+ pclm = 0.5999999
+ cjswg = 4.43205e-10
+ mjswg = 0.3683619
+ wvoff = -1.320298e-9
+ weta0 = 0
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ wvsat = 0.0
+ keta = 0.04310941
+ pscbe1 = 199999970.0
+ pscbe2 = 5e-7
+ wvth0 = 8.154323e-9
+ dsub = 0.0
+ nqsmod = 0
+ tpbswg = 0.001572025
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ noimod = 2
+ voff = -0.1261533
+ ldif = 9e-8
+ a0 = 0.8704194
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ at = 10000.0
+ cf = 0
+ cj = 0.00117705
+ ef = 1.064
+ k1 = 0.5421249
+ k2 = 0.04121244
+ k3 = 0.0
+ em = 30000000.0
+ ags = 0.02
+ eta0 = 5e-5
+ js = 2.5e-7
+ ll = 0.0
+ mj = 0.4476
+ lw = 0.0
+ pvag = 0.0
+ etab = -5e-5
+ u0 = 0.0096929738
+ pb = 0.895226
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ vsat = 149999.98
+ xpart = 1
+ ua = 1.2584637e-9
+ ub = 4.999999e-20
+ uc = -1.6065008e-10
+ wint = 5e-9
+ wl = 0.0
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ cit = -0.0001
+ vth0 = -0.4721925
+ rdsw = 530.0
+ dlc = 2e-9
+ wkt1 = 3.830554e-9
+ wkt2 = 1.9527771e-9
+ k3b = 0.0
+ lint = 1.4999999e-8
+ pbswg = 0.895226
+ dwb = 0.0
+ wmax = 5e-7
+ dwg = 0.0
+ nfactor = 1.0
+ wmin = 2.2e-7
+ lvoff = -1.5817200000000002e-9
+ lmax = 2.0001e-5
+ lmin = 1e-5
+ capmod = 3
+ beta0 = 22.67827
+ leta0 = 1.8966694548261387e-18
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.001
+ pdiblcb = 0.01
+ jsw = 1.2e-12
+ kt1 = -0.2247607
+ kt2 = -0.027069092
+ lk2 = 1.18629e-9
+ lvth0 = -3.9543e-9
+ llc = -0.039
+ lln = -1
+ lu0 = -7.9086e-11
+ wub1 = 2.1644123e-27
+ wuc1 = -1.2526765e-17
+ nch = 3.9e+17
+ mobmod = 1
+ lwl = 0.0
+ lwn = 1.0
+ delta = 0.01
+ hdif = 2e-7
+ nlx = 0.0
+ pnfactor = 0
+ binunit = 2
+ wute = 6.898109e-9
+ mjsw = 0.3683619
+ wnfactor = 0.0
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ pu0 = 0.0
+ prt = 0
+ rsh = 7.2
+ tcj = 0.0009739001
+ ua1 = 1.224e-9
+ ub1 = -1.3041941e-18
+ uc1 = 6.665171e-11
+ cdsc = 0.0
+ tpb = 0.001572025
+ tox = 4.08e-9
+ wa0 = 8.951166e-8
+ lnfactor = -3.9543e-9
+ cgdo = 3.28e-10
+ ute = -0.7678431
+ wk1 = 3.561511e-9
+ wk2 = -4.719829e-9
+ wln = 1.0
+ cgso = 3.28e-10
+ wu0 = -6.011836e-11
+ wua = -2.3131395e-16
+ wuc = -1.2695932e-17
+ wwl = 0.0
+ wwn = 1.0
+ xti = 3
+ tcjsw = 0.0004130718
+ tcjswg = 0.0004130718
+ version = 3.24
+ cjsw = 2.60505e-10
+ pvoff = 0.0
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 1.8966694548261387e-25
+ tnom = 25.0
+ )

.model pch_fs_14 pmos (
+ level = 49
+ tpbswg = 0.001572025
+ noimod = 2
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0004772729
+ cit = -0.0001
+ wub1 = -3.0198158e-27
+ wuc1 = -1.0513175e-17
+ pdiblcb = 0.01
+ lpscbe1 = 195.04262
+ dlc = 2e-9
+ hdif = 2e-7
+ k3b = 0.0
+ lub1 = -2.0820251e-25
+ dwb = 0.0
+ dwg = 0.0
+ luc1 = 9.921307e-17
+ wute = 1.1298283e-8
+ mjsw = 0.3683619
+ binunit = 2
+ lketa = -4.562476e-8
+ lute = 2.2927659e-7
+ xpart = 1
+ la0 = 5.081137e-7
+ cdsc = 0.0
+ jsw = 1.2e-12
+ kt1 = -0.2237138
+ lk1 = -4.88067e-8
+ kt2 = -0.026908273
+ lk2 = 2.4488488e-8
+ llc = -0.039
+ lln = -1
+ cgdo = 3.28e-10
+ lu0 = -3.7909119e-10
+ pbswg = 0.895226
+ lua = -3.24011e-17
+ lub = -3.941427e-28
+ luc = -6.882293e-17
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ cgso = 3.28e-10
+ pa0 = -1.854315e-13
+ lvoff = -3.9703229000000005e-9
+ nlx = 0.0
+ capmod = 3
+ pk1 = 3.786126e-14
+ pk2 = -1.6169635e-14
+ beta0 = 22.67827
+ pu0 = -6.225135e-16
+ leta0 = 1.8966694548261387e-18
+ prt = 0
+ pua = -1.3939852e-23
+ pub = 1.1764949e-34
+ puc = 1.4094153e-23
+ cjsw = 2.60505e-10
+ lvsat = -0.013002842
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ lvth0 = -8.562635e-9
+ version = 3.24
+ rsh = 7.2
+ tcj = 0.0009739001
+ mobmod = 1
+ ua1 = 1.224e-9
+ ub1 = -1.2832692e-18
+ uc1 = 5.668055e-11
+ tpb = 0.001572025
+ tox = 4.08e-9
+ delta = 0.01
+ wa0 = 1.0814799e-7
+ tnom = 25.0
+ ute = -0.790886
+ wk1 = -2.4364055e-10
+ wk2 = -3.0947396e-9
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ wln = 1.0
+ wu0 = 2.4458129999999986e-12
+ toxm = 4.08e-9
+ wua = -2.2991296e-16
+ wub = -1.1822094e-29
+ wuc = -1.4112429e-17
+ wwl = 0.0
+ wwn = 1.0
+ pbsw = 0.895226
+ xti = 3
+ pclm = 0.5738635
+ pketa = 1.7549415e-14
+ a0 = 0.8193527
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ at = 10000.0
+ cf = 0
+ cj = 0.00117705
+ ef = 1.064
+ k1 = 0.5470301
+ k2 = 0.038870510000000004
+ k3 = 0.0
+ em = 30000000.0
+ js = 2.5e-7
+ ll = 0.0
+ mj = 0.4476
+ lw = 0.0
+ u0 = 0.0097231258
+ pb = 0.895226
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ua = 1.2617201e-9
+ ub = 5.00396e-20
+ uc = -1.5373321e-10
+ wl = 0.0
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -2e-8
+ ww = 0.0
+ tcjswg = 0.0004130718
+ xw = 0.0
+ tcjsw = 0.0004130718
+ pkt1 = 2.5501714e-15
+ pkt2 = -4.817884e-16
+ keta = 0.04769481
+ pvoff = 2.6840621e-15
+ dsub = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 1.8966694548261387e-25
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ pnfactor = 0
+ wketa = -8.167253e-9
+ pvth0 = -4.826672e-15
+ wnfactor = 0.0
+ voff = -0.1259132
+ drout = 0.0
+ ldif = 9e-8
+ tpbsw = 0.001572025
+ kt1l = 0.0
+ prwb = 0.0
+ pub1 = 5.158311e-32
+ prwg = 0.0
+ puc1 = -2.0035212e-23
+ eta0 = 5e-5
+ cjswg = 4.43205e-10
+ pvag = 0.0
+ etab = -5e-5
+ vsat = 151306.8
+ mjswg = 0.3683619
+ wint = 5e-9
+ pute = -4.378173e-14
+ vth0 = -0.4717293
+ rdsw = 530.0
+ lnfactor = -3.9543e-9
+ wvoff = -1.590053e-9
+ wkt1 = 3.574256e-9
+ wkt2 = 2.0011981e-9
+ lint = 1.4999999e-8
+ wmax = 5e-7
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ wmin = 2.2e-7
+ lkt1 = -1.0417262e-8
+ lkt2 = -1.6001408e-9
+ weta0 = 0
+ nfactor = 1.0
+ lmax = 1e-5
+ pscbe1 = 180397700.0
+ pscbe2 = 5e-7
+ wvsat = 0.0
+ lmin = 1.2e-6
+ lpclm = 2.6005691e-7
+ wvth0 = 8.52019e-9
+ lpdiblc2 = 5.201136e-9
+ ags = 0.02
+ nqsmod = 0
+ )

.model pch_fs_15 pmos (
+ level = 49
+ ute = -0.5904401
+ wk1 = 4.182789e-8
+ wk2 = -2.2085489e-8
+ beta0 = 22.67827
+ wln = 1.0
+ wu0 = -4.185056e-10
+ pkt1 = -8.599671e-15
+ pkt2 = 1.9347028e-16
+ lpdiblc2 = 3.696429e-9
+ keta = 0.0004484208
+ wua = -1.9008923e-16
+ leta0 = 3.6964281896669455e-11
+ wub = 8.369847e-27
+ wuc = 5.370726e-18
+ wwl = 0.0
+ wwn = 1.0
+ letab = -3.696428e-11
+ xti = 3
+ mobmod = 1
+ lvsat = -0.007392816
+ dsub = 0.0
+ lvth0 = -1.9486833e-8
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ delta = 0.01
+ lcit = 2.2622144e-10
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ voff = -0.1186655
+ ldif = 9e-8
+ kt1l = 0.0
+ prwb = 0.0
+ pub1 = -1.2589071e-33
+ prwg = 0.0
+ puc1 = 4.27717e-24
+ eta0 = 1.7857146e-5
+ pvag = 0.0
+ etab = -1.7857146e-5
+ vsat = 146428.52
+ wint = 5e-9
+ pute = -8.783067e-15
+ vth0 = -0.46223000000000003
+ rdsw = 530.0
+ pketa = -5.090041e-15
+ wkt1 = 1.3269771e-8
+ wkt2 = 1.4140165e-9
+ lint = 1.4999999e-8
+ wmax = 5e-7
+ tcjswg = 0.0004130718
+ wmin = 2.2e-7
+ lkt1 = 1.1386779e-8
+ lkt2 = -8.841858e-10
+ lmax = 1.2e-6
+ lmin = 5e-7
+ tcjsw = 0.0004130718
+ nfactor = 1.0
+ pvoff = 3.95383e-15
+ wub1 = 4.292976e-26
+ cdscb = 0.0
+ wuc1 = -3.165437e-17
+ cdscd = 0.0
+ peta0 = 1.8966694548261387e-25
+ hdif = 2e-7
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0017857139
+ pdiblcb = 0.01
+ lub1 = -9.299159e-27
+ wketa = 1.1519229e-8
+ luc1 = 4.434689e-18
+ pvth0 = -4.239814e-16
+ wute = -1.9135335e-8
+ mjsw = 0.3683619
+ drout = 0.0
+ tpbsw = 0.001572025
+ lute = -1.2362289e-9
+ cjswg = 4.43205e-10
+ binunit = 2
+ mjswg = 0.3683619
+ ags = 0.02
+ cdsc = 0.0
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ wvoff = -2.6941984e-9
+ cit = -0.00029671428
+ cgdo = 3.28e-10
+ pscbe1 = 349999900.0
+ pscbe2 = 5e-7
+ dlc = 2e-9
+ cgso = 3.28e-10
+ k3b = 0.0
+ weta0 = 0
+ dwb = 0.0
+ dwg = 0.0
+ wvsat = 0.0
+ lpclm = 1.4785714e-7
+ wvth0 = 4.691763999999999e-9
+ nqsmod = 0
+ a0 = 1.1508681
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ tpbswg = 0.001572025
+ cjsw = 2.60505e-10
+ noimod = 2
+ at = 10000.0
+ cf = 0
+ cj = 0.00117705
+ ef = 1.064
+ k1 = 0.510219
+ k2 = 0.0596423
+ k3 = 0.0
+ em = 30000000.0
+ js = 2.5e-7
+ ll = 0.0
+ noia = 9.5e+18
+ mj = 0.4476
+ noib = 100000.0
+ noic = 1.4e-12
+ lw = 0.0
+ u0 = 0.0091479268
+ pb = 0.895226
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ua = 1.0922192e-9
+ ub = 2.0536515e-20
+ uc = -2.183638e-10
+ la0 = 1.2687106e-7
+ wl = 0.0
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ jsw = 1.2e-12
+ version = 3.24
+ kt1 = -0.2426738
+ lk1 = -6.473878e-9
+ kt2 = -0.027530843
+ lk2 = 6.009272e-10
+ llc = -0.039
+ lln = -1
+ pnfactor = 0
+ lu0 = 2.823877e-10
+ tnom = 25.0
+ lua = 1.6252487e-16
+ lub = 3.353441e-26
+ luc = 5.502275e-18
+ nch = 3.9e+17
+ wnfactor = 0.0
+ lwl = 0.0
+ lwn = 1.0
+ pa0 = 5.971399e-14
+ nlx = 0.0
+ toxm = 4.08e-9
+ lketa = 8.708591e-9
+ pk1 = -1.0521005e-14
+ pk2 = 5.669729e-15
+ pbsw = 0.895226
+ pclm = 0.6714286
+ pu0 = -1.384194e-16
+ xpart = 1
+ prt = 0
+ pua = -5.973716e-23
+ pub = -9.521269e-33
+ puc = -8.311478e-24
+ rsh = 7.2
+ lnfactor = -3.9543e-9
+ tcj = 0.0009739001
+ ua1 = 1.224e-9
+ ub1 = -1.4562286e-18
+ uc1 = 1.3909653e-10
+ pbswg = 0.895226
+ capmod = 3
+ tpb = 0.001572025
+ tox = 4.08e-9
+ wa0 = -1.0502199e-7
+ lvoff = -1.2305139000000001e-8
+ )

.model pch_fs_16 pmos (
+ level = 49
+ cdsc = 0.0
+ binunit = 2
+ pketa = 7.45672e-16
+ lnfactor = -3.9543e-9
+ tcjswg = 0.0004130718
+ cgdo = 3.28e-10
+ wpclm = 4.634222e-9
+ cgso = 3.28e-10
+ tcjsw = 0.0004130718
+ lpdiblc2 = 1.8281252e-9
+ cjsw = 2.60505e-10
+ pvoff = 1.4541431e-15
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ wcdscd = -1.4183201e-11
+ ags = 0.03625
+ cdscb = 0.0
+ cdscd = -6.449223e-5
+ peta0 = 1.8966694548261387e-25
+ cit = 8.534377e-5
+ tnom = 25.0
+ wketa = -1.4490222e-9
+ pvth0 = -1.47043808e-15
+ version = 3.24
+ dlc = 2e-9
+ drout = 0.0
+ pcdscd = 6.382441e-18
+ tpbsw = 0.001572025
+ k3b = 0.0
+ toxm = 4.08e-9
+ dwb = 0.0
+ dwg = 0.0
+ pbsw = 0.895226
+ pclm = 0.9648299
+ cjswg = 4.43205e-10
+ mjswg = 0.3683619
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ wvoff = 2.8606606e-9
+ pscbe1 = 350000000.0
+ pscbe2 = 5e-7
+ la0 = 7.233052e-9
+ jsw = 1.2e-12
+ kt1 = -0.2130934
+ lk1 = 1.3789155e-8
+ kt2 = -0.03589084
+ lk2 = -1.920656e-9
+ llc = -0.039
+ weta0 = 0
+ lln = -1
+ lu0 = -4.357122e-10
+ nqsmod = 0
+ lua = -2.6402067e-16
+ lub = 2.6345733e-25
+ luc = 3.340897e-17
+ nch = 3.9e+17
+ wvsat = 0.0
+ tpbswg = 0.001572025
+ lwl = 0.0
+ lwn = 1.0
+ noimod = 2
+ lpclm = 1.5826547e-8
+ pa0 = -6.072043e-15
+ wvth0 = 7.017223000000001e-9
+ nlx = 0.0
+ pkt1 = -9.758805e-16
+ pkt2 = -1.0643102e-15
+ keta = 0.03159368
+ pk1 = 4.122718e-15
+ pk2 = -2.3103772e-15
+ dsub = 0.0
+ pu0 = 1.3574996e-16
+ prt = 0
+ pua = 6.304761e-23
+ pub = -7.522618e-32
+ puc = -8.758834e-24
+ lags = -7.312499e-9
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ rsh = 7.2
+ tcj = 0.0009739001
+ ua1 = 1.224e-9
+ ub1 = -1.4433942e-18
+ uc1 = 2.0396977e-10
+ tpb = 0.001572025
+ tox = 4.08e-9
+ lcit = 5.429531e-11
+ voff = -0.1287204
+ wa0 = 4.116919e-8
+ lcdscd = 2.9021494e-11
+ ldif = 9e-8
+ ute = -0.5893072
+ wk1 = 9.286284e-9
+ kt1l = 0.0
+ wk2 = -4.351921e-9
+ prwb = 0.0
+ pub1 = 1.9106841e-32
+ prwg = 0.0
+ lketa = -5.306775e-9
+ puc1 = 6.153712e-24
+ wln = 1.0
+ wu0 = -1.0277709000000001e-9
+ eta0 = -0.0004687502
+ wua = -4.629443e-16
+ pvag = 0.0
+ wub = 1.5438073e-25
+ wuc = 6.364847e-18
+ etab = 0.0006718753
+ xpart = 1
+ wwl = 0.0
+ wwn = 1.0
+ vsat = 130812.55
+ xti = 3
+ wint = 5e-9
+ pute = 5.968411e-15
+ vth0 = -0.47511210000000004
+ capmod = 3
+ rdsw = 530.0
+ wkt1 = -3.671987e-9
+ wkt2 = 4.209085e-9
+ pbswg = 0.895226
+ lint = 1.4999999e-8
+ wmax = 5e-7
+ wmin = 2.2e-7
+ lvoff = -7.780439e-9
+ lkt1 = -1.9244071e-9
+ lkt2 = 2.877812e-9
+ lmax = 5e-7
+ beta0 = 22.67827
+ lmin = 1.8e-7
+ mobmod = 1
+ leta0 = 2.559375818966695e-10
+ letab = -3.473438e-10
+ lvsat = -0.0003656336
+ nfactor = 1.0
+ lvth0 = -1.3689881e-8
+ ppclm = -2.0853998e-15
+ wub1 = -2.3274574e-27
+ wuc1 = -3.582447e-17
+ delta = 0.01
+ hdif = 2e-7
+ a0 = 1.4167303
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ pnfactor = 0
+ lub1 = -1.5074642e-26
+ luc1 = -2.4758267e-17
+ at = 10000.0
+ cf = 0
+ cj = 0.00117705
+ ef = 1.064
+ k1 = 0.46519
+ dvt0w = 0.0
+ k2 = 0.06524582
+ k3 = 0.0
+ em = 30000000.0
+ wnfactor = 0.0
+ wute = -5.191639e-8
+ dvt1w = 0.0
+ dvt2w = 0.0
+ mjsw = 0.3683619
+ js = 2.5e-7
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.005937499
+ ll = 0.0
+ mj = 0.4476
+ lw = 0.0
+ u0 = 0.0107437038
+ pb = 0.895226
+ w0 = 0.0
+ rd = 0
+ pdiblcb = 0.01
+ rs = 0
+ ua = 2.0400983e-9
+ ub = -4.904033e-19
+ uc = -2.8037866e-10
+ wl = 0.0
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -2e-8
+ ww = 0.0
+ lute = -1.7460413e-9
+ xw = 0.0
+ )

.model pch_sf_1 pmos (
+ level = 49
+ lvth0 = 3.9543e-9
+ cdsc = 0.0
+ binunit = 2
+ pnfactor = 0
+ cgdo = 3.28e-10
+ delta = 0.01
+ wnfactor = 0.0
+ cgso = 3.28e-10
+ dvt0w = 0.0
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ dvt1w = 0.0
+ dvt2w = 0.0
+ pscbe1 = 199999970.0
+ pscbe2 = 5e-7
+ cjsw = 2.35695e-10
+ ags = 0.02
+ lnfactor = 3.9543e-9
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ nqsmod = 0
+ tpbswg = 0.001572025
+ noimod = 2
+ cit = -0.0001
+ dlc = 2e-9
+ tnom = 25.0
+ version = 3.24
+ k3b = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ toxm = 4.08e-9
+ tcjsw = 0.0004130718
+ pbsw = 0.895226
+ pclm = 0.6000001
+ pvoff = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ jsw = 1.2e-12
+ peta0 = 4.7451600189666944e-17
+ kt1 = -0.2311294
+ lk2 = -1.18629e-9
+ kt2 = -0.02433992
+ llc = -0.039
+ lln = -1
+ lu0 = 7.9086e-11
+ nch = 3.9e+17
+ pvth0 = 1.18629e-15
+ lwl = 0.0
+ lwn = 1.0
+ drout = 0.0
+ nlx = 0.0
+ tpbsw = 0.001572025
+ capmod = 3
+ keta = 0.026632193
+ pu0 = 0.0
+ cjswg = 4.00995e-10
+ prt = 0
+ dsub = 0.0
+ mjswg = 0.3683619
+ rsh = 7.2
+ tcj = 0.0009739001
+ ua1 = 1.224e-9
+ ub1 = -1.3928839e-18
+ uc1 = -4.59467e-12
+ wvoff = 0.0
+ mobmod = 1
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ tpb = 0.001572025
+ tox = 4.08e-9
+ ute = -0.8288856
+ voff = -0.1275921
+ weta0 = 0
+ ldif = 9e-8
+ wvsat = 0.0
+ wln = 1.0
+ kt1l = 0.0
+ prwb = 0.0
+ wu0 = 1.97715e-11
+ prwg = 0.0
+ wvth0 = 1.18629e-9
+ wwl = 0.0
+ wwn = 1.0
+ eta0 = 5e-5
+ xti = 3
+ pvag = 0.0
+ etab = -5e-5
+ vsat = 149999.98
+ wint = 5e-9
+ vth0 = -0.4147553
+ rdsw = 530.0
+ lint = 1.4999999e-8
+ wmax = 0.000900001
+ wmin = 1e-5
+ a0 = 1.0461572
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ lmax = 2.0001e-5
+ at = 10000.0
+ cf = 0
+ cj = 0.00106495
+ lmin = 1e-5
+ ef = 1.064
+ k1 = 0.5375325
+ k2 = 0.029496539999999998
+ k3 = 0.0
+ em = 30000000.0
+ tcjswg = 0.0004130718
+ js = 2.5e-7
+ ll = 0.0
+ mj = 0.4476
+ lw = 0.0
+ u0 = 0.0109204782
+ pb = 0.895226
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ua = 8.23294e-10
+ ub = 6.854322e-19
+ uc = -8.655411e-11
+ wl = 0.0
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ xpart = 1
+ nfactor = 1.0
+ pbswg = 0.895226
+ hdif = 2e-7
+ lvoff = 1.5817200000000002e-9
+ mjsw = 0.3683619
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0010000003
+ pdiblcb = 0.01
+ beta0 = 22.67827
+ leta0 = 4.745160018966694e-10
+ )

.model pch_sf_2 pmos (
+ level = 49
+ mj = 0.4476
+ lw = 0.0
+ kt1 = -0.2295883
+ lk1 = 1.8783622e-8
+ kt2 = -0.024031118
+ lk2 = -6.673462e-9
+ u0 = 0.0110505252
+ pb = 0.895226
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ua = 8.625313e-10
+ ub = 6.401998e-19
+ uc = -8.855145e-11
+ llc = -0.039
+ lln = -1
+ wl = 0.0
+ lu0 = -1.2148829000000001e-9
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ voff = -0.1274002
+ lua = -3.904111e-16
+ lub = 4.500626e-25
+ luc = 1.9873557e-17
+ ldif = 9e-8
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ kt1l = 0.0
+ tcjsw = 0.0004130718
+ prwb = 0.0
+ prwg = 0.0
+ nlx = 0.0
+ eta0 = 5e-5
+ pvag = 0.0
+ etab = -5e-5
+ pvoff = 0.0
+ vsat = 151306.8
+ pu0 = 0.0
+ wint = 5e-9
+ prt = 0
+ vth0 = -0.4122614
+ rdsw = 530.0
+ pnfactor = 0
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 4.7451600189666944e-17
+ lint = 1.4999999e-8
+ rsh = 7.2
+ tcj = 0.0009739001
+ ua1 = 1.224e-9
+ wnfactor = 0.0
+ wmax = 0.000900001
+ ub1 = -1.3977103e-18
+ uc1 = -6.694918e-12
+ wmin = 1e-5
+ tpb = 0.001572025
+ capmod = 3
+ pvth0 = 1.18629e-15
+ tox = 4.08e-9
+ lkt1 = -1.5333228e-8
+ lkt2 = -3.0725886e-9
+ drout = 0.0
+ lmax = 1e-5
+ tpbsw = 0.001572025
+ ute = -0.8385549
+ lmin = 1.2e-6
+ wln = 1.0
+ wu0 = 1.97715e-11
+ cjswg = 4.00995e-10
+ wwl = 0.0
+ wwn = 1.0
+ mjswg = 0.3683619
+ lnfactor = 3.9543e-9
+ xti = 3
+ mobmod = 1
+ nfactor = 1.0
+ wvoff = 0.0
+ hdif = 2e-7
+ lub1 = 4.802326e-26
+ luc1 = 2.0897466e-17
+ weta0 = 0
+ mjsw = 0.3683619
+ lpdiblc2 = 5.201137e-9
+ wvsat = 0.0
+ lute = 9.620972e-8
+ lpclm = 2.6005682e-7
+ wvth0 = 1.18629e-9
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0004772727
+ pdiblcb = 0.01
+ lpscbe1 = 195.04263
+ cdsc = 0.0
+ cgdo = 3.28e-10
+ binunit = 2
+ cgso = 3.28e-10
+ tcjswg = 0.0004130718
+ lketa = -2.0462676e-9
+ cjsw = 2.35695e-10
+ xpart = 1
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ pbswg = 0.895226
+ tnom = 25.0
+ lvoff = -3.274108999999997e-10
+ toxm = 4.08e-9
+ beta0 = 22.67827
+ version = 3.24
+ pbsw = 0.895226
+ pclm = 0.5738637
+ leta0 = 4.745160018966694e-10
+ lvsat = -0.013002843
+ lvth0 = -2.0859753e-8
+ ags = 0.02
+ delta = 0.01
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ cit = -0.0001
+ dlc = 2e-9
+ dvt0w = 0.0
+ dvt1w = 0.0
+ pscbe1 = 180397680.0
+ pscbe2 = 5e-7
+ dvt2w = 0.0
+ k3b = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ keta = 0.026837848
+ nqsmod = 0
+ tpbswg = 0.001572025
+ dsub = 0.0
+ noimod = 2
+ a0 = 1.0385712
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ at = 10000.0
+ cf = 0
+ cj = 0.00106495
+ la0 = 7.548124e-8
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ ef = 1.064
+ k1 = 0.5356447
+ k2 = 0.030048010000000003
+ k3 = 0.0
+ em = 30000000.0
+ js = 2.5e-7
+ jsw = 1.2e-12
+ ll = 0.0
+ )

.model pch_sf_3 pmos (
+ level = 49
+ cjswg = 4.00995e-10
+ mjswg = 0.3683619
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ wvoff = 0.0
+ tnom = 25.0
+ weta0 = 0
+ wvsat = 0.0
+ toxm = 4.08e-9
+ a0 = 1.0045335
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ lpclm = 1.4785704e-7
+ wvth0 = 1.18629e-9
+ pbsw = 0.895226
+ pclm = 0.6714287
+ at = 10000.0
+ cf = 0
+ cj = 0.00106495
+ ef = 1.064
+ k1 = 0.5405614
+ k2 = 0.02936555
+ k3 = 0.0
+ em = 30000000.0
+ js = 2.5e-7
+ version = 3.24
+ ll = 0.0
+ mj = 0.4476
+ lw = 0.0
+ u0 = 0.0102799442
+ pb = 0.895226
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ua = 5.26694e-10
+ ub = 1.1734415e-18
+ uc = -4.332115e-11
+ wl = 0.0
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ pnfactor = 0
+ wnfactor = 0.0
+ tcjswg = 0.0004130718
+ lketa = -8.158225e-9
+ keta = 0.03215259
+ xpart = 1
+ dsub = 0.0
+ lnfactor = 3.9543e-9
+ ags = 0.02
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ pbswg = 0.895226
+ lvoff = 6.329375000000001e-10
+ lcit = 2.2402701e-10
+ cit = -0.00029480609
+ voff = -0.1282353
+ lpdiblc2 = 3.696428e-9
+ ldif = 9e-8
+ dlc = 2e-9
+ beta0 = 22.67827
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ k3b = 0.0
+ dwb = 0.0
+ leta0 = 5.114802818966694e-10
+ dwg = 0.0
+ eta0 = 1.7857143e-5
+ letab = -3.696428e-11
+ pvag = 0.0
+ etab = -1.7857143e-5
+ lvsat = -0.007392833
+ vsat = 146428.53
+ wint = 5e-9
+ lvth0 = -2.735142e-9
+ vth0 = -0.42802199999999996
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ rdsw = 530.0
+ delta = 0.01
+ lint = 1.4999999e-8
+ wmax = 0.000900001
+ pscbe1 = 349999900.0
+ pscbe2 = 5e-7
+ la0 = 1.146246e-7
+ wmin = 1e-5
+ jsw = 1.2e-12
+ lkt1 = 1.5747348e-9
+ lkt2 = 9.740028e-10
+ kt1 = -0.2442909
+ lk1 = 1.3129389e-8
+ kt2 = -0.027549893
+ lk2 = -5.888625e-9
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ lmax = 1.2e-6
+ llc = -0.039
+ lln = -1
+ lu0 = -3.287146e-10
+ lmin = 5e-7
+ lua = -4.198125e-18
+ lub = -1.631654e-25
+ luc = -3.214129e-17
+ nch = 3.9e+17
+ nqsmod = 0
+ lwl = 0.0
+ lwn = 1.0
+ tpbswg = 0.001572025
+ noimod = 2
+ nlx = 0.0
+ pu0 = 0.0
+ prt = 0
+ hdif = 2e-7
+ rsh = 7.2
+ tcj = 0.0009739001
+ nfactor = 1.0
+ ua1 = 1.224e-9
+ lub1 = 3.0810812e-26
+ ub1 = -1.3827429e-18
+ luc1 = 2.9752128e-17
+ uc1 = -1.4394627e-11
+ mjsw = 0.3683619
+ tpb = 0.001572025
+ tox = 4.08e-9
+ tcjsw = 0.0004130718
+ lute = 3.654092e-8
+ ute = -0.786669
+ wln = 1.0
+ pvoff = 0.0
+ wu0 = 1.97715e-11
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0017857148
+ wwl = 0.0
+ wwn = 1.0
+ pdiblcb = 0.01
+ cdsc = 0.0
+ xti = 3
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 4.7451600189666944e-17
+ capmod = 3
+ cgdo = 3.28e-10
+ pvth0 = 1.18629e-15
+ cgso = 3.28e-10
+ drout = 0.0
+ binunit = 2
+ tpbsw = 0.001572025
+ cjsw = 2.35695e-10
+ mobmod = 1
+ )

.model pch_sf_4 pmos (
+ level = 49
+ wmin = 1e-5
+ lkt1 = -2.665e-9
+ lkt2 = -2.325577e-10
+ lmax = 5e-7
+ cit = -4.054396e-5
+ lmin = 1.8e-7
+ lketa = -8.307595e-10
+ dlc = 2e-9
+ k3b = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ xpart = 1
+ pbswg = 0.895226
+ hdif = 2e-7
+ lub1 = 2.883988e-26
+ luc1 = -6.846759e-18
+ lvoff = 1.5460040800000002e-9
+ la0 = 1.6196543e-8
+ mjsw = 0.3683619
+ jsw = 1.2e-12
+ kt1 = -0.2348693
+ lk1 = 1.6807924e-8
+ kt2 = -0.024868647
+ lk2 = -7.0625049999999995e-9
+ beta0 = 22.67827
+ nfactor = 1.0
+ llc = -0.039
+ lln = -1
+ lu0 = -1.9861809999999995e-11
+ lute = 1.6013461e-9
+ leta0 = 7.304535218966694e-10
+ lua = -1.5999061e-16
+ lub = 1.2197973e-25
+ luc = 1.8500639e-17
+ nch = 3.9e+17
+ letab = -5.298917e-10
+ lwl = 0.0
+ lwn = 1.0
+ lvsat = -0.0003656265
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ nlx = 0.0
+ lvth0 = -4.286252e-9
+ cdsc = 0.0
+ pscbe1 = 350000000.0
+ pscbe2 = 5e-7
+ pnfactor = 0
+ pu0 = 0.0
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.00796875
+ delta = 0.01
+ a0 = 1.2232625
+ a1 = 0.0
+ a2 = 0.4
+ prt = 0
+ b0 = 0.0
+ b1 = 0.0
+ cgdo = 3.28e-10
+ wnfactor = 0.0
+ pdiblcb = 0.01
+ at = 10000.0
+ cf = 0
+ cj = 0.00106495
+ ef = 1.064
+ k1 = 0.5323869
+ k2 = 0.031974169999999996
+ k3 = 0.0
+ em = 30000000.0
+ cgso = 3.28e-10
+ js = 2.5e-7
+ dvt0w = 0.0
+ dvt1w = 0.0
+ ll = 0.0
+ rsh = 7.2
+ mj = 0.4476
+ dvt2w = 0.0
+ lw = 0.0
+ u0 = 0.0095936042
+ tcj = 0.0009739001
+ nqsmod = 0
+ pb = 0.895226
+ ua1 = 1.224e-9
+ w0 = 0.0
+ ub1 = -1.3783631e-18
+ rd = 0
+ uc1 = 6.693623e-11
+ tpbswg = 0.001572025
+ rs = 0
+ ua = 8.728995e-10
+ ub = 5.397856e-19
+ uc = -1.5585878e-10
+ noimod = 2
+ wl = 0.0
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ tpb = 0.001572025
+ tox = 4.08e-9
+ binunit = 2
+ cjsw = 2.35695e-10
+ ute = -0.7090256
+ lnfactor = 3.9543e-9
+ wln = 1.0
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ wu0 = 1.97715e-11
+ wwl = 0.0
+ wwn = 1.0
+ xti = 3
+ tnom = 25.0
+ lcdscd = 3.65625e-11
+ lpdiblc2 = 9.140626e-10
+ toxm = 4.08e-9
+ tcjsw = 0.0004130718
+ pbsw = 0.895226
+ pclm = 0.9102259
+ pvoff = 0.0
+ capmod = 3
+ version = 3.24
+ cdscb = 0.0
+ cdscd = -8.125e-5
+ peta0 = 4.7451600189666944e-17
+ pvth0 = 1.18629e-15
+ drout = 0.0
+ tpbsw = 0.001572025
+ mobmod = 1
+ keta = 0.015869336
+ cjswg = 4.00995e-10
+ mjswg = 0.3683619
+ dsub = 0.0
+ wvoff = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ weta0 = 0
+ lcit = 1.0960905e-10
+ voff = -0.1302643
+ ldif = 9e-8
+ wvsat = 0.0
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ lpclm = 4.03983e-8
+ wvth0 = 1.18629e-9
+ eta0 = -0.0004687502
+ pvag = 0.0
+ etab = 0.0010775371
+ vsat = 130812.52
+ wint = 5e-9
+ vth0 = -0.4245751
+ rdsw = 530.0
+ tcjswg = 0.0004130718
+ lint = 1.4999999e-8
+ wmax = 0.000900001
+ ags = 0.02
+ )

.model pch_sf_5 pmos (
+ level = 49
+ wa0 = -4.787191e-8
+ pscbe1 = 199999970.0
+ pscbe2 = 5e-7
+ ute = -0.8394966
+ lvth0 = 3.9543e-9
+ wk1 = 1.2456701e-8
+ wk2 = -5.940143e-9
+ wln = 1.0
+ wu0 = -1.2297032e-9
+ delta = 0.01
+ wua = 1.7543858e-16
+ wub = -6.530953e-25
+ wuc = -7.950096e-17
+ wwl = 0.0
+ wwn = 1.0
+ nqsmod = 0
+ xti = 3
+ version = 3.24
+ tpbswg = 0.001572025
+ noimod = 2
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ keta = 0.02600144
+ dsub = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ voff = -0.1274889
+ ldif = 9e-8
+ tcjsw = 0.0004130718
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ eta0 = 5e-5
+ pvoff = 0.0
+ capmod = 3
+ pvag = 0.0
+ etab = -5e-5
+ vsat = 149999.98
+ wint = 5e-9
+ vth0 = -0.41604359999999996
+ cdscb = 0.0
+ rdsw = 530.0
+ cdscd = 0.0
+ pnfactor = 0
+ peta0 = 4.7451600189666944e-17
+ wkt1 = 8.228274e-9
+ wkt2 = 1.4868883e-9
+ lint = 1.4999999e-8
+ wnfactor = 0.0
+ wmax = 1e-5
+ wketa = 6.301227e-9
+ wmin = 1.2e-6
+ pvth0 = 1.18629e-15
+ mobmod = 1
+ drout = 0.0
+ tpbsw = 0.001572025
+ lmax = 2.0001e-5
+ lmin = 1e-5
+ cjswg = 4.00995e-10
+ a0 = 1.0509492
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ at = 10000.0
+ mjswg = 0.3683619
+ cf = 0
+ cj = 0.00106495
+ lnfactor = 3.9543e-9
+ ef = 1.064
+ k1 = 0.5362856
+ k2 = 0.03009115
+ k3 = 0.0
+ em = 30000000.0
+ js = 2.5e-7
+ ll = 0.0
+ mj = 0.4476
+ lw = 0.0
+ u0 = 0.0110455512
+ pb = 0.895226
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ wvoff = -1.0305298e-9
+ ua = 8.057326e-10
+ ub = 7.508071e-19
+ uc = -7.859605e-11
+ wub1 = 6.909715e-26
+ wuc1 = 3.0354498e-17
+ wl = 0.0
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ hdif = 2e-7
+ weta0 = 0
+ ags = 0.02
+ wute = 1.0600407e-7
+ mjsw = 0.3683619
+ wvsat = 0.0
+ wvth0 = 1.4056747999999999e-8
+ cit = -0.0001
+ dlc = 2e-9
+ nfactor = 1.0
+ k3b = 0.0
+ tcjswg = 0.0004130718
+ dwb = 0.0
+ dwg = 0.0
+ cdsc = 0.0
+ cgdo = 3.28e-10
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0010000004
+ cgso = 3.28e-10
+ pdiblcb = 0.01
+ jsw = 1.2e-12
+ kt1 = -0.231953
+ kt2 = -0.024488758
+ lk2 = -1.18629e-9
+ llc = -0.039
+ lln = -1
+ cjsw = 2.35695e-10
+ lu0 = 7.9086e-11
+ xpart = 1
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ binunit = 2
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ nlx = 0.0
+ pbswg = 0.895226
+ pu0 = 0.0
+ prt = 0
+ tnom = 25.0
+ lvoff = 1.5817200000000002e-9
+ rsh = 7.2
+ beta0 = 22.67827
+ toxm = 4.08e-9
+ tcj = 0.0009739001
+ ua1 = 1.224e-9
+ ub1 = -1.3998005e-18
+ uc1 = -7.633158e-12
+ leta0 = 4.745160018966694e-10
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ pbsw = 0.895226
+ pclm = 0.6000001
+ tpb = 0.001572025
+ tox = 4.08e-9
+ )

.model pch_sf_6 pmos (
+ level = 49
+ lub1 = 5.442727e-26
+ luc1 = 1.8276951e-17
+ wute = 1.0644106e-7
+ mjsw = 0.3683619
+ tcjsw = 0.0004130718
+ capmod = 3
+ lute = 9.664497e-8
+ pvoff = -4.403278e-15
+ nfactor = 1.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 4.7451600189666944e-17
+ mobmod = 1
+ cgdo = 3.28e-10
+ wketa = 7.084359e-9
+ pvth0 = -4.150182e-15
+ cgso = 3.28e-10
+ drout = 0.0
+ tpbsw = 0.001572025
+ ags = 0.02
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0004772728
+ pdiblcb = 0.01
+ lpscbe1 = 195.04262
+ cjswg = 4.00995e-10
+ cit = -0.0001
+ cjsw = 2.35695e-10
+ mjswg = 0.3683619
+ dlc = 2e-9
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ k3b = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ wvoff = -5.879894e-10
+ binunit = 2
+ tnom = 25.0
+ weta0 = 0
+ wvsat = 0.0
+ toxm = 4.08e-9
+ lpclm = 2.6005682e-7
+ wvth0 = 1.4593076e-8
+ la0 = 6.878132e-8
+ pbsw = 0.895226
+ tcjswg = 0.0004130718
+ pclm = 0.5738637
+ jsw = 1.2e-12
+ kt1 = -0.2303147
+ lk1 = 1.8184398e-8
+ kt2 = -0.024155809
+ lk2 = -6.466925e-9
+ llc = -0.039
+ lln = -1
+ lu0 = -1.2264377e-9
+ lua = -3.935608e-16
+ lub = 4.219459e-25
+ luc = 1.8883157e-17
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ pnfactor = 0
+ pa0 = 6.693222e-14
+ nlx = 0.0
+ wnfactor = 0.0
+ pk1 = 5.986243e-15
+ pk2 = -2.063307e-15
+ pu0 = 1.1543239e-16
+ prt = 0
+ pua = 3.1465633e-23
+ pub = 2.8088595e-31
+ puc = 9.8941e-24
+ version = 3.24
+ lketa = -1.2662711e-9
+ rsh = 7.2
+ pkt1 = 9.666697e-15
+ tcj = 0.0009739001
+ pkt2 = 2.4000725e-15
+ ua1 = 1.224e-9
+ keta = 0.026128704
+ ub1 = -1.4052706e-18
+ uc1 = -9.470036e-12
+ xpart = 1
+ tpb = 0.001572025
+ lnfactor = 3.9543e-9
+ tox = 4.08e-9
+ dsub = 0.0
+ wa0 = -5.459876e-8
+ ute = -0.8492097
+ wk1 = 1.185507e-8
+ wk2 = -5.732776e-9
+ pbswg = 0.895226
+ wln = 1.0
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ wu0 = -1.2413044999999998e-9
+ wua = 1.7227619e-16
+ wub = -6.81325e-25
+ wuc = -8.049533e-17
+ wwl = 0.0
+ wwn = 1.0
+ a0 = 1.0440365
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ lvoff = 1.1335760000000018e-10
+ xti = 3
+ at = 10000.0
+ cf = 0
+ lpdiblc2 = 5.201137e-9
+ cj = 0.00106495
+ voff = -0.1273414
+ ef = 1.064
+ k1 = 0.534458
+ k2 = 0.03062187
+ k3 = 0.0
+ em = 30000000.0
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ ldif = 9e-8
+ beta0 = 22.67827
+ js = 2.5e-7
+ ll = 0.0
+ mj = 0.4476
+ lw = 0.0
+ u0 = 0.0111767602
+ pb = 0.895226
+ kt1l = 0.0
+ w0 = 0.0
+ prwb = 0.0
+ rd = 0
+ pub1 = -6.397619e-32
+ prwg = 0.0
+ leta0 = 4.745160018966694e-10
+ puc1 = 2.6178952e-23
+ rs = 0
+ ua = 8.452865e-10
+ ub = 7.084005e-19
+ uc = -8.049386e-11
+ pscbe1 = 180397700.0
+ pscbe2 = 5e-7
+ wl = 0.0
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ eta0 = 5e-5
+ lvsat = -0.013002842
+ pvag = 0.0
+ etab = -5e-5
+ vsat = 151306.8
+ lvth0 = -2.0325569e-8
+ wint = 5e-9
+ pute = -4.348101e-15
+ vth0 = -0.41360349999999996
+ nqsmod = 0
+ rdsw = 530.0
+ tpbswg = 0.001572025
+ delta = 0.01
+ wkt1 = 7.256747e-9
+ wkt2 = 1.245675e-9
+ noimod = 2
+ lint = 1.4999999e-8
+ wmax = 1e-5
+ wmin = 1.2e-6
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ lkt1 = -1.6300865e-8
+ lkt2 = -3.312836e-9
+ lmax = 1e-5
+ lmin = 1.2e-6
+ pketa = -7.792167e-15
+ wub1 = 7.552692e-26
+ wuc1 = 2.7723443e-17
+ hdif = 2e-7
+ )

.model pch_sf_7 pmos (
+ level = 49
+ mjswg = 0.3683619
+ jsw = 1.2e-12
+ kt1 = -0.2459144
+ lk1 = 8.371453e-9
+ kt2 = -0.027846618
+ lk2 = -4.402144e-9
+ dsub = 0.0
+ llc = -0.039
+ lln = -1
+ lu0 = -2.666366e-10
+ wvoff = -7.866491e-9
+ lua = 3.0792715e-17
+ lub = -1.9665828e-25
+ luc = -3.700045e-17
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ wcit = -1.788104e-11
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ pa0 = -1.2519753e-13
+ nlx = 0.0
+ weta0 = 0
+ pk1 = 4.753178e-14
+ pk2 = -1.4849934e-14
+ lcit = 2.2196864e-10
+ voff = -0.1274479
+ pu0 = -6.201592e-16
+ wvsat = 0.0
+ ldif = 9e-8
+ tcjswg = 0.0004130718
+ prt = 0
+ pua = -3.495584e-22
+ pub = 3.345938e-31
+ puc = 4.854297e-23
+ lpclm = 1.4785702e-7
+ wvth0 = 1.1317e-8
+ kt1l = 0.0
+ prwb = 0.0
+ pub1 = -1.382964e-31
+ prwg = 0.0
+ puc1 = -5.043768e-23
+ eta0 = 1.7857139e-5
+ rsh = 7.2
+ tcj = 0.0009739001
+ ua1 = 1.224e-9
+ pvag = 0.0
+ ub1 = -1.3967723e-18
+ etab = -1.7857139e-5
+ uc1 = -2.3838735e-11
+ vsat = 146428.53
+ wint = 5e-9
+ pute = 2.0900147e-14
+ tpb = 0.001572025
+ tox = 4.08e-9
+ vth0 = -0.4290361
+ wa0 = 1.1247056e-7
+ rdsw = 530.0
+ ute = -0.7951261
+ wkt1 = 1.6218328e-8
+ wkt2 = 2.9642964e-9
+ wk1 = -2.4271484e-8
+ wk2 = 5.386031e-9
+ lint = 1.4999999e-8
+ wmax = 1e-5
+ wln = 1.0
+ wu0 = -6.016596e-10
+ wmin = 1.2e-6
+ wua = 5.036014e-16
+ wub = -7.280275e-25
+ wuc = -1.1410304e-16
+ lkt1 = 1.6387112e-9
+ lkt2 = 9.315946e-10
+ wwl = 0.0
+ wwn = 1.0
+ xti = 3
+ lmax = 1.2e-6
+ lketa = -8.380984e-9
+ lmin = 5e-7
+ xpart = 1
+ wub1 = 1.4015321e-25
+ pbswg = 0.895226
+ wuc1 = 9.434661e-17
+ hdif = 2e-7
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ lvoff = 2.3584050000000025e-10
+ lub1 = 4.46543e-26
+ luc1 = 3.480094e-17
+ wute = 8.448607e-8
+ mjsw = 0.3683619
+ pscbe1 = 349999900.0
+ pscbe2 = 5e-7
+ beta0 = 22.67827
+ leta0 = 5.114802918966694e-10
+ lute = 3.444881e-8
+ letab = -3.696429e-11
+ lvsat = -0.007392833
+ lvth0 = -2.5780870000000004e-9
+ nqsmod = 0
+ tpbswg = 0.001572025
+ noimod = 2
+ cdsc = 0.0
+ pnfactor = 0
+ delta = 0.01
+ wnfactor = 0.0
+ cgdo = 3.28e-10
+ nfactor = 1.0
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ cgso = 3.28e-10
+ cjsw = 2.35695e-10
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0017857144
+ lnfactor = 3.9543e-9
+ pdiblcb = 0.01
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ pketa = 2.2253538e-15
+ tnom = 25.0
+ binunit = 2
+ capmod = 3
+ lpdiblc2 = 3.696428e-9
+ tcjsw = 0.0004130718
+ toxm = 4.08e-9
+ ags = 0.02
+ pcit = 2.0563189e-17
+ pbsw = 0.895226
+ pclm = 0.6714287
+ pvoff = 3.966999e-15
+ cit = -0.0002930162
+ a0 = 0.9932752
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ at = 10000.0
+ mobmod = 1
+ cf = 0
+ dlc = 2e-9
+ cj = 0.00106495
+ ef = 1.064
+ k1 = 0.542991
+ k2 = 0.0288264
+ k3 = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ em = 30000000.0
+ peta0 = 4.7451600189666944e-17
+ k3b = 0.0
+ js = 2.5e-7
+ ll = 0.0
+ mj = 0.4476
+ lw = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ u0 = 0.0103421492
+ pb = 0.895226
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ua = 4.762835e-10
+ ub = 1.2463172e-18
+ uc = -3.189942e-11
+ wl = 0.0
+ wr = 1.0
+ xj = 1.7000001e-7
+ wketa = -1.6265284e-9
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ pvth0 = -3.826928e-16
+ drout = 0.0
+ tpbsw = 0.001572025
+ pkt1 = -6.391237e-16
+ pkt2 = 4.236579e-16
+ keta = 0.03231541
+ cjswg = 4.00995e-10
+ version = 3.24
+ la0 = 1.2715688e-7
+ )

.model pch_sf_8 pmos (
+ level = 49
+ cgso = 3.28e-10
+ nfactor = 1.0
+ a0 = 1.2640158
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ lketa = -5.872592e-10
+ at = 10000.0
+ cf = 0
+ cj = 0.00106495
+ ef = 1.064
+ k1 = 0.5203763
+ k2 = 0.036403239999999996
+ k3 = 0.0
+ em = 30000000.0
+ pcdscd = -7.408954e-18
+ js = 2.5e-7
+ ll = 0.0
+ mj = 0.4476
+ lw = 0.0
+ u0 = 0.0098511212
+ pb = 0.895226
+ xpart = 1
+ w0 = 0.0
+ rd = 0
+ cjsw = 2.35695e-10
+ rs = 0
+ ua = 9.357863e-10
+ ub = 5.091257e-19
+ uc = -1.5731644e-10
+ wl = 0.0
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.007987866
+ pbswg = 0.895226
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ pdiblcb = 0.01
+ pscbe1 = 350000000.0
+ pscbe2 = 5e-7
+ lvoff = 1.7452549500000003e-9
+ tnom = 25.0
+ pags = -6.875222e-16
+ beta0 = 22.67827
+ toxm = 4.08e-9
+ binunit = 2
+ leta0 = 7.304535218966694e-10
+ letab = -5.545772e-10
+ nqsmod = 0
+ pcit = -7.907631e-17
+ pbsw = 0.895226
+ pclm = 0.9107697
+ tpbswg = 0.001572025
+ lvsat = -0.0003656271
+ noimod = 2
+ lvth0 = -4.173726e-9
+ ppclm = 2.4445072e-15
+ delta = 0.01
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ lcdscd = 3.730414e-11
+ pkt1 = -1.8229216e-15
+ pkt2 = -1.2254391e-15
+ keta = 0.014996022
+ ags = 0.019847063
+ wags = 1.5278273e-9
+ dsub = 0.0
+ version = 3.24
+ cit = -6.09184e-5
+ pketa = -2.4325694e-15
+ dlc = 2e-9
+ lags = 6.882101e-11
+ wcit = 2.0354016e-10
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ k3b = 0.0
+ capmod = 3
+ dwb = 0.0
+ dwg = 0.0
+ wpclm = -5.432238e-9
+ lcit = 1.1752459e-10
+ voff = -0.1308021
+ tcjsw = 0.0004130718
+ ldif = 9e-8
+ kt1l = 0.0
+ prwb = 0.0
+ pub1 = 2.7781507e-32
+ prwg = 0.0
+ puc1 = 8.113434e-24
+ pvoff = -1.9905158e-15
+ eta0 = -0.0004687502
+ mobmod = 1
+ pvag = 0.0
+ etab = 0.0011323938
+ la0 = 5.323636e-9
+ vsat = 130812.52
+ wint = 5e-9
+ pute = 9.798417e-15
+ jsw = 1.2e-12
+ kt1 = -0.2367561
+ lk1 = 1.854804e-8
+ kt2 = -0.025532207
+ lk2 = -7.811716e-9
+ vth0 = -0.4254902
+ cdscb = 0.0
+ cdscd = -8.289813e-5
+ pnfactor = 0
+ peta0 = 4.7451600189666944e-17
+ llc = -0.039
+ rdsw = 530.0
+ lln = -1
+ lu0 = -4.5673330000000005e-11
+ petab = 2.4660761e-16
+ wnfactor = 0.0
+ wkt1 = 1.8848993e-8
+ wkt2 = 6.628956e-9
+ lua = -1.759835e-16
+ lub = 1.3507784e-25
+ luc = 1.9437196e-17
+ lint = 1.4999999e-8
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ wmax = 1e-5
+ wketa = 8.724413e-9
+ pvth0 = 6.215440000000003e-17
+ pa0 = 1.0862038e-13
+ nlx = 0.0
+ wmin = 1.2e-6
+ drout = 0.0
+ lkt1 = -2.4825255e-9
+ lkt2 = -1.0989117e-10
+ tpbsw = 0.001572025
+ pk1 = -1.7383759e-14
+ pk2 = 7.484627e-15
+ lmax = 5e-7
+ pu0 = 2.5785697e-16
+ lmin = 1.8e-7
+ ppdiblc2 = 8.594017e-17
+ prt = 0
+ pua = 1.5976873e-22
+ pub = -1.3085017e-31
+ puc = -9.356197e-24
+ cjswg = 4.00995e-10
+ wpdiblc2 = -1.9097854e-10
+ mjswg = 0.3683619
+ lnfactor = 3.9543e-9
+ rsh = 7.2
+ tcj = 0.0009739001
+ ua1 = 1.224e-9
+ ub1 = -1.3554493e-18
+ uc1 = 7.051652e-11
+ wvoff = 5.372431e-9
+ tpb = 0.001572025
+ tox = 4.08e-9
+ wub1 = -2.2890885e-25
+ wuc1 = -3.576699e-17
+ wa0 = -4.071248e-7
+ hdif = 2e-7
+ ute = -0.7199521
+ wk1 = 1.1998529e-7
+ wk2 = -4.424634e-8
+ weta0 = 0
+ tcjswg = 0.0004130718
+ lub1 = 2.6058948e-26
+ luc1 = -7.658915e-18
+ wln = 1.0
+ wetab = -5.480169e-10
+ lpdiblc2 = 9.0546e-10
+ wu0 = -2.5528067e-9
+ wute = 1.0915658e-7
+ mjsw = 0.3683619
+ wvsat = 0.0
+ wua = -6.282368e-16
+ wub = 3.0629255e-25
+ wuc = 1.4561782e-17
+ wwl = 0.0
+ wwn = 1.0
+ lpclm = 4.015361e-8
+ wvth0 = 1.0328453999999999e-8
+ xti = 3
+ lute = 6.205235e-10
+ cdsc = 0.0
+ wcdscd = 1.6464351e-11
+ cgdo = 3.28e-10
+ )

.model pch_sf_9 pmos (
+ level = 49
+ pvag = 0.0
+ etab = -5e-5
+ lvth0 = 3.9543e-9
+ ags = 0.02
+ vsat = 149999.98
+ wint = 5e-9
+ vth0 = -0.40491299999999997
+ delta = 0.01
+ rdsw = 530.0
+ cit = -0.0001
+ wkt1 = 6.74333e-9
+ wkt2 = 1.2948118e-10
+ lint = 1.4999999e-8
+ dlc = 2e-9
+ wmax = 1.2e-6
+ dvt0w = 0.0
+ k3b = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ wmin = 5e-7
+ dwb = 0.0
+ dwg = 0.0
+ lmax = 2.0001e-5
+ lmin = 1e-5
+ capmod = 3
+ a0 = 0.9810578
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ jsw = 1.2e-12
+ kt1 = -0.2307052
+ kt2 = -0.02334808
+ lk2 = -1.18629e-9
+ wub1 = 3.495163e-26
+ wuc1 = 1.9335648e-17
+ at = 10000.0
+ cf = 0
+ cj = 0.00106495
+ ef = 1.064
+ k1 = 0.5449055
+ k2 = 0.02831336
+ k3 = 0.0
+ em = 30000000.0
+ llc = -0.039
+ lln = -1
+ lu0 = 7.9086e-11
+ hdif = 2e-7
+ js = 2.5e-7
+ ll = 0.0
+ mj = 0.4476
+ lw = 0.0
+ u0 = 0.0101875252
+ nch = 3.9e+17
+ pb = 0.895226
+ w0 = 0.0
+ rd = 0
+ lwl = 0.0
+ lwn = 1.0
+ rs = 0
+ ua = 1.0698959e-9
+ ub = 3.0837888e-19
+ uc = -1.1659398e-10
+ wl = 0.0
+ wute = -2.7886795e-9
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ mjsw = 0.3683619
+ nlx = 0.0
+ tcjsw = 0.0004130718
+ mobmod = 1
+ pu0 = 0.0
+ pvoff = 0.0
+ prt = 0
+ rsh = 7.2
+ cdscb = 0.0
+ cdscd = 0.0
+ tcj = 0.0009739001
+ peta0 = 4.7451600189666944e-17
+ cdsc = 0.0
+ ua1 = 1.224e-9
+ ub1 = -1.3711068e-18
+ uc1 = 1.6263793e-12
+ tpb = 0.001572025
+ tox = 4.08e-9
+ cgdo = 3.28e-10
+ wketa = -1.0458587e-9
+ wa0 = 3.529885e-8
+ pvth0 = 1.18629e-15
+ drout = 0.0
+ ute = -0.7480742
+ wk1 = 2.1990281e-9
+ cgso = 3.28e-10
+ wk2 = -3.824582e-9
+ tpbsw = 0.001572025
+ wln = 1.0
+ wu0 = -2.086521e-10
+ wua = -1.3891575e-16
+ wub = -1.2660565e-25
+ wuc = -3.428342e-17
+ wwl = 0.0
+ wwn = 1.0
+ cjswg = 4.00995e-10
+ nfactor = 1.0
+ xti = 3
+ cjsw = 2.35695e-10
+ mjswg = 0.3683619
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ wvoff = -4.105241e-10
+ tcjswg = 0.0004130718
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0009999998
+ weta0 = 0
+ tnom = 25.0
+ pdiblcb = 0.01
+ wvsat = 0.0
+ wvth0 = 8.112289000000001e-10
+ toxm = 4.08e-9
+ pbsw = 0.895226
+ pclm = 0.6
+ binunit = 2
+ pnfactor = 0
+ wnfactor = 0.0
+ keta = 0.03217546
+ xpart = 1
+ lnfactor = 3.9543e-9
+ alpha0 = 0.0
+ dsub = 0.0
+ alpha1 = 6.8730453846
+ pbswg = 0.895226
+ pscbe1 = 199999970.0
+ pscbe2 = 5e-7
+ dvt0 = 0.0
+ version = 3.24
+ dvt1 = 0.0
+ dvt2 = 0.0
+ lvoff = 1.5817200000000002e-9
+ voff = -0.12801
+ beta0 = 22.67827
+ nqsmod = 0
+ ldif = 9e-8
+ tpbswg = 0.001572025
+ noimod = 2
+ leta0 = 4.745160018966694e-10
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ eta0 = 5e-5
+ )

.model pch_sf_10 pmos (
+ level = 49
+ dsub = 0.0
+ wk1 = 1.7598129e-9
+ wk2 = -3.600003e-9
+ wln = 1.0
+ wu0 = -1.7835274000000001e-10
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ wua = -1.6455617e-16
+ wub = -7.150721e-26
+ wuc = -2.8652769e-17
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ wwl = 0.0
+ wwn = 1.0
+ xti = 3
+ pscbe1 = 180397680.0
+ pscbe2 = 5e-7
+ voff = -0.1269095
+ ldif = 9e-8
+ nfactor = 1.0
+ kt1l = 0.0
+ prwb = 0.0
+ pub1 = -8.629597e-32
+ prwg = 0.0
+ puc1 = 1.5034668e-23
+ nqsmod = 0
+ tpbswg = 0.001572025
+ lketa = -6.417587e-9
+ eta0 = 5e-5
+ noimod = 2
+ pvag = 0.0
+ etab = -5e-5
+ vsat = 151306.8
+ wint = 5e-9
+ pute = 3.909688e-14
+ xpart = 1
+ vth0 = -0.40084529999999996
+ rdsw = 530.0
+ wkt1 = 6.495125e-9
+ wkt2 = 2.3726165e-10
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0004772722
+ lint = 1.4999999e-8
+ pdiblcb = 0.01
+ lpscbe1 = 195.04263
+ wmax = 1.2e-6
+ pbswg = 0.895226
+ wmin = 5e-7
+ lkt1 = -1.0252924e-8
+ lkt2 = -3.947785e-10
+ lmax = 1e-5
+ lvoff = -9.367244999999999e-9
+ lmin = 1.2e-6
+ beta0 = 22.67827
+ binunit = 2
+ leta0 = 4.745160018966694e-10
+ lvsat = -0.013002842
+ lvth0 = -3.651863e-8
+ wub1 = 4.362458e-26
+ wuc1 = 1.7824627e-17
+ capmod = 3
+ hdif = 2e-7
+ delta = 0.01
+ lub1 = 7.318341e-26
+ luc1 = 2.7641896e-17
+ pnfactor = 0
+ wute = -6.718015e-9
+ mjsw = 0.3683619
+ wnfactor = 0.0
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ lute = 6.013659e-8
+ mobmod = 1
+ cdsc = 0.0
+ version = 3.24
+ lnfactor = 3.9543e-9
+ pketa = -1.6621007e-15
+ cgdo = 3.28e-10
+ ags = 0.02
+ cgso = 3.28e-10
+ cit = -0.0001
+ tcjsw = 0.0004130718
+ dlc = 2e-9
+ lpdiblc2 = 5.201137e-9
+ cjsw = 2.35695e-10
+ k3b = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ pvoff = 6.87864e-15
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 4.7451600189666944e-17
+ tcjswg = 0.0004130718
+ tnom = 25.0
+ wketa = -8.788133e-10
+ pvth0 = 1.511956e-14
+ la0 = 1.2176828e-7
+ drout = 0.0
+ toxm = 4.08e-9
+ jsw = 1.2e-12
+ kt1 = -0.2296747
+ lk1 = 1.9542425e-8
+ kt2 = -0.023308404
+ lk2 = -6.323008999999999e-9
+ tpbsw = 0.001572025
+ pbsw = 0.895226
+ llc = -0.039
+ pclm = 0.5738636
+ lln = -1
+ lu0 = -8.760922000000001e-10
+ lua = -5.815077e-16
+ lub = 1.1186816e-24
+ luc = 7.427734e-17
+ nch = 3.9e+17
+ a0 = 0.9688198
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ lwl = 0.0
+ lwn = 1.0
+ cjswg = 4.00995e-10
+ at = 10000.0
+ cf = 0
+ cj = 0.00106495
+ pa0 = 3.87773e-15
+ nlx = 0.0
+ ef = 1.064
+ k1 = 0.5429414
+ k2 = 0.028829620000000004
+ k3 = 0.0
+ em = 30000000.0
+ mjswg = 0.3683619
+ js = 2.5e-7
+ ll = 0.0
+ mj = 0.4476
+ lw = 0.0
+ pk1 = 4.370194e-15
+ pk2 = -2.2345663e-15
+ u0 = 0.0102835232
+ pb = 0.895226
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ua = 1.1283389e-9
+ ub = 1.9594849e-19
+ uc = -1.2405904e-10
+ wvoff = -1.1018445e-9
+ wl = 0.0
+ pu0 = -3.0147877e-16
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ prt = 0
+ pua = 2.5512236e-22
+ pub = -5.482294e-31
+ puc = -5.602498e-23
+ weta0 = 0
+ rsh = 7.2
+ tcj = 0.0009739001
+ ua1 = 1.224e-9
+ ub1 = -1.3784619e-18
+ uc1 = -1.1517035e-12
+ wvsat = 0.0
+ pkt1 = 2.469645e-15
+ pkt2 = -1.0724159e-15
+ keta = 0.03282044
+ tpb = 0.001572025
+ tox = 4.08e-9
+ lpclm = 2.6005682e-7
+ wvth0 = -5.891015e-10
+ wa0 = 3.490912e-8
+ ute = -0.754118
+ )

.model pch_sf_11 pmos (
+ level = 49
+ cgso = 3.28e-10
+ a0 = 1.1936638
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ lvoff = 6.818931000000001e-9
+ at = 10000.0
+ cf = 0
+ cj = 0.00106495
+ ef = 1.064
+ k1 = 0.4715038
+ k2 = 0.05425073
+ k3 = 0.0
+ em = 30000000.0
+ js = 2.5e-7
+ ll = 0.0
+ mj = 0.4476
+ lw = 0.0
+ beta0 = 22.67827
+ u0 = 0.0107824642
+ pb = 0.895226
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ua = 1.036115e-9
+ ub = 1.0523674e-18
+ uc = -7.205117e-11
+ cjsw = 2.35695e-10
+ leta0 = 5.114802618966694e-10
+ wl = 0.0
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ letab = -3.696426e-11
+ lvsat = -0.007392855
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ capmod = 3
+ lvth0 = 3.9159799999999995e-10
+ delta = 0.01
+ tnom = 25.0
+ ags = 0.02
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ toxm = 4.08e-9
+ mobmod = 1
+ pcit = -1.0851648e-17
+ pbsw = 0.895226
+ pclm = 0.6714286
+ cit = -0.00031597191
+ dlc = 2e-9
+ k3b = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ pketa = 4.024799e-15
+ la0 = -1.3680231e-7
+ pkt1 = -6.051915e-15
+ pkt2 = -1.4802061e-15
+ tcjsw = 0.0004130718
+ keta = 0.03584265
+ jsw = 1.2e-12
+ kt1 = -0.2439705
+ lk1 = 1.0169572e-7
+ kt2 = -0.025852976
+ lk2 = -3.555729e-8
+ llc = -0.039
+ lln = -1
+ lu0 = -1.4498735e-9
+ dsub = 0.0
+ pvoff = -3.866879e-15
+ lua = -4.754501e-16
+ lub = 1.337998e-25
+ luc = 1.4468274e-17
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ pa0 = 1.8891395e-13
+ nlx = 0.0
+ tcjswg = 0.0004130718
+ wcit = 9.436221e-12
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ pk1 = -6.35241e-14
+ pk2 = 2.2224691e-14
+ peta0 = 4.7451600189666944e-17
+ pu0 = 7.878928e-16
+ pnfactor = 0
+ prt = 0
+ lcit = 2.4836766e-10
+ pua = 2.5287059e-22
+ pub = -5.865131e-32
+ puc = -1.2704817e-23
+ wketa = -5.823942e-9
+ voff = -0.1409845
+ pvth0 = -3.9166180000000005e-15
+ wnfactor = 0.0
+ ldif = 9e-8
+ drout = 0.0
+ kt1l = 0.0
+ tpbsw = 0.001572025
+ prwb = 0.0
+ pub1 = 4.97241e-32
+ prwg = 0.0
+ rsh = 7.2
+ puc1 = 1.7282469e-23
+ tcj = 0.0009739001
+ ua1 = 1.224e-9
+ ub1 = -1.2162624e-18
+ uc1 = 4.210797e-11
+ eta0 = 1.7857154e-5
+ nfactor = 1.0
+ pvag = 0.0
+ etab = -1.7857154e-5
+ tpb = 0.001572025
+ tox = 4.08e-9
+ cjswg = 4.00995e-10
+ vsat = 146428.56
+ wa0 = -1.2599192e-7
+ wint = 5e-9
+ pute = -5.928695e-14
+ mjswg = 0.3683619
+ vth0 = -0.43294119999999997
+ ute = -0.7903757
+ wk1 = 6.079834e-8
+ wk2 = -2.4868919e-8
+ rdsw = 530.0
+ wln = 1.0
+ wkt1 = 1.3905176e-8
+ wkt2 = 5.918618e-10
+ lnfactor = 3.9543e-9
+ wu0 = -1.1256324e-9
+ lint = 1.4999999e-8
+ wvoff = 8.242083e-9
+ wua = -1.625981e-16
+ wmax = 1.2e-6
+ wub = -4.972273e-25
+ wuc = -6.632247e-17
+ wwl = 0.0
+ wwn = 1.0
+ wmin = 5e-7
+ xti = 3
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0017857137
+ lkt1 = 6.187276e-9
+ lkt2 = 2.5314804e-9
+ pdiblcb = 0.01
+ weta0 = 0
+ lmax = 1.2e-6
+ lmin = 5e-7
+ wvsat = 0.0
+ lpclm = 1.4785714e-7
+ wvth0 = 1.5964097e-8
+ lpdiblc2 = 3.696429e-9
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ binunit = 2
+ pscbe1 = 349999900.0
+ pscbe2 = 5e-7
+ wub1 = -7.465372e-26
+ wuc1 = 1.5870021e-17
+ hdif = 2e-7
+ lub1 = -1.133461e-25
+ luc1 = -2.2106738e-17
+ wute = 7.883313e-8
+ mjsw = 0.3683619
+ nqsmod = 0
+ tpbswg = 0.001572025
+ noimod = 2
+ lute = 1.0183292e-7
+ lketa = -9.893122e-9
+ xpart = 1
+ cdsc = 0.0
+ cgdo = 3.28e-10
+ pbswg = 0.895226
+ version = 3.24
+ )

.model pch_sf_12 pmos (
+ level = 49
+ wint = 5e-9
+ llc = -0.039
+ pute = 1.3160581e-15
+ lln = -1
+ lu0 = 2.9107207000000003e-10
+ vth0 = -0.42263
+ nfactor = 1.0
+ lua = 2.3815556e-17
+ lub = -3.425063e-26
+ luc = 8.803578e-18
+ nch = 3.9e+17
+ rdsw = 530.0
+ lwl = 0.0
+ lwn = 1.0
+ pketa = -9.609158e-16
+ wkt1 = 2.7434011e-10
+ wkt2 = -6.113567e-9
+ lint = 1.4999999e-8
+ pa0 = -8.476619e-14
+ nlx = 0.0
+ wmax = 1.2e-6
+ pk1 = 1.5213101e-14
+ pk2 = -6.235986e-15
+ wmin = 5e-7
+ lkt1 = -4.083267e-9
+ lkt2 = -2.4314675e-9
+ wpclm = 5.671285e-8
+ pu0 = -1.4287007e-16
+ lmax = 5e-7
+ prt = 0
+ pua = -7.799214e-23
+ pub = 7.065072e-32
+ puc = 3.297807e-24
+ lmin = 1.8e-7
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.009150297
+ tcjsw = 0.0004130718
+ pdiblcb = 0.01
+ rsh = 7.2
+ tcj = 0.0009739001
+ ua1 = 1.224e-9
+ ub1 = -1.6175756e-18
+ uc1 = -2.2818641e-11
+ pvoff = -1.4343533e-15
+ tcjswg = 0.0004130718
+ tpb = 0.001572025
+ tox = 4.08e-9
+ a0 = 0.5166956
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ wa0 = 4.821862e-7
+ at = 10000.0
+ cf = 0
+ cj = 0.00106495
+ wub1 = 8.30214e-26
+ ute = -0.5812994
+ wuc1 = 7.530186e-17
+ ef = 1.064
+ k1 = 0.7171482
+ k2 = -0.033028159
+ k3 = 0.0
+ em = 30000000.0
+ wk1 = -1.1417325e-7
+ wk2 = 3.837703e-8
+ binunit = 2
+ cdscb = 0.0
+ cdscd = -5.200001e-5
+ peta0 = 4.7451600189666944e-17
+ js = 2.5e-7
+ ll = 0.0
+ mj = 0.4476
+ hdif = 2e-7
+ lw = 0.0
+ u0 = 0.0069136952
+ wln = 1.0
+ pb = 0.895226
+ w0 = 0.0
+ wu0 = 9.427299e-10
+ rd = 0
+ rs = 0
+ ua = -7.336427e-11
+ ub = 1.4258127e-18
+ uc = -5.946296e-11
+ lub1 = 6.724484e-26
+ wua = 5.726523e-16
+ wub = -7.845651e-25
+ wuc = -1.0188386e-16
+ wl = 0.0
+ luc1 = 7.110234e-18
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ wwl = 0.0
+ wwn = 1.0
+ wute = -5.584022e-8
+ wketa = 5.255423e-9
+ mjsw = 0.3683619
+ pvth0 = 1.5103980000000002e-16
+ xti = 3
+ drout = 0.0
+ tpbsw = 0.001572025
+ lute = 7.748556e-9
+ wcdscd = -2.0304376e-11
+ cjswg = 4.00995e-10
+ mjswg = 0.3683619
+ cdsc = 0.0
+ wvoff = 2.8364715e-9
+ cgdo = 3.28e-10
+ pcdscd = 9.13697e-18
+ cgso = 3.28e-10
+ weta0 = 0
+ version = 3.24
+ wvsat = 0.0
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ lpclm = 6.365384e-8
+ wvth0 = 6.924854999999999e-9
+ cjsw = 2.35695e-10
+ pscbe1 = 350000000.0
+ pscbe2 = 5e-7
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ nqsmod = 0
+ tpbswg = 0.001572025
+ tnom = 25.0
+ pnfactor = 0
+ noimod = 2
+ pags = -5.667374e-15
+ wnfactor = 0.0
+ toxm = 4.08e-9
+ pcit = 2.6834248e-18
+ pbsw = 0.895226
+ lketa = -1.8239428e-9
+ pclm = 0.858547
+ xpart = 1
+ ppdiblc2 = 7.08422e-16
+ wpdiblc2 = -1.5742713e-9
+ lnfactor = 3.9543e-9
+ pbswg = 0.895226
+ lcdscd = 2.3400004e-11
+ lvoff = 1.2778913700000001e-9
+ ags = 0.010547621
+ beta0 = 22.67827
+ pkt1 = 8.196091e-17
+ pkt2 = 1.5372367e-15
+ keta = 0.01791114
+ lpdiblc2 = 3.823661e-10
+ leta0 = 7.304534718966694e-10
+ capmod = 3
+ letab = -3.473438e-10
+ cit = 0.00012746976
+ wags = 1.2594167e-8
+ lvsat = -0.0003656142
+ dsub = 0.0
+ dlc = 2e-9
+ lvth0 = -4.248419000000001e-9
+ k3b = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ lags = 4.253569e-9
+ wcit = -2.0641719e-11
+ ppclm = -2.5520774e-14
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ delta = 0.01
+ mobmod = 1
+ lcit = 4.881893e-11
+ voff = -0.1286711
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ ldif = 9e-8
+ kt1l = 0.0
+ prwb = 0.0
+ pub1 = -2.1229706e-32
+ prwg = 0.0
+ puc1 = -9.461855e-24
+ la0 = 1.6783336e-7
+ eta0 = -0.00046875
+ pvag = 0.0
+ jsw = 1.2e-12
+ etab = 0.0006718753
+ kt1 = -0.2211471
+ lk1 = -8.844278e-9
+ kt2 = -0.014824204
+ lk2 = 3.718209e-9
+ vsat = 130812.46
+ )

.model pch_sf_13 pmos (
+ level = 49
+ wketa = -6.403492e-9
+ pvth0 = 1.18629e-15
+ drout = 0.0
+ toxm = 4.08e-9
+ tpbsw = 0.001572025
+ pbsw = 0.895226
+ pclm = 0.5999999
+ cjswg = 4.00995e-10
+ mjswg = 0.3683619
+ wvoff = -1.320298e-9
+ weta0 = 0
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ wvsat = 0.0
+ keta = 0.04310941
+ pscbe1 = 199999970.0
+ pscbe2 = 5e-7
+ wvth0 = 1.0526903e-8
+ dsub = 0.0
+ nqsmod = 0
+ tpbswg = 0.001572025
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ noimod = 2
+ voff = -0.1261533
+ ldif = 9e-8
+ a0 = 0.8704194
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ at = 10000.0
+ cf = 0
+ cj = 0.00106495
+ ef = 1.064
+ k1 = 0.5421249
+ k2 = 0.0301404
+ k3 = 0.0
+ em = 30000000.0
+ ags = 0.02
+ eta0 = 5e-5
+ js = 2.5e-7
+ ll = 0.0
+ mj = 0.4476
+ lw = 0.0
+ pvag = 0.0
+ etab = -5e-5
+ u0 = 0.009803694200000001
+ pb = 0.895226
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ vsat = 149999.98
+ xpart = 1
+ ua = 1.2584637e-9
+ ub = 4.999999e-20
+ uc = -1.6065008e-10
+ wint = 5e-9
+ wl = 0.0
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ cit = -0.0001
+ vth0 = -0.4247409
+ rdsw = 530.0
+ dlc = 2e-9
+ wkt1 = 3.830554e-9
+ wkt2 = 1.9527771e-9
+ k3b = 0.0
+ lint = 1.4999999e-8
+ pbswg = 0.895226
+ dwb = 0.0
+ wmax = 5e-7
+ dwg = 0.0
+ nfactor = 1.0
+ wmin = 2.2e-7
+ lvoff = 1.5817200000000002e-9
+ lmax = 2.0001e-5
+ lmin = 1e-5
+ capmod = 3
+ beta0 = 22.67827
+ leta0 = 4.745160018966694e-10
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.001
+ pdiblcb = 0.01
+ jsw = 1.2e-12
+ kt1 = -0.2247607
+ kt2 = -0.027069092
+ lk2 = -1.18629e-9
+ lvth0 = 3.9543e-9
+ llc = -0.039
+ lln = -1
+ lu0 = 7.9086e-11
+ wub1 = 2.1644123e-27
+ wuc1 = -1.2526765e-17
+ nch = 3.9e+17
+ mobmod = 1
+ lwl = 0.0
+ lwn = 1.0
+ delta = 0.01
+ hdif = 2e-7
+ nlx = 0.0
+ pnfactor = 0
+ binunit = 2
+ wute = 6.898109e-9
+ mjsw = 0.3683619
+ wnfactor = 0.0
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ pu0 = 0.0
+ prt = 0
+ rsh = 7.2
+ tcj = 0.0009739001
+ ua1 = 1.224e-9
+ ub1 = -1.3041941e-18
+ uc1 = 6.665171e-11
+ cdsc = 0.0
+ tpb = 0.001572025
+ tox = 4.08e-9
+ wa0 = 8.951166e-8
+ lnfactor = 3.9543e-9
+ cgdo = 3.28e-10
+ ute = -0.7678431
+ wk1 = 3.561511e-9
+ wk2 = -4.719829e-9
+ wln = 1.0
+ cgso = 3.28e-10
+ wu0 = -2.057536e-11
+ wua = -2.3131395e-16
+ wuc = -1.2695932e-17
+ wwl = 0.0
+ wwn = 1.0
+ xti = 3
+ tcjsw = 0.0004130718
+ tcjswg = 0.0004130718
+ version = 3.24
+ cjsw = 2.35695e-10
+ pvoff = 0.0
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 4.7451600189666944e-17
+ tnom = 25.0
+ )

.model pch_sf_14 pmos (
+ level = 49
+ tpbswg = 0.001572025
+ noimod = 2
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0004772729
+ cit = -0.0001
+ wub1 = -3.0198158e-27
+ wuc1 = -1.0513175e-17
+ pdiblcb = 0.01
+ lpscbe1 = 195.04262
+ dlc = 2e-9
+ hdif = 2e-7
+ k3b = 0.0
+ lub1 = -2.0820251e-25
+ dwb = 0.0
+ dwg = 0.0
+ luc1 = 9.921307e-17
+ wute = 1.1298283e-8
+ mjsw = 0.3683619
+ binunit = 2
+ lketa = -4.562476e-8
+ lute = 2.2927659e-7
+ xpart = 1
+ la0 = 5.081137e-7
+ cdsc = 0.0
+ jsw = 1.2e-12
+ kt1 = -0.2237138
+ lk1 = -4.88067e-8
+ kt2 = -0.026908273
+ lk2 = 2.2115907999999998e-8
+ llc = -0.039
+ lln = -1
+ cgdo = 3.28e-10
+ lu0 = -2.2091919e-10
+ pbswg = 0.895226
+ lua = -3.24011e-17
+ lub = -3.941427e-28
+ luc = -6.882293e-17
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ cgso = 3.28e-10
+ pa0 = -1.854315e-13
+ lvoff = -8.068828999999997e-10
+ nlx = 0.0
+ capmod = 3
+ pk1 = 3.786126e-14
+ pk2 = -1.6169635e-14
+ beta0 = 22.67827
+ pu0 = -6.225135e-16
+ leta0 = 4.745160018966694e-10
+ prt = 0
+ pua = -1.3939852e-23
+ pub = 1.1764949e-34
+ puc = 1.4094153e-23
+ cjsw = 2.35695e-10
+ lvsat = -0.013002842
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ lvth0 = -6.54035e-10
+ version = 3.24
+ rsh = 7.2
+ tcj = 0.0009739001
+ mobmod = 1
+ ua1 = 1.224e-9
+ ub1 = -1.2832692e-18
+ uc1 = 5.668055e-11
+ tpb = 0.001572025
+ tox = 4.08e-9
+ delta = 0.01
+ wa0 = 1.0814799e-7
+ tnom = 25.0
+ ute = -0.790886
+ wk1 = -2.4364055e-10
+ wk2 = -3.0947396e-9
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ wln = 1.0
+ wu0 = 4.1988812999999995e-11
+ toxm = 4.08e-9
+ wua = -2.2991296e-16
+ wub = -1.1822094e-29
+ wuc = -1.4112429e-17
+ wwl = 0.0
+ wwn = 1.0
+ pbsw = 0.895226
+ xti = 3
+ pclm = 0.5738635
+ pketa = 1.7549415e-14
+ a0 = 0.8193527
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ at = 10000.0
+ cf = 0
+ cj = 0.00106495
+ ef = 1.064
+ k1 = 0.5470301
+ k2 = 0.027798470000000002
+ k3 = 0.0
+ em = 30000000.0
+ js = 2.5e-7
+ ll = 0.0
+ mj = 0.4476
+ lw = 0.0
+ u0 = 0.0098338462
+ pb = 0.895226
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ua = 1.2617201e-9
+ ub = 5.00396e-20
+ uc = -1.5373321e-10
+ wl = 0.0
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -2e-8
+ ww = 0.0
+ tcjswg = 0.0004130718
+ xw = 0.0
+ tcjsw = 0.0004130718
+ pkt1 = 2.5501714e-15
+ pkt2 = -4.817884e-16
+ keta = 0.04769481
+ pvoff = 2.6840621e-15
+ dsub = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 4.7451600189666944e-17
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ pnfactor = 0
+ wketa = -8.167253e-9
+ pvth0 = -2.454092e-15
+ wnfactor = 0.0
+ voff = -0.1259132
+ drout = 0.0
+ ldif = 9e-8
+ tpbsw = 0.001572025
+ kt1l = 0.0
+ prwb = 0.0
+ pub1 = 5.158311e-32
+ prwg = 0.0
+ puc1 = -2.0035212e-23
+ eta0 = 5e-5
+ cjswg = 4.00995e-10
+ pvag = 0.0
+ etab = -5e-5
+ vsat = 151306.8
+ mjswg = 0.3683619
+ wint = 5e-9
+ pute = -4.378173e-14
+ vth0 = -0.4242777
+ rdsw = 530.0
+ lnfactor = 3.9543e-9
+ wvoff = -1.590053e-9
+ wkt1 = 3.574256e-9
+ wkt2 = 2.0011981e-9
+ lint = 1.4999999e-8
+ wmax = 5e-7
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ wmin = 2.2e-7
+ lkt1 = -1.0417262e-8
+ lkt2 = -1.6001408e-9
+ weta0 = 0
+ nfactor = 1.0
+ lmax = 1e-5
+ pscbe1 = 180397700.0
+ pscbe2 = 5e-7
+ wvsat = 0.0
+ lmin = 1.2e-6
+ lpclm = 2.6005691e-7
+ wvth0 = 1.089277e-8
+ lpdiblc2 = 5.201136e-9
+ ags = 0.02
+ nqsmod = 0
+ )

.model pch_sf_15 pmos (
+ level = 49
+ ute = -0.5904401
+ wk1 = 4.182789e-8
+ wk2 = -2.2085489e-8
+ beta0 = 22.67827
+ wln = 1.0
+ wu0 = -3.789626e-10
+ pkt1 = -8.599671e-15
+ pkt2 = 1.9347028e-16
+ lpdiblc2 = 3.696429e-9
+ keta = 0.0004484208
+ wua = -1.9008923e-16
+ leta0 = 5.114802818966694e-10
+ wub = 8.369847e-27
+ wuc = 5.370726e-18
+ wwl = 0.0
+ wwn = 1.0
+ letab = -3.696428e-11
+ xti = 3
+ mobmod = 1
+ lvsat = -0.007392816
+ dsub = 0.0
+ lvth0 = -1.1578233000000001e-8
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ delta = 0.01
+ lcit = 2.2622144e-10
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ voff = -0.1186655
+ ldif = 9e-8
+ kt1l = 0.0
+ prwb = 0.0
+ pub1 = -1.2589071e-33
+ prwg = 0.0
+ puc1 = 4.27717e-24
+ eta0 = 1.7857146e-5
+ pvag = 0.0
+ etab = -1.7857146e-5
+ vsat = 146428.52
+ wint = 5e-9
+ pute = -8.783067e-15
+ vth0 = -0.4147784
+ rdsw = 530.0
+ pketa = -5.090041e-15
+ wkt1 = 1.3269771e-8
+ wkt2 = 1.4140165e-9
+ lint = 1.4999999e-8
+ wmax = 5e-7
+ tcjswg = 0.0004130718
+ wmin = 2.2e-7
+ lkt1 = 1.1386779e-8
+ lkt2 = -8.841858e-10
+ lmax = 1.2e-6
+ lmin = 5e-7
+ tcjsw = 0.0004130718
+ nfactor = 1.0
+ pvoff = 3.95383e-15
+ wub1 = 4.292976e-26
+ cdscb = 0.0
+ wuc1 = -3.165437e-17
+ cdscd = 0.0
+ peta0 = 4.7451600189666944e-17
+ hdif = 2e-7
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0017857139
+ pdiblcb = 0.01
+ lub1 = -9.299159e-27
+ wketa = 1.1519229e-8
+ luc1 = 4.434689e-18
+ pvth0 = 1.9485986e-15
+ wute = -1.9135335e-8
+ mjsw = 0.3683619
+ drout = 0.0
+ tpbsw = 0.001572025
+ lute = -1.2362289e-9
+ cjswg = 4.00995e-10
+ binunit = 2
+ mjswg = 0.3683619
+ ags = 0.02
+ cdsc = 0.0
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ wvoff = -2.6941984e-9
+ cit = -0.00029671428
+ cgdo = 3.28e-10
+ pscbe1 = 349999900.0
+ pscbe2 = 5e-7
+ dlc = 2e-9
+ cgso = 3.28e-10
+ k3b = 0.0
+ weta0 = 0
+ dwb = 0.0
+ dwg = 0.0
+ wvsat = 0.0
+ lpclm = 1.4785714e-7
+ wvth0 = 7.064344e-9
+ nqsmod = 0
+ a0 = 1.1508681
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ tpbswg = 0.001572025
+ cjsw = 2.35695e-10
+ noimod = 2
+ at = 10000.0
+ cf = 0
+ cj = 0.00106495
+ ef = 1.064
+ k1 = 0.510219
+ k2 = 0.04857026
+ k3 = 0.0
+ em = 30000000.0
+ js = 2.5e-7
+ ll = 0.0
+ noia = 9.5e+18
+ mj = 0.4476
+ noib = 100000.0
+ noic = 1.4e-12
+ lw = 0.0
+ u0 = 0.0092586472
+ pb = 0.895226
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ua = 1.0922192e-9
+ ub = 2.0536515e-20
+ uc = -2.183638e-10
+ la0 = 1.2687106e-7
+ wl = 0.0
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ jsw = 1.2e-12
+ version = 3.24
+ kt1 = -0.2426738
+ lk1 = -6.473878e-9
+ kt2 = -0.027530843
+ lk2 = -1.7716528e-9
+ llc = -0.039
+ lln = -1
+ pnfactor = 0
+ lu0 = 4.405597e-10
+ tnom = 25.0
+ lua = 1.6252487e-16
+ lub = 3.353441e-26
+ luc = 5.502275e-18
+ nch = 3.9e+17
+ wnfactor = 0.0
+ lwl = 0.0
+ lwn = 1.0
+ pa0 = 5.971399e-14
+ nlx = 0.0
+ toxm = 4.08e-9
+ lketa = 8.708591e-9
+ pk1 = -1.0521005e-14
+ pk2 = 5.669729e-15
+ pbsw = 0.895226
+ pclm = 0.6714286
+ pu0 = -1.384194e-16
+ xpart = 1
+ prt = 0
+ pua = -5.973716e-23
+ pub = -9.521269e-33
+ puc = -8.311478e-24
+ rsh = 7.2
+ lnfactor = 3.9543e-9
+ tcj = 0.0009739001
+ ua1 = 1.224e-9
+ ub1 = -1.4562286e-18
+ uc1 = 1.3909653e-10
+ pbswg = 0.895226
+ capmod = 3
+ tpb = 0.001572025
+ tox = 4.08e-9
+ wa0 = -1.0502199e-7
+ lvoff = -9.141699e-9
+ )

.model pch_sf_16 pmos (
+ level = 49
+ cdsc = 0.0
+ binunit = 2
+ pketa = 7.45672e-16
+ lnfactor = 3.9543e-9
+ tcjswg = 0.0004130718
+ cgdo = 3.28e-10
+ wpclm = 4.634222e-9
+ cgso = 3.28e-10
+ tcjsw = 0.0004130718
+ lpdiblc2 = 1.8281252e-9
+ cjsw = 2.35695e-10
+ pvoff = 1.4541431e-15
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ wcdscd = -1.4183201e-11
+ ags = 0.03625
+ cdscb = 0.0
+ cdscd = -6.449223e-5
+ peta0 = 4.7451600189666944e-17
+ cit = 8.534377e-5
+ tnom = 25.0
+ wketa = -1.4490222e-9
+ pvth0 = 9.0214192e-16
+ version = 3.24
+ dlc = 2e-9
+ drout = 0.0
+ pcdscd = 6.382441e-18
+ tpbsw = 0.001572025
+ k3b = 0.0
+ toxm = 4.08e-9
+ dwb = 0.0
+ dwg = 0.0
+ pbsw = 0.895226
+ pclm = 0.9648299
+ cjswg = 4.00995e-10
+ mjswg = 0.3683619
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ wvoff = 2.8606606e-9
+ pscbe1 = 350000000.0
+ pscbe2 = 5e-7
+ la0 = 7.233052e-9
+ jsw = 1.2e-12
+ kt1 = -0.2130934
+ lk1 = 1.3789155e-8
+ kt2 = -0.03589084
+ lk2 = -4.293236e-9
+ llc = -0.039
+ weta0 = 0
+ lln = -1
+ lu0 = -2.775402e-10
+ nqsmod = 0
+ lua = -2.6402067e-16
+ lub = 2.6345733e-25
+ luc = 3.340897e-17
+ nch = 3.9e+17
+ wvsat = 0.0
+ tpbswg = 0.001572025
+ lwl = 0.0
+ lwn = 1.0
+ noimod = 2
+ lpclm = 1.5826547e-8
+ pa0 = -6.072043e-15
+ wvth0 = 9.389803e-9
+ nlx = 0.0
+ pkt1 = -9.758805e-16
+ pkt2 = -1.0643102e-15
+ keta = 0.03159368
+ pk1 = 4.122718e-15
+ pk2 = -2.3103772e-15
+ dsub = 0.0
+ pu0 = 1.3574996e-16
+ prt = 0
+ pua = 6.304761e-23
+ pub = -7.522618e-32
+ puc = -8.758834e-24
+ lags = -7.312499e-9
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ rsh = 7.2
+ tcj = 0.0009739001
+ ua1 = 1.224e-9
+ ub1 = -1.4433942e-18
+ uc1 = 2.0396977e-10
+ tpb = 0.001572025
+ tox = 4.08e-9
+ lcit = 5.429531e-11
+ voff = -0.1287204
+ wa0 = 4.116919e-8
+ lcdscd = 2.9021494e-11
+ ldif = 9e-8
+ ute = -0.5893072
+ wk1 = 9.286284e-9
+ kt1l = 0.0
+ wk2 = -4.351921e-9
+ prwb = 0.0
+ pub1 = 1.9106841e-32
+ prwg = 0.0
+ lketa = -5.306775e-9
+ puc1 = 6.153712e-24
+ wln = 1.0
+ wu0 = -9.882279e-10
+ eta0 = -0.0004687502
+ wua = -4.629443e-16
+ pvag = 0.0
+ wub = 1.5438073e-25
+ wuc = 6.364847e-18
+ etab = 0.0006718753
+ xpart = 1
+ wwl = 0.0
+ wwn = 1.0
+ vsat = 130812.55
+ xti = 3
+ wint = 5e-9
+ pute = 5.968411e-15
+ vth0 = -0.4276605
+ capmod = 3
+ rdsw = 530.0
+ wkt1 = -3.671987e-9
+ wkt2 = 4.209085e-9
+ pbswg = 0.895226
+ lint = 1.4999999e-8
+ wmax = 5e-7
+ wmin = 2.2e-7
+ lvoff = -4.616999000000001e-9
+ lkt1 = -1.9244071e-9
+ lkt2 = 2.877812e-9
+ lmax = 5e-7
+ beta0 = 22.67827
+ lmin = 1.8e-7
+ mobmod = 1
+ leta0 = 7.304535818966694e-10
+ letab = -3.473438e-10
+ lvsat = -0.0003656336
+ nfactor = 1.0
+ lvth0 = -5.781281000000001e-9
+ ppclm = -2.0853998e-15
+ wub1 = -2.3274574e-27
+ wuc1 = -3.582447e-17
+ delta = 0.01
+ hdif = 2e-7
+ a0 = 1.4167303
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ pnfactor = 0
+ lub1 = -1.5074642e-26
+ luc1 = -2.4758267e-17
+ at = 10000.0
+ cf = 0
+ cj = 0.00106495
+ ef = 1.064
+ k1 = 0.46519
+ dvt0w = 0.0
+ k2 = 0.05417378
+ k3 = 0.0
+ em = 30000000.0
+ wnfactor = 0.0
+ wute = -5.191639e-8
+ dvt1w = 0.0
+ dvt2w = 0.0
+ mjsw = 0.3683619
+ js = 2.5e-7
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.005937499
+ ll = 0.0
+ mj = 0.4476
+ lw = 0.0
+ u0 = 0.0108544242
+ pb = 0.895226
+ w0 = 0.0
+ rd = 0
+ pdiblcb = 0.01
+ rs = 0
+ ua = 2.0400983e-9
+ ub = -4.904033e-19
+ uc = -2.8037866e-10
+ wl = 0.0
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -2e-8
+ ww = 0.0
+ lute = -1.7460413e-9
+ xw = 0.0
+ )

.model pch_mc_1 pmos (
+ level = 49
+ lvth0 = 0.0
+ cdsc = 0.0
+ binunit = 2
+ pnfactor = 0
+ cgdo = 3.28e-10
+ delta = 0.01
+ wnfactor = 0.0
+ cgso = 3.28e-10
+ dvt0w = 0.0
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ dvt1w = 0.0
+ dvt2w = 0.0
+ pscbe1 = 199999970.0
+ pscbe2 = 5e-7
+ cjsw = 2.481e-10
+ ags = 0.02
+ lnfactor = 0.0
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ nqsmod = 0
+ tpbswg = 0.001572025
+ noimod = 2
+ cit = -0.0001
+ dlc = 2e-9
+ tnom = 25.0
+ version = 3.24
+ k3b = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ toxm = 4.08e-9
+ tcjsw = 0.0004130718
+ pbsw = 0.895226
+ pclm = 0.6000001
+ pvoff = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ jsw = 1.2e-12
+ peta0 = 5.5000000000000005e-21
+ kt1 = -0.2311294
+ lk2 = 0.0
+ kt2 = -0.02433992
+ llc = -0.039
+ lln = -1
+ lu0 = 0.0
+ nch = 3.9e+17
+ pvth0 = 0.0
+ lwl = 0.0
+ lwn = 1.0
+ drout = 0.0
+ nlx = 0.0
+ tpbsw = 0.001572025
+ capmod = 3
+ keta = 0.026632193
+ pu0 = 0.0
+ cjswg = 4.221e-10
+ prt = 0
+ dsub = 0.0
+ mjswg = 0.3683619
+ rsh = 7.2
+ tcj = 0.0009739001
+ ua1 = 1.224e-9
+ ub1 = -1.3928839e-18
+ uc1 = -4.59467e-12
+ wvoff = 0.0
+ mobmod = 1
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ tpb = 0.001572025
+ tox = 4.08e-9
+ ute = -0.8288856
+ voff = -0.1275921
+ weta0 = 0
+ ldif = 9e-8
+ wvsat = 0.0
+ wln = 1.0
+ kt1l = 0.0
+ prwb = 0.0
+ wu0 = 0.0
+ prwg = 0.0
+ wvth0 = 0.0
+ wwl = 0.0
+ wwn = 1.0
+ eta0 = 5e-5
+ xti = 3
+ pvag = 0.0
+ etab = -5e-5
+ vsat = 149999.98
+ wint = 5e-9
+ vth0 = -0.4384811
+ rdsw = 530.0
+ lint = 1.4999999e-8
+ wmax = 0.000900001
+ wmin = 1e-5
+ a0 = 1.0461572
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ lmax = 2.0001e-5
+ at = 10000.0
+ cf = 0
+ cj = 0.001121
+ lmin = 1e-5
+ ef = 1.064
+ k1 = 0.5375325
+ k2 = 0.03503256
+ k3 = 0.0
+ em = 30000000.0
+ tcjswg = 0.0004130718
+ js = 2.5e-7
+ ll = 0.0
+ mj = 0.4476
+ lw = 0.0
+ u0 = 0.010865118
+ pb = 0.895226
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ua = 8.23294e-10
+ ub = 6.854322e-19
+ uc = -8.655411e-11
+ wl = 0.0
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ xpart = 1
+ nfactor = 1.0
+ pbswg = 0.895226
+ hdif = 2e-7
+ lvoff = 0.0
+ mjsw = 0.3683619
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0010000003
+ pdiblcb = 0.01
+ beta0 = 22.67827
+ leta0 = 8e-15
+ )

.model pch_mc_2 pmos (
+ level = 49
+ mj = 0.4476
+ lw = 0.0
+ kt1 = -0.2295883
+ lk1 = 1.8783622e-8
+ kt2 = -0.024031118
+ lk2 = -5.487172e-9
+ u0 = 0.010995165
+ pb = 0.895226
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ua = 8.625313e-10
+ ub = 6.401998e-19
+ uc = -8.855145e-11
+ llc = -0.039
+ lln = -1
+ wl = 0.0
+ lu0 = -1.2939689e-9
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ voff = -0.1274002
+ lua = -3.904111e-16
+ lub = 4.500626e-25
+ luc = 1.9873557e-17
+ ldif = 9e-8
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ kt1l = 0.0
+ tcjsw = 0.0004130718
+ prwb = 0.0
+ prwg = 0.0
+ nlx = 0.0
+ eta0 = 5e-5
+ pvag = 0.0
+ etab = -5e-5
+ pvoff = 0.0
+ vsat = 151306.8
+ pu0 = 0.0
+ wint = 5e-9
+ prt = 0
+ vth0 = -0.4359872
+ rdsw = 530.0
+ pnfactor = 0
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 5.5000000000000005e-21
+ lint = 1.4999999e-8
+ rsh = 7.2
+ tcj = 0.0009739001
+ ua1 = 1.224e-9
+ wnfactor = 0.0
+ wmax = 0.000900001
+ ub1 = -1.3977103e-18
+ uc1 = -6.694918e-12
+ wmin = 1e-5
+ tpb = 0.001572025
+ capmod = 3
+ pvth0 = 0.0
+ tox = 4.08e-9
+ lkt1 = -1.5333228e-8
+ lkt2 = -3.0725886e-9
+ drout = 0.0
+ lmax = 1e-5
+ tpbsw = 0.001572025
+ ute = -0.8385549
+ lmin = 1.2e-6
+ wln = 1.0
+ wu0 = 0.0
+ cjswg = 4.221e-10
+ wwl = 0.0
+ wwn = 1.0
+ mjswg = 0.3683619
+ lnfactor = 0.0
+ xti = 3
+ mobmod = 1
+ nfactor = 1.0
+ wvoff = 0.0
+ hdif = 2e-7
+ lub1 = 4.802326e-26
+ luc1 = 2.0897466e-17
+ weta0 = 0
+ mjsw = 0.3683619
+ lpdiblc2 = 5.201137e-9
+ wvsat = 0.0
+ lute = 9.620972e-8
+ lpclm = 2.6005682e-7
+ wvth0 = 0.0
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0004772727
+ pdiblcb = 0.01
+ lpscbe1 = 195.04263
+ cdsc = 0.0
+ cgdo = 3.28e-10
+ binunit = 2
+ cgso = 3.28e-10
+ tcjswg = 0.0004130718
+ lketa = -2.0462676e-9
+ cjsw = 2.481e-10
+ xpart = 1
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ pbswg = 0.895226
+ tnom = 25.0
+ lvoff = -1.9091309e-9
+ toxm = 4.08e-9
+ beta0 = 22.67827
+ version = 3.24
+ pbsw = 0.895226
+ pclm = 0.5738637
+ leta0 = 8e-15
+ lvsat = -0.013002843
+ lvth0 = -2.4814053e-8
+ ags = 0.02
+ delta = 0.01
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ cit = -0.0001
+ dlc = 2e-9
+ dvt0w = 0.0
+ dvt1w = 0.0
+ pscbe1 = 180397680.0
+ pscbe2 = 5e-7
+ dvt2w = 0.0
+ k3b = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ keta = 0.026837848
+ nqsmod = 0
+ tpbswg = 0.001572025
+ dsub = 0.0
+ noimod = 2
+ a0 = 1.0385712
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ at = 10000.0
+ cf = 0
+ cj = 0.001121
+ la0 = 7.548124e-8
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ ef = 1.064
+ k1 = 0.5356447
+ k2 = 0.03558403
+ k3 = 0.0
+ em = 30000000.0
+ js = 2.5e-7
+ jsw = 1.2e-12
+ ll = 0.0
+ )

.model pch_mc_3 pmos (
+ level = 49
+ cjswg = 4.221e-10
+ mjswg = 0.3683619
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ wvoff = 0.0
+ tnom = 25.0
+ weta0 = 0
+ wvsat = 0.0
+ toxm = 4.08e-9
+ a0 = 1.0045335
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ lpclm = 1.4785704e-7
+ wvth0 = 0.0
+ pbsw = 0.895226
+ pclm = 0.6714287
+ at = 10000.0
+ cf = 0
+ cj = 0.001121
+ ef = 1.064
+ k1 = 0.5405614
+ k2 = 0.03490157
+ k3 = 0.0
+ em = 30000000.0
+ js = 2.5e-7
+ version = 3.24
+ ll = 0.0
+ mj = 0.4476
+ lw = 0.0
+ u0 = 0.010224584
+ pb = 0.895226
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ua = 5.26694e-10
+ ub = 1.1734415e-18
+ uc = -4.332115e-11
+ wl = 0.0
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ pnfactor = 0
+ wnfactor = 0.0
+ tcjswg = 0.0004130718
+ lketa = -8.158225e-9
+ keta = 0.03215259
+ xpart = 1
+ dsub = 0.0
+ lnfactor = 0.0
+ ags = 0.02
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ pbswg = 0.895226
+ lvoff = -9.487825e-10
+ lcit = 2.2402701e-10
+ cit = -0.00029480609
+ voff = -0.1282353
+ lpdiblc2 = 3.696428e-9
+ ldif = 9e-8
+ dlc = 2e-9
+ beta0 = 22.67827
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ k3b = 0.0
+ dwb = 0.0
+ leta0 = 3.697228e-11
+ dwg = 0.0
+ eta0 = 1.7857143e-5
+ letab = -3.696428e-11
+ pvag = 0.0
+ etab = -1.7857143e-5
+ lvsat = -0.007392833
+ vsat = 146428.53
+ wint = 5e-9
+ lvth0 = -6.689442e-9
+ vth0 = -0.4517478
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ rdsw = 530.0
+ delta = 0.01
+ lint = 1.4999999e-8
+ wmax = 0.000900001
+ pscbe1 = 349999900.0
+ pscbe2 = 5e-7
+ la0 = 1.146246e-7
+ wmin = 1e-5
+ jsw = 1.2e-12
+ lkt1 = 1.5747348e-9
+ lkt2 = 9.740028e-10
+ kt1 = -0.2442909
+ lk1 = 1.3129389e-8
+ kt2 = -0.027549893
+ lk2 = -4.702335e-9
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ lmax = 1.2e-6
+ llc = -0.039
+ lln = -1
+ lu0 = -4.078006e-10
+ lmin = 5e-7
+ lua = -4.198125e-18
+ lub = -1.631654e-25
+ luc = -3.214129e-17
+ nch = 3.9e+17
+ nqsmod = 0
+ lwl = 0.0
+ lwn = 1.0
+ tpbswg = 0.001572025
+ noimod = 2
+ nlx = 0.0
+ pu0 = 0.0
+ prt = 0
+ hdif = 2e-7
+ rsh = 7.2
+ tcj = 0.0009739001
+ nfactor = 1.0
+ ua1 = 1.224e-9
+ lub1 = 3.0810812e-26
+ ub1 = -1.3827429e-18
+ luc1 = 2.9752128e-17
+ uc1 = -1.4394627e-11
+ mjsw = 0.3683619
+ tpb = 0.001572025
+ tox = 4.08e-9
+ tcjsw = 0.0004130718
+ lute = 3.654092e-8
+ ute = -0.786669
+ wln = 1.0
+ pvoff = 0.0
+ wu0 = 0.0
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0017857148
+ wwl = 0.0
+ wwn = 1.0
+ pdiblcb = 0.01
+ cdsc = 0.0
+ xti = 3
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 5.5000000000000005e-21
+ capmod = 3
+ cgdo = 3.28e-10
+ pvth0 = 0.0
+ cgso = 3.28e-10
+ drout = 0.0
+ binunit = 2
+ tpbsw = 0.001572025
+ cjsw = 2.481e-10
+ mobmod = 1
+ )

.model pch_mc_4 pmos (
+ level = 49
+ wmin = 1e-5
+ lkt1 = -2.665e-9
+ lkt2 = -2.325577e-10
+ lmax = 5e-7
+ cit = -4.054396e-5
+ lmin = 1.8e-7
+ lketa = -8.307595e-10
+ dlc = 2e-9
+ k3b = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ xpart = 1
+ pbswg = 0.895226
+ hdif = 2e-7
+ lub1 = 2.883988e-26
+ luc1 = -6.846759e-18
+ lvoff = -3.571592e-11
+ la0 = 1.6196543e-8
+ mjsw = 0.3683619
+ jsw = 1.2e-12
+ kt1 = -0.2348693
+ lk1 = 1.6807924e-8
+ kt2 = -0.024868647
+ lk2 = -5.876215e-9
+ beta0 = 22.67827
+ nfactor = 1.0
+ llc = -0.039
+ lln = -1
+ lu0 = -9.894781e-11
+ lute = 1.6013461e-9
+ leta0 = 2.5594552000000003e-10
+ lua = -1.5999061e-16
+ lub = 1.2197973e-25
+ luc = 1.8500639e-17
+ nch = 3.9e+17
+ letab = -5.298917e-10
+ lwl = 0.0
+ lwn = 1.0
+ lvsat = -0.0003656265
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ nlx = 0.0
+ lvth0 = -8.240552e-9
+ cdsc = 0.0
+ pscbe1 = 350000000.0
+ pscbe2 = 5e-7
+ pnfactor = 0
+ pu0 = 0.0
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.00796875
+ delta = 0.01
+ a0 = 1.2232625
+ a1 = 0.0
+ a2 = 0.4
+ prt = 0
+ b0 = 0.0
+ b1 = 0.0
+ cgdo = 3.28e-10
+ wnfactor = 0.0
+ pdiblcb = 0.01
+ at = 10000.0
+ cf = 0
+ cj = 0.001121
+ ef = 1.064
+ k1 = 0.5323869
+ k2 = 0.03751019
+ k3 = 0.0
+ em = 30000000.0
+ cgso = 3.28e-10
+ js = 2.5e-7
+ dvt0w = 0.0
+ dvt1w = 0.0
+ ll = 0.0
+ rsh = 7.2
+ mj = 0.4476
+ dvt2w = 0.0
+ lw = 0.0
+ u0 = 0.009538244
+ tcj = 0.0009739001
+ nqsmod = 0
+ pb = 0.895226
+ ua1 = 1.224e-9
+ w0 = 0.0
+ ub1 = -1.3783631e-18
+ rd = 0
+ uc1 = 6.693623e-11
+ tpbswg = 0.001572025
+ rs = 0
+ ua = 8.728995e-10
+ ub = 5.397856e-19
+ uc = -1.5585878e-10
+ noimod = 2
+ wl = 0.0
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ tpb = 0.001572025
+ tox = 4.08e-9
+ binunit = 2
+ cjsw = 2.481e-10
+ ute = -0.7090256
+ lnfactor = 0.0
+ wln = 1.0
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ wu0 = 0.0
+ wwl = 0.0
+ wwn = 1.0
+ xti = 3
+ tnom = 25.0
+ lcdscd = 3.65625e-11
+ lpdiblc2 = 9.140626e-10
+ toxm = 4.08e-9
+ tcjsw = 0.0004130718
+ pbsw = 0.895226
+ pclm = 0.9102259
+ pvoff = 0.0
+ capmod = 3
+ version = 3.24
+ cdscb = 0.0
+ cdscd = -8.125e-5
+ peta0 = 5.5000000000000005e-21
+ pvth0 = 0.0
+ drout = 0.0
+ tpbsw = 0.001572025
+ mobmod = 1
+ keta = 0.015869336
+ cjswg = 4.221e-10
+ mjswg = 0.3683619
+ dsub = 0.0
+ wvoff = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ weta0 = 0
+ lcit = 1.0960905e-10
+ voff = -0.1302643
+ ldif = 9e-8
+ wvsat = 0.0
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ lpclm = 4.03983e-8
+ wvth0 = 0.0
+ eta0 = -0.0004687502
+ pvag = 0.0
+ etab = 0.0010775371
+ vsat = 130812.52
+ wint = 5e-9
+ vth0 = -0.4483009
+ rdsw = 530.0
+ tcjswg = 0.0004130718
+ lint = 1.4999999e-8
+ wmax = 0.000900001
+ ags = 0.02
+ )

.model pch_mc_5 pmos (
+ level = 49
+ wa0 = -4.787191e-8
+ pscbe1 = 199999970.0
+ pscbe2 = 5e-7
+ ute = -0.8394966
+ lvth0 = 0.0
+ wk1 = 1.2456701e-8
+ wk2 = -5.940143e-9
+ wln = 1.0
+ wu0 = -1.2494747e-9
+ delta = 0.01
+ wua = 1.7543858e-16
+ wub = -6.530953e-25
+ wuc = -7.950096e-17
+ wwl = 0.0
+ wwn = 1.0
+ nqsmod = 0
+ xti = 3
+ version = 3.24
+ tpbswg = 0.001572025
+ noimod = 2
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ keta = 0.02600144
+ dsub = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ voff = -0.1274889
+ ldif = 9e-8
+ tcjsw = 0.0004130718
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ eta0 = 5e-5
+ pvoff = 0.0
+ capmod = 3
+ pvag = 0.0
+ etab = -5e-5
+ vsat = 149999.98
+ wint = 5e-9
+ vth0 = -0.4397694
+ cdscb = 0.0
+ rdsw = 530.0
+ cdscd = 0.0
+ pnfactor = 0
+ peta0 = 5.5000000000000005e-21
+ wkt1 = 8.228274e-9
+ wkt2 = 1.4868883e-9
+ lint = 1.4999999e-8
+ wnfactor = 0.0
+ wmax = 1e-5
+ wketa = 6.301227e-9
+ wmin = 1.2e-6
+ pvth0 = 0.0
+ mobmod = 1
+ drout = 0.0
+ tpbsw = 0.001572025
+ lmax = 2.0001e-5
+ lmin = 1e-5
+ cjswg = 4.221e-10
+ a0 = 1.0509492
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ at = 10000.0
+ mjswg = 0.3683619
+ cf = 0
+ cj = 0.001121
+ lnfactor = 0.0
+ ef = 1.064
+ k1 = 0.5362856
+ k2 = 0.03562717
+ k3 = 0.0
+ em = 30000000.0
+ js = 2.5e-7
+ ll = 0.0
+ mj = 0.4476
+ lw = 0.0
+ u0 = 0.010990191
+ pb = 0.895226
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ wvoff = -1.0305298e-9
+ ua = 8.057326e-10
+ ub = 7.508071e-19
+ uc = -7.859605e-11
+ wub1 = 6.909715e-26
+ wuc1 = 3.0354498e-17
+ wl = 0.0
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ hdif = 2e-7
+ weta0 = 0
+ ags = 0.02
+ wute = 1.0600407e-7
+ mjsw = 0.3683619
+ wvsat = 0.0
+ wvth0 = 1.2870458e-8
+ cit = -0.0001
+ dlc = 2e-9
+ nfactor = 1.0
+ k3b = 0.0
+ tcjswg = 0.0004130718
+ dwb = 0.0
+ dwg = 0.0
+ cdsc = 0.0
+ cgdo = 3.28e-10
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0010000004
+ cgso = 3.28e-10
+ pdiblcb = 0.01
+ jsw = 1.2e-12
+ kt1 = -0.231953
+ kt2 = -0.024488758
+ lk2 = 0.0
+ llc = -0.039
+ lln = -1
+ cjsw = 2.481e-10
+ lu0 = 0.0
+ xpart = 1
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ binunit = 2
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ nlx = 0.0
+ pbswg = 0.895226
+ pu0 = 0.0
+ prt = 0
+ tnom = 25.0
+ lvoff = 0.0
+ rsh = 7.2
+ beta0 = 22.67827
+ toxm = 4.08e-9
+ tcj = 0.0009739001
+ ua1 = 1.224e-9
+ ub1 = -1.3998005e-18
+ uc1 = -7.633158e-12
+ leta0 = 8e-15
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ pbsw = 0.895226
+ pclm = 0.6000001
+ tpb = 0.001572025
+ tox = 4.08e-9
+ )

.model pch_mc_6 pmos (
+ level = 49
+ lub1 = 5.442727e-26
+ luc1 = 1.8276951e-17
+ wute = 1.0644106e-7
+ mjsw = 0.3683619
+ tcjsw = 0.0004130718
+ capmod = 3
+ lute = 9.664497e-8
+ pvoff = -4.403278e-15
+ nfactor = 1.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 5.5000000000000005e-21
+ mobmod = 1
+ cgdo = 3.28e-10
+ wketa = 7.084359e-9
+ pvth0 = -5.336472e-15
+ cgso = 3.28e-10
+ drout = 0.0
+ tpbsw = 0.001572025
+ ags = 0.02
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0004772728
+ pdiblcb = 0.01
+ lpscbe1 = 195.04262
+ cjswg = 4.221e-10
+ cit = -0.0001
+ cjsw = 2.481e-10
+ mjswg = 0.3683619
+ dlc = 2e-9
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ k3b = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ wvoff = -5.879894e-10
+ binunit = 2
+ tnom = 25.0
+ weta0 = 0
+ wvsat = 0.0
+ toxm = 4.08e-9
+ lpclm = 2.6005682e-7
+ wvth0 = 1.3406786e-8
+ la0 = 6.878132e-8
+ pbsw = 0.895226
+ tcjswg = 0.0004130718
+ pclm = 0.5738637
+ jsw = 1.2e-12
+ kt1 = -0.2303147
+ lk1 = 1.8184398e-8
+ kt2 = -0.024155809
+ lk2 = -5.280635e-9
+ llc = -0.039
+ lln = -1
+ lu0 = -1.3055237e-9
+ lua = -3.935608e-16
+ lub = 4.219459e-25
+ luc = 1.8883157e-17
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ pnfactor = 0
+ pa0 = 6.693222e-14
+ nlx = 0.0
+ wnfactor = 0.0
+ pk1 = 5.986243e-15
+ pk2 = -2.063307e-15
+ pu0 = 1.1543239e-16
+ prt = 0
+ pua = 3.1465633e-23
+ pub = 2.8088595e-31
+ puc = 9.8941e-24
+ version = 3.24
+ lketa = -1.2662711e-9
+ rsh = 7.2
+ pkt1 = 9.666697e-15
+ tcj = 0.0009739001
+ pkt2 = 2.4000725e-15
+ ua1 = 1.224e-9
+ keta = 0.026128704
+ ub1 = -1.4052706e-18
+ uc1 = -9.470036e-12
+ xpart = 1
+ tpb = 0.001572025
+ lnfactor = 0.0
+ tox = 4.08e-9
+ dsub = 0.0
+ wa0 = -5.459876e-8
+ ute = -0.8492097
+ wk1 = 1.185507e-8
+ wk2 = -5.732776e-9
+ pbswg = 0.895226
+ wln = 1.0
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ wu0 = -1.261076e-9
+ wua = 1.7227619e-16
+ wub = -6.81325e-25
+ wuc = -8.049533e-17
+ wwl = 0.0
+ wwn = 1.0
+ a0 = 1.0440365
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ lvoff = -1.4683624e-9
+ xti = 3
+ at = 10000.0
+ cf = 0
+ lpdiblc2 = 5.201137e-9
+ cj = 0.001121
+ voff = -0.1273414
+ ef = 1.064
+ k1 = 0.534458
+ k2 = 0.03615789
+ k3 = 0.0
+ em = 30000000.0
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ ldif = 9e-8
+ beta0 = 22.67827
+ js = 2.5e-7
+ ll = 0.0
+ mj = 0.4476
+ lw = 0.0
+ u0 = 0.0111214
+ pb = 0.895226
+ kt1l = 0.0
+ w0 = 0.0
+ prwb = 0.0
+ rd = 0
+ pub1 = -6.397619e-32
+ prwg = 0.0
+ leta0 = 8e-15
+ puc1 = 2.6178952e-23
+ rs = 0
+ ua = 8.452865e-10
+ ub = 7.084005e-19
+ uc = -8.049386e-11
+ pscbe1 = 180397700.0
+ pscbe2 = 5e-7
+ wl = 0.0
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ eta0 = 5e-5
+ lvsat = -0.013002842
+ pvag = 0.0
+ etab = -5e-5
+ vsat = 151306.8
+ lvth0 = -2.4279869e-8
+ wint = 5e-9
+ pute = -4.348101e-15
+ vth0 = -0.4373293
+ nqsmod = 0
+ rdsw = 530.0
+ tpbswg = 0.001572025
+ delta = 0.01
+ wkt1 = 7.256747e-9
+ wkt2 = 1.245675e-9
+ noimod = 2
+ lint = 1.4999999e-8
+ wmax = 1e-5
+ wmin = 1.2e-6
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ lkt1 = -1.6300865e-8
+ lkt2 = -3.312836e-9
+ lmax = 1e-5
+ lmin = 1.2e-6
+ pketa = -7.792167e-15
+ wub1 = 7.552692e-26
+ wuc1 = 2.7723443e-17
+ hdif = 2e-7
+ )

.model pch_mc_7 pmos (
+ level = 49
+ mjswg = 0.3683619
+ jsw = 1.2e-12
+ kt1 = -0.2459144
+ lk1 = 8.371453e-9
+ kt2 = -0.027846618
+ lk2 = -3.215854e-9
+ dsub = 0.0
+ llc = -0.039
+ lln = -1
+ lu0 = -3.457226e-10
+ wvoff = -7.866491e-9
+ lua = 3.0792715e-17
+ lub = -1.9665828e-25
+ luc = -3.700045e-17
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ wcit = -1.788104e-11
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ pa0 = -1.2519753e-13
+ nlx = 0.0
+ weta0 = 0
+ pk1 = 4.753178e-14
+ pk2 = -1.4849934e-14
+ lcit = 2.2196864e-10
+ voff = -0.1274479
+ pu0 = -6.201592e-16
+ wvsat = 0.0
+ ldif = 9e-8
+ tcjswg = 0.0004130718
+ prt = 0
+ pua = -3.495584e-22
+ pub = 3.345938e-31
+ puc = 4.854297e-23
+ lpclm = 1.4785702e-7
+ wvth0 = 1.013071e-8
+ kt1l = 0.0
+ prwb = 0.0
+ pub1 = -1.382964e-31
+ prwg = 0.0
+ puc1 = -5.043768e-23
+ eta0 = 1.7857139e-5
+ rsh = 7.2
+ tcj = 0.0009739001
+ ua1 = 1.224e-9
+ pvag = 0.0
+ ub1 = -1.3967723e-18
+ etab = -1.7857139e-5
+ uc1 = -2.3838735e-11
+ vsat = 146428.53
+ wint = 5e-9
+ pute = 2.0900147e-14
+ tpb = 0.001572025
+ tox = 4.08e-9
+ vth0 = -0.4527619
+ wa0 = 1.1247056e-7
+ rdsw = 530.0
+ ute = -0.7951261
+ wkt1 = 1.6218328e-8
+ wkt2 = 2.9642964e-9
+ wk1 = -2.4271484e-8
+ wk2 = 5.386031e-9
+ lint = 1.4999999e-8
+ wmax = 1e-5
+ wln = 1.0
+ wu0 = -6.214311e-10
+ wmin = 1.2e-6
+ wua = 5.036014e-16
+ wub = -7.280275e-25
+ wuc = -1.1410304e-16
+ lkt1 = 1.6387112e-9
+ lkt2 = 9.315946e-10
+ wwl = 0.0
+ wwn = 1.0
+ xti = 3
+ lmax = 1.2e-6
+ lketa = -8.380984e-9
+ lmin = 5e-7
+ xpart = 1
+ wub1 = 1.4015321e-25
+ pbswg = 0.895226
+ wuc1 = 9.434661e-17
+ hdif = 2e-7
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ lvoff = -1.3458795e-9
+ lub1 = 4.46543e-26
+ luc1 = 3.480094e-17
+ wute = 8.448607e-8
+ mjsw = 0.3683619
+ pscbe1 = 349999900.0
+ pscbe2 = 5e-7
+ beta0 = 22.67827
+ leta0 = 3.697229e-11
+ lute = 3.444881e-8
+ letab = -3.696429e-11
+ lvsat = -0.007392833
+ lvth0 = -6.532387e-9
+ nqsmod = 0
+ tpbswg = 0.001572025
+ noimod = 2
+ cdsc = 0.0
+ pnfactor = 0
+ delta = 0.01
+ wnfactor = 0.0
+ cgdo = 3.28e-10
+ nfactor = 1.0
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ cgso = 3.28e-10
+ cjsw = 2.481e-10
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0017857144
+ lnfactor = 0.0
+ pdiblcb = 0.01
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ pketa = 2.2253538e-15
+ tnom = 25.0
+ binunit = 2
+ capmod = 3
+ lpdiblc2 = 3.696428e-9
+ tcjsw = 0.0004130718
+ toxm = 4.08e-9
+ ags = 0.02
+ pcit = 2.0563189e-17
+ pbsw = 0.895226
+ pclm = 0.6714287
+ pvoff = 3.966999e-15
+ cit = -0.0002930162
+ a0 = 0.9932752
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ at = 10000.0
+ mobmod = 1
+ cf = 0
+ dlc = 2e-9
+ cj = 0.001121
+ ef = 1.064
+ k1 = 0.542991
+ k2 = 0.03436242
+ k3 = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ em = 30000000.0
+ peta0 = 5.5000000000000005e-21
+ k3b = 0.0
+ js = 2.5e-7
+ ll = 0.0
+ mj = 0.4476
+ lw = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ u0 = 0.010286789
+ pb = 0.895226
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ua = 4.762835e-10
+ ub = 1.2463172e-18
+ uc = -3.189942e-11
+ wl = 0.0
+ wr = 1.0
+ xj = 1.7000001e-7
+ wketa = -1.6265284e-9
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ pvth0 = -1.5689828e-15
+ drout = 0.0
+ tpbsw = 0.001572025
+ pkt1 = -6.391237e-16
+ pkt2 = 4.236579e-16
+ keta = 0.03231541
+ cjswg = 4.221e-10
+ version = 3.24
+ la0 = 1.2715688e-7
+ )

.model pch_mc_8 pmos (
+ level = 49
+ cgso = 3.28e-10
+ nfactor = 1.0
+ a0 = 1.2640158
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ lketa = -5.872592e-10
+ at = 10000.0
+ cf = 0
+ cj = 0.001121
+ ef = 1.064
+ k1 = 0.5203763
+ k2 = 0.04193926
+ k3 = 0.0
+ em = 30000000.0
+ pcdscd = -7.408954e-18
+ js = 2.5e-7
+ ll = 0.0
+ mj = 0.4476
+ lw = 0.0
+ u0 = 0.009795761
+ pb = 0.895226
+ xpart = 1
+ w0 = 0.0
+ rd = 0
+ cjsw = 2.481e-10
+ rs = 0
+ ua = 9.357863e-10
+ ub = 5.091257e-19
+ uc = -1.5731644e-10
+ wl = 0.0
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.007987866
+ pbswg = 0.895226
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ pdiblcb = 0.01
+ pscbe1 = 350000000.0
+ pscbe2 = 5e-7
+ lvoff = 1.6353495e-10
+ tnom = 25.0
+ pags = -6.875222e-16
+ beta0 = 22.67827
+ toxm = 4.08e-9
+ binunit = 2
+ leta0 = 2.5594552000000003e-10
+ letab = -5.545772e-10
+ nqsmod = 0
+ pcit = -7.907631e-17
+ pbsw = 0.895226
+ pclm = 0.9107697
+ tpbswg = 0.001572025
+ lvsat = -0.0003656271
+ noimod = 2
+ lvth0 = -8.128026e-9
+ ppclm = 2.4445072e-15
+ delta = 0.01
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ lcdscd = 3.730414e-11
+ pkt1 = -1.8229216e-15
+ pkt2 = -1.2254391e-15
+ keta = 0.014996022
+ ags = 0.019847063
+ wags = 1.5278273e-9
+ dsub = 0.0
+ version = 3.24
+ cit = -6.09184e-5
+ pketa = -2.4325694e-15
+ dlc = 2e-9
+ lags = 6.882101e-11
+ wcit = 2.0354016e-10
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ k3b = 0.0
+ capmod = 3
+ dwb = 0.0
+ dwg = 0.0
+ wpclm = -5.432238e-9
+ lcit = 1.1752459e-10
+ voff = -0.1308021
+ tcjsw = 0.0004130718
+ ldif = 9e-8
+ kt1l = 0.0
+ prwb = 0.0
+ pub1 = 2.7781507e-32
+ prwg = 0.0
+ puc1 = 8.113434e-24
+ pvoff = -1.9905158e-15
+ eta0 = -0.0004687502
+ mobmod = 1
+ pvag = 0.0
+ etab = 0.0011323938
+ la0 = 5.323636e-9
+ vsat = 130812.52
+ wint = 5e-9
+ pute = 9.798417e-15
+ jsw = 1.2e-12
+ kt1 = -0.2367561
+ lk1 = 1.854804e-8
+ kt2 = -0.025532207
+ lk2 = -6.625426e-9
+ vth0 = -0.449216
+ cdscb = 0.0
+ cdscd = -8.289813e-5
+ pnfactor = 0
+ peta0 = 5.5000000000000005e-21
+ llc = -0.039
+ rdsw = 530.0
+ lln = -1
+ lu0 = -1.2475933e-10
+ petab = 2.4660761e-16
+ wnfactor = 0.0
+ wkt1 = 1.8848993e-8
+ wkt2 = 6.628956e-9
+ lua = -1.759835e-16
+ lub = 1.3507784e-25
+ luc = 1.9437196e-17
+ lint = 1.4999999e-8
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ wmax = 1e-5
+ wketa = 8.724413e-9
+ pvth0 = -1.1241356e-15
+ pa0 = 1.0862038e-13
+ nlx = 0.0
+ wmin = 1.2e-6
+ drout = 0.0
+ lkt1 = -2.4825255e-9
+ lkt2 = -1.0989117e-10
+ tpbsw = 0.001572025
+ pk1 = -1.7383759e-14
+ pk2 = 7.484627e-15
+ lmax = 5e-7
+ pu0 = 2.5785697e-16
+ lmin = 1.8e-7
+ ppdiblc2 = 8.594017e-17
+ prt = 0
+ pua = 1.5976873e-22
+ pub = -1.3085017e-31
+ puc = -9.356197e-24
+ cjswg = 4.221e-10
+ wpdiblc2 = -1.9097854e-10
+ mjswg = 0.3683619
+ lnfactor = 0.0
+ rsh = 7.2
+ tcj = 0.0009739001
+ ua1 = 1.224e-9
+ ub1 = -1.3554493e-18
+ uc1 = 7.051652e-11
+ wvoff = 5.372431e-9
+ tpb = 0.001572025
+ tox = 4.08e-9
+ wub1 = -2.2890885e-25
+ wuc1 = -3.576699e-17
+ wa0 = -4.071248e-7
+ hdif = 2e-7
+ ute = -0.7199521
+ wk1 = 1.1998529e-7
+ wk2 = -4.424634e-8
+ weta0 = 0
+ tcjswg = 0.0004130718
+ lub1 = 2.6058948e-26
+ luc1 = -7.658915e-18
+ wln = 1.0
+ wetab = -5.480169e-10
+ lpdiblc2 = 9.0546e-10
+ wu0 = -2.5725782e-9
+ wute = 1.0915658e-7
+ mjsw = 0.3683619
+ wvsat = 0.0
+ wua = -6.282368e-16
+ wub = 3.0629255e-25
+ wuc = 1.4561782e-17
+ wwl = 0.0
+ wwn = 1.0
+ lpclm = 4.015361e-8
+ wvth0 = 9.142164e-9
+ xti = 3
+ lute = 6.205235e-10
+ cdsc = 0.0
+ wcdscd = 1.6464351e-11
+ cgdo = 3.28e-10
+ )

.model pch_mc_9 pmos (
+ level = 49
+ pvag = 0.0
+ etab = -5e-5
+ lvth0 = 0.0
+ ags = 0.02
+ vsat = 149999.98
+ wint = 5e-9
+ vth0 = -0.4286388
+ delta = 0.01
+ rdsw = 530.0
+ cit = -0.0001
+ wkt1 = 6.74333e-9
+ wkt2 = 1.2948118e-10
+ lint = 1.4999999e-8
+ dlc = 2e-9
+ wmax = 1.2e-6
+ dvt0w = 0.0
+ k3b = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ wmin = 5e-7
+ dwb = 0.0
+ dwg = 0.0
+ lmax = 2.0001e-5
+ lmin = 1e-5
+ capmod = 3
+ a0 = 0.9810578
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ jsw = 1.2e-12
+ kt1 = -0.2307052
+ kt2 = -0.02334808
+ lk2 = 0.0
+ wub1 = 3.495163e-26
+ wuc1 = 1.9335648e-17
+ at = 10000.0
+ cf = 0
+ cj = 0.001121
+ ef = 1.064
+ k1 = 0.5449055
+ k2 = 0.03384938
+ k3 = 0.0
+ em = 30000000.0
+ llc = -0.039
+ lln = -1
+ lu0 = 0.0
+ hdif = 2e-7
+ js = 2.5e-7
+ ll = 0.0
+ mj = 0.4476
+ lw = 0.0
+ u0 = 0.010132165
+ nch = 3.9e+17
+ pb = 0.895226
+ w0 = 0.0
+ rd = 0
+ lwl = 0.0
+ lwn = 1.0
+ rs = 0
+ ua = 1.0698959e-9
+ ub = 3.0837888e-19
+ uc = -1.1659398e-10
+ wl = 0.0
+ wute = -2.7886795e-9
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ mjsw = 0.3683619
+ nlx = 0.0
+ tcjsw = 0.0004130718
+ mobmod = 1
+ pu0 = 0.0
+ pvoff = 0.0
+ prt = 0
+ rsh = 7.2
+ cdscb = 0.0
+ cdscd = 0.0
+ tcj = 0.0009739001
+ peta0 = 5.5000000000000005e-21
+ cdsc = 0.0
+ ua1 = 1.224e-9
+ ub1 = -1.3711068e-18
+ uc1 = 1.6263793e-12
+ tpb = 0.001572025
+ tox = 4.08e-9
+ cgdo = 3.28e-10
+ wketa = -1.0458587e-9
+ wa0 = 3.529885e-8
+ pvth0 = 0.0
+ drout = 0.0
+ ute = -0.7480742
+ wk1 = 2.1990281e-9
+ cgso = 3.28e-10
+ wk2 = -3.824582e-9
+ tpbsw = 0.001572025
+ wln = 1.0
+ wu0 = -2.284236e-10
+ wua = -1.3891575e-16
+ wub = -1.2660565e-25
+ wuc = -3.428342e-17
+ wwl = 0.0
+ wwn = 1.0
+ cjswg = 4.221e-10
+ nfactor = 1.0
+ xti = 3
+ cjsw = 2.481e-10
+ mjswg = 0.3683619
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ wvoff = -4.105241e-10
+ tcjswg = 0.0004130718
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0009999998
+ weta0 = 0
+ tnom = 25.0
+ pdiblcb = 0.01
+ wvsat = 0.0
+ wvth0 = -3.750611e-10
+ toxm = 4.08e-9
+ pbsw = 0.895226
+ pclm = 0.6
+ binunit = 2
+ pnfactor = 0
+ wnfactor = 0.0
+ keta = 0.03217546
+ xpart = 1
+ lnfactor = 0.0
+ alpha0 = 0.0
+ dsub = 0.0
+ alpha1 = 6.8730453846
+ pbswg = 0.895226
+ pscbe1 = 199999970.0
+ pscbe2 = 5e-7
+ dvt0 = 0.0
+ version = 3.24
+ dvt1 = 0.0
+ dvt2 = 0.0
+ lvoff = 0.0
+ voff = -0.12801
+ beta0 = 22.67827
+ nqsmod = 0
+ ldif = 9e-8
+ tpbswg = 0.001572025
+ noimod = 2
+ leta0 = 8e-15
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ eta0 = 5e-5
+ )

.model pch_mc_10 pmos (
+ level = 49
+ dsub = 0.0
+ wk1 = 1.7598129e-9
+ wk2 = -3.600003e-9
+ wln = 1.0
+ wu0 = -1.9812424e-10
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ wua = -1.6455617e-16
+ wub = -7.150721e-26
+ wuc = -2.8652769e-17
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ wwl = 0.0
+ wwn = 1.0
+ xti = 3
+ pscbe1 = 180397680.0
+ pscbe2 = 5e-7
+ voff = -0.1269095
+ ldif = 9e-8
+ nfactor = 1.0
+ kt1l = 0.0
+ prwb = 0.0
+ pub1 = -8.629597e-32
+ prwg = 0.0
+ puc1 = 1.5034668e-23
+ nqsmod = 0
+ tpbswg = 0.001572025
+ lketa = -6.417587e-9
+ eta0 = 5e-5
+ noimod = 2
+ pvag = 0.0
+ etab = -5e-5
+ vsat = 151306.8
+ wint = 5e-9
+ pute = 3.909688e-14
+ xpart = 1
+ vth0 = -0.4245711
+ rdsw = 530.0
+ wkt1 = 6.495125e-9
+ wkt2 = 2.3726165e-10
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0004772722
+ lint = 1.4999999e-8
+ pdiblcb = 0.01
+ lpscbe1 = 195.04263
+ wmax = 1.2e-6
+ pbswg = 0.895226
+ wmin = 5e-7
+ lkt1 = -1.0252924e-8
+ lkt2 = -3.947785e-10
+ lmax = 1e-5
+ lvoff = -1.0948965e-8
+ lmin = 1.2e-6
+ beta0 = 22.67827
+ binunit = 2
+ leta0 = 8e-15
+ lvsat = -0.013002842
+ lvth0 = -4.047293e-8
+ wub1 = 4.362458e-26
+ wuc1 = 1.7824627e-17
+ capmod = 3
+ hdif = 2e-7
+ delta = 0.01
+ lub1 = 7.318341e-26
+ luc1 = 2.7641896e-17
+ pnfactor = 0
+ wute = -6.718015e-9
+ mjsw = 0.3683619
+ wnfactor = 0.0
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ lute = 6.013659e-8
+ mobmod = 1
+ cdsc = 0.0
+ version = 3.24
+ lnfactor = 0.0
+ pketa = -1.6621007e-15
+ cgdo = 3.28e-10
+ ags = 0.02
+ cgso = 3.28e-10
+ cit = -0.0001
+ tcjsw = 0.0004130718
+ dlc = 2e-9
+ lpdiblc2 = 5.201137e-9
+ cjsw = 2.481e-10
+ k3b = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ pvoff = 6.87864e-15
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 5.5000000000000005e-21
+ tcjswg = 0.0004130718
+ tnom = 25.0
+ wketa = -8.788133e-10
+ pvth0 = 1.393327e-14
+ la0 = 1.2176828e-7
+ drout = 0.0
+ toxm = 4.08e-9
+ jsw = 1.2e-12
+ kt1 = -0.2296747
+ lk1 = 1.9542425e-8
+ kt2 = -0.023308404
+ lk2 = -5.136719e-9
+ tpbsw = 0.001572025
+ pbsw = 0.895226
+ llc = -0.039
+ pclm = 0.5738636
+ lln = -1
+ lu0 = -9.551782e-10
+ lua = -5.815077e-16
+ lub = 1.1186816e-24
+ luc = 7.427734e-17
+ nch = 3.9e+17
+ a0 = 0.9688198
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ lwl = 0.0
+ lwn = 1.0
+ cjswg = 4.221e-10
+ at = 10000.0
+ cf = 0
+ cj = 0.001121
+ pa0 = 3.87773e-15
+ nlx = 0.0
+ ef = 1.064
+ k1 = 0.5429414
+ k2 = 0.03436564
+ k3 = 0.0
+ em = 30000000.0
+ mjswg = 0.3683619
+ js = 2.5e-7
+ ll = 0.0
+ mj = 0.4476
+ lw = 0.0
+ pk1 = 4.370194e-15
+ pk2 = -2.2345663e-15
+ u0 = 0.010228163
+ pb = 0.895226
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ua = 1.1283389e-9
+ ub = 1.9594849e-19
+ uc = -1.2405904e-10
+ wvoff = -1.1018445e-9
+ wl = 0.0
+ pu0 = -3.0147877e-16
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ prt = 0
+ pua = 2.5512236e-22
+ pub = -5.482294e-31
+ puc = -5.602498e-23
+ weta0 = 0
+ rsh = 7.2
+ tcj = 0.0009739001
+ ua1 = 1.224e-9
+ ub1 = -1.3784619e-18
+ uc1 = -1.1517035e-12
+ wvsat = 0.0
+ pkt1 = 2.469645e-15
+ pkt2 = -1.0724159e-15
+ keta = 0.03282044
+ tpb = 0.001572025
+ tox = 4.08e-9
+ lpclm = 2.6005682e-7
+ wvth0 = -1.7753915e-9
+ wa0 = 3.490912e-8
+ ute = -0.754118
+ )

.model pch_mc_11 pmos (
+ level = 49
+ cgso = 3.28e-10
+ a0 = 1.1936638
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ lvoff = 5.237211e-9
+ at = 10000.0
+ cf = 0
+ cj = 0.001121
+ ef = 1.064
+ k1 = 0.4715038
+ k2 = 0.05978675
+ k3 = 0.0
+ em = 30000000.0
+ js = 2.5e-7
+ ll = 0.0
+ mj = 0.4476
+ lw = 0.0
+ beta0 = 22.67827
+ u0 = 0.010727104
+ pb = 0.895226
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ua = 1.036115e-9
+ ub = 1.0523674e-18
+ uc = -7.205117e-11
+ cjsw = 2.481e-10
+ leta0 = 3.6972259999999995e-11
+ wl = 0.0
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ letab = -3.696426e-11
+ lvsat = -0.007392855
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ capmod = 3
+ lvth0 = -3.562702e-9
+ delta = 0.01
+ tnom = 25.0
+ ags = 0.02
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ toxm = 4.08e-9
+ mobmod = 1
+ pcit = -1.0851648e-17
+ pbsw = 0.895226
+ pclm = 0.6714286
+ cit = -0.00031597191
+ dlc = 2e-9
+ k3b = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ pketa = 4.024799e-15
+ la0 = -1.3680231e-7
+ pkt1 = -6.051915e-15
+ pkt2 = -1.4802061e-15
+ tcjsw = 0.0004130718
+ keta = 0.03584265
+ jsw = 1.2e-12
+ kt1 = -0.2439705
+ lk1 = 1.0169572e-7
+ kt2 = -0.025852976
+ lk2 = -3.4371e-8
+ llc = -0.039
+ lln = -1
+ lu0 = -1.5289595e-9
+ dsub = 0.0
+ pvoff = -3.866879e-15
+ lua = -4.754501e-16
+ lub = 1.337998e-25
+ luc = 1.4468274e-17
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ pa0 = 1.8891395e-13
+ nlx = 0.0
+ tcjswg = 0.0004130718
+ wcit = 9.436221e-12
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ pk1 = -6.35241e-14
+ pk2 = 2.2224691e-14
+ peta0 = 5.5000000000000005e-21
+ pu0 = 7.878928e-16
+ pnfactor = 0
+ prt = 0
+ lcit = 2.4836766e-10
+ pua = 2.5287059e-22
+ pub = -5.865131e-32
+ puc = -1.2704817e-23
+ wketa = -5.823942e-9
+ voff = -0.1409845
+ pvth0 = -5.102908e-15
+ wnfactor = 0.0
+ ldif = 9e-8
+ drout = 0.0
+ kt1l = 0.0
+ tpbsw = 0.001572025
+ prwb = 0.0
+ pub1 = 4.97241e-32
+ prwg = 0.0
+ rsh = 7.2
+ puc1 = 1.7282469e-23
+ tcj = 0.0009739001
+ ua1 = 1.224e-9
+ ub1 = -1.2162624e-18
+ uc1 = 4.210797e-11
+ eta0 = 1.7857154e-5
+ nfactor = 1.0
+ pvag = 0.0
+ etab = -1.7857154e-5
+ tpb = 0.001572025
+ tox = 4.08e-9
+ cjswg = 4.221e-10
+ vsat = 146428.56
+ wa0 = -1.2599192e-7
+ wint = 5e-9
+ pute = -5.928695e-14
+ mjswg = 0.3683619
+ vth0 = -0.456667
+ ute = -0.7903757
+ wk1 = 6.079834e-8
+ wk2 = -2.4868919e-8
+ rdsw = 530.0
+ wln = 1.0
+ wkt1 = 1.3905176e-8
+ wkt2 = 5.918618e-10
+ lnfactor = 0.0
+ wu0 = -1.1454039e-9
+ lint = 1.4999999e-8
+ wvoff = 8.242083e-9
+ wua = -1.625981e-16
+ wmax = 1.2e-6
+ wub = -4.972273e-25
+ wuc = -6.632247e-17
+ wwl = 0.0
+ wwn = 1.0
+ wmin = 5e-7
+ xti = 3
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0017857137
+ lkt1 = 6.187276e-9
+ lkt2 = 2.5314804e-9
+ pdiblcb = 0.01
+ weta0 = 0
+ lmax = 1.2e-6
+ lmin = 5e-7
+ wvsat = 0.0
+ lpclm = 1.4785714e-7
+ wvth0 = 1.4777807e-8
+ lpdiblc2 = 3.696429e-9
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ binunit = 2
+ pscbe1 = 349999900.0
+ pscbe2 = 5e-7
+ wub1 = -7.465372e-26
+ wuc1 = 1.5870021e-17
+ hdif = 2e-7
+ lub1 = -1.133461e-25
+ luc1 = -2.2106738e-17
+ wute = 7.883313e-8
+ mjsw = 0.3683619
+ nqsmod = 0
+ tpbswg = 0.001572025
+ noimod = 2
+ lute = 1.0183292e-7
+ lketa = -9.893122e-9
+ xpart = 1
+ cdsc = 0.0
+ cgdo = 3.28e-10
+ pbswg = 0.895226
+ version = 3.24
+ )

.model pch_mc_12 pmos (
+ level = 49
+ wint = 5e-9
+ llc = -0.039
+ pute = 1.3160581e-15
+ lln = -1
+ lu0 = 2.1198607e-10
+ vth0 = -0.4463558
+ nfactor = 1.0
+ lua = 2.3815556e-17
+ lub = -3.425063e-26
+ luc = 8.803578e-18
+ nch = 3.9e+17
+ rdsw = 530.0
+ lwl = 0.0
+ lwn = 1.0
+ pketa = -9.609158e-16
+ wkt1 = 2.7434011e-10
+ wkt2 = -6.113567e-9
+ lint = 1.4999999e-8
+ pa0 = -8.476619e-14
+ nlx = 0.0
+ wmax = 1.2e-6
+ pk1 = 1.5213101e-14
+ pk2 = -6.235986e-15
+ wmin = 5e-7
+ lkt1 = -4.083267e-9
+ lkt2 = -2.4314675e-9
+ wpclm = 5.671285e-8
+ pu0 = -1.4287007e-16
+ lmax = 5e-7
+ prt = 0
+ pua = -7.799214e-23
+ pub = 7.065072e-32
+ puc = 3.297807e-24
+ lmin = 1.8e-7
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.009150297
+ tcjsw = 0.0004130718
+ pdiblcb = 0.01
+ rsh = 7.2
+ tcj = 0.0009739001
+ ua1 = 1.224e-9
+ ub1 = -1.6175756e-18
+ uc1 = -2.2818641e-11
+ pvoff = -1.4343533e-15
+ tcjswg = 0.0004130718
+ tpb = 0.001572025
+ tox = 4.08e-9
+ a0 = 0.5166956
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ wa0 = 4.821862e-7
+ at = 10000.0
+ cf = 0
+ cj = 0.001121
+ wub1 = 8.30214e-26
+ ute = -0.5812994
+ wuc1 = 7.530186e-17
+ ef = 1.064
+ k1 = 0.7171482
+ k2 = -0.027492139
+ k3 = 0.0
+ em = 30000000.0
+ wk1 = -1.1417325e-7
+ wk2 = 3.837703e-8
+ binunit = 2
+ cdscb = 0.0
+ cdscd = -5.200001e-5
+ peta0 = 5.5000000000000005e-21
+ js = 2.5e-7
+ ll = 0.0
+ mj = 0.4476
+ hdif = 2e-7
+ lw = 0.0
+ u0 = 0.006858335
+ wln = 1.0
+ pb = 0.895226
+ w0 = 0.0
+ wu0 = 9.229584e-10
+ rd = 0
+ rs = 0
+ ua = -7.336427e-11
+ ub = 1.4258127e-18
+ uc = -5.946296e-11
+ lub1 = 6.724484e-26
+ wua = 5.726523e-16
+ wub = -7.845651e-25
+ wuc = -1.0188386e-16
+ wl = 0.0
+ luc1 = 7.110234e-18
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ wwl = 0.0
+ wwn = 1.0
+ wute = -5.584022e-8
+ wketa = 5.255423e-9
+ mjsw = 0.3683619
+ pvth0 = -1.0352502e-15
+ xti = 3
+ drout = 0.0
+ tpbsw = 0.001572025
+ lute = 7.748556e-9
+ wcdscd = -2.0304376e-11
+ cjswg = 4.221e-10
+ mjswg = 0.3683619
+ cdsc = 0.0
+ wvoff = 2.8364715e-9
+ cgdo = 3.28e-10
+ pcdscd = 9.13697e-18
+ cgso = 3.28e-10
+ weta0 = 0
+ version = 3.24
+ wvsat = 0.0
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ lpclm = 6.365384e-8
+ wvth0 = 5.738565e-9
+ cjsw = 2.481e-10
+ pscbe1 = 350000000.0
+ pscbe2 = 5e-7
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ nqsmod = 0
+ tpbswg = 0.001572025
+ tnom = 25.0
+ pnfactor = 0
+ noimod = 2
+ pags = -5.667374e-15
+ wnfactor = 0.0
+ toxm = 4.08e-9
+ pcit = 2.6834248e-18
+ pbsw = 0.895226
+ lketa = -1.8239428e-9
+ pclm = 0.858547
+ xpart = 1
+ ppdiblc2 = 7.08422e-16
+ wpdiblc2 = -1.5742713e-9
+ lnfactor = 0.0
+ pbswg = 0.895226
+ lcdscd = 2.3400004e-11
+ lvoff = -3.0382863e-10
+ ags = 0.010547621
+ beta0 = 22.67827
+ pkt1 = 8.196091e-17
+ pkt2 = 1.5372367e-15
+ keta = 0.01791114
+ lpdiblc2 = 3.823661e-10
+ leta0 = 2.5594547e-10
+ capmod = 3
+ letab = -3.473438e-10
+ cit = 0.00012746976
+ wags = 1.2594167e-8
+ lvsat = -0.0003656142
+ dsub = 0.0
+ dlc = 2e-9
+ lvth0 = -8.202719e-9
+ k3b = 0.0
+ dwb = 0.0
+ dwg = 0.0
+ lags = 4.253569e-9
+ wcit = -2.0641719e-11
+ ppclm = -2.5520774e-14
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ delta = 0.01
+ mobmod = 1
+ lcit = 4.881893e-11
+ voff = -0.1286711
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ ldif = 9e-8
+ kt1l = 0.0
+ prwb = 0.0
+ pub1 = -2.1229706e-32
+ prwg = 0.0
+ puc1 = -9.461855e-24
+ la0 = 1.6783336e-7
+ eta0 = -0.00046875
+ pvag = 0.0
+ jsw = 1.2e-12
+ etab = 0.0006718753
+ kt1 = -0.2211471
+ lk1 = -8.844278e-9
+ kt2 = -0.014824204
+ lk2 = 4.904499e-9
+ vsat = 130812.46
+ )

.model pch_mc_13 pmos (
+ level = 49
+ wketa = -6.403492e-9
+ pvth0 = 0.0
+ drout = 0.0
+ toxm = 4.08e-9
+ tpbsw = 0.001572025
+ pbsw = 0.895226
+ pclm = 0.5999999
+ cjswg = 4.221e-10
+ mjswg = 0.3683619
+ wvoff = -1.320298e-9
+ weta0 = 0
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ wvsat = 0.0
+ keta = 0.04310941
+ pscbe1 = 199999970.0
+ pscbe2 = 5e-7
+ wvth0 = 9.340613e-9
+ dsub = 0.0
+ nqsmod = 0
+ tpbswg = 0.001572025
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ noimod = 2
+ voff = -0.1261533
+ ldif = 9e-8
+ a0 = 0.8704194
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ kt1l = 0.0
+ prwb = 0.0
+ prwg = 0.0
+ at = 10000.0
+ cf = 0
+ cj = 0.001121
+ ef = 1.064
+ k1 = 0.5421249
+ k2 = 0.03567642
+ k3 = 0.0
+ em = 30000000.0
+ ags = 0.02
+ eta0 = 5e-5
+ js = 2.5e-7
+ ll = 0.0
+ mj = 0.4476
+ lw = 0.0
+ pvag = 0.0
+ etab = -5e-5
+ u0 = 0.009748334
+ pb = 0.895226
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ vsat = 149999.98
+ xpart = 1
+ ua = 1.2584637e-9
+ ub = 4.999999e-20
+ uc = -1.6065008e-10
+ wint = 5e-9
+ wl = 0.0
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ cit = -0.0001
+ vth0 = -0.4484667
+ rdsw = 530.0
+ dlc = 2e-9
+ wkt1 = 3.830554e-9
+ wkt2 = 1.9527771e-9
+ k3b = 0.0
+ lint = 1.4999999e-8
+ pbswg = 0.895226
+ dwb = 0.0
+ wmax = 5e-7
+ dwg = 0.0
+ nfactor = 1.0
+ wmin = 2.2e-7
+ lvoff = 0.0
+ lmax = 2.0001e-5
+ lmin = 1e-5
+ capmod = 3
+ beta0 = 22.67827
+ leta0 = 8e-15
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.001
+ pdiblcb = 0.01
+ jsw = 1.2e-12
+ kt1 = -0.2247607
+ kt2 = -0.027069092
+ lk2 = 0.0
+ lvth0 = 0.0
+ llc = -0.039
+ lln = -1
+ lu0 = 0.0
+ wub1 = 2.1644123e-27
+ wuc1 = -1.2526765e-17
+ nch = 3.9e+17
+ mobmod = 1
+ lwl = 0.0
+ lwn = 1.0
+ delta = 0.01
+ hdif = 2e-7
+ nlx = 0.0
+ pnfactor = 0
+ binunit = 2
+ wute = 6.898109e-9
+ mjsw = 0.3683619
+ wnfactor = 0.0
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ pu0 = 0.0
+ prt = 0
+ rsh = 7.2
+ tcj = 0.0009739001
+ ua1 = 1.224e-9
+ ub1 = -1.3041941e-18
+ uc1 = 6.665171e-11
+ cdsc = 0.0
+ tpb = 0.001572025
+ tox = 4.08e-9
+ wa0 = 8.951166e-8
+ lnfactor = 0.0
+ cgdo = 3.28e-10
+ ute = -0.7678431
+ wk1 = 3.561511e-9
+ wk2 = -4.719829e-9
+ wln = 1.0
+ cgso = 3.28e-10
+ wu0 = -4.034686e-11
+ wua = -2.3131395e-16
+ wuc = -1.2695932e-17
+ wwl = 0.0
+ wwn = 1.0
+ xti = 3
+ tcjsw = 0.0004130718
+ tcjswg = 0.0004130718
+ version = 3.24
+ cjsw = 2.481e-10
+ pvoff = 0.0
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 5.5000000000000005e-21
+ tnom = 25.0
+ )

.model pch_mc_14 pmos (
+ level = 49
+ tpbswg = 0.001572025
+ noimod = 2
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0004772729
+ cit = -0.0001
+ wub1 = -3.0198158e-27
+ wuc1 = -1.0513175e-17
+ pdiblcb = 0.01
+ lpscbe1 = 195.04262
+ dlc = 2e-9
+ hdif = 2e-7
+ k3b = 0.0
+ lub1 = -2.0820251e-25
+ dwb = 0.0
+ dwg = 0.0
+ luc1 = 9.921307e-17
+ wute = 1.1298283e-8
+ mjsw = 0.3683619
+ binunit = 2
+ lketa = -4.562476e-8
+ lute = 2.2927659e-7
+ xpart = 1
+ la0 = 5.081137e-7
+ cdsc = 0.0
+ jsw = 1.2e-12
+ kt1 = -0.2237138
+ lk1 = -4.88067e-8
+ kt2 = -0.026908273
+ lk2 = 2.3302198e-8
+ llc = -0.039
+ lln = -1
+ cgdo = 3.28e-10
+ lu0 = -3.0000519e-10
+ pbswg = 0.895226
+ lua = -3.24011e-17
+ lub = -3.941427e-28
+ luc = -6.882293e-17
+ nch = 3.9e+17
+ lwl = 0.0
+ lwn = 1.0
+ cgso = 3.28e-10
+ pa0 = -1.854315e-13
+ lvoff = -2.3886029e-9
+ nlx = 0.0
+ capmod = 3
+ pk1 = 3.786126e-14
+ pk2 = -1.6169635e-14
+ beta0 = 22.67827
+ pu0 = -6.225135e-16
+ leta0 = 8e-15
+ prt = 0
+ pua = -1.3939852e-23
+ pub = 1.1764949e-34
+ puc = 1.4094153e-23
+ cjsw = 2.481e-10
+ lvsat = -0.013002842
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ lvth0 = -4.608335e-9
+ version = 3.24
+ rsh = 7.2
+ tcj = 0.0009739001
+ mobmod = 1
+ ua1 = 1.224e-9
+ ub1 = -1.2832692e-18
+ uc1 = 5.668055e-11
+ tpb = 0.001572025
+ tox = 4.08e-9
+ delta = 0.01
+ wa0 = 1.0814799e-7
+ tnom = 25.0
+ ute = -0.790886
+ wk1 = -2.4364055e-10
+ wk2 = -3.0947396e-9
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ wln = 1.0
+ wu0 = 2.2217313e-11
+ toxm = 4.08e-9
+ wua = -2.2991296e-16
+ wub = -1.1822094e-29
+ wuc = -1.4112429e-17
+ wwl = 0.0
+ wwn = 1.0
+ pbsw = 0.895226
+ xti = 3
+ pclm = 0.5738635
+ pketa = 1.7549415e-14
+ a0 = 0.8193527
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ at = 10000.0
+ cf = 0
+ cj = 0.001121
+ ef = 1.064
+ k1 = 0.5470301
+ k2 = 0.03333449
+ k3 = 0.0
+ em = 30000000.0
+ js = 2.5e-7
+ ll = 0.0
+ mj = 0.4476
+ lw = 0.0
+ u0 = 0.009778486
+ pb = 0.895226
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ua = 1.2617201e-9
+ ub = 5.00396e-20
+ uc = -1.5373321e-10
+ wl = 0.0
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -2e-8
+ ww = 0.0
+ tcjswg = 0.0004130718
+ xw = 0.0
+ tcjsw = 0.0004130718
+ pkt1 = 2.5501714e-15
+ pkt2 = -4.817884e-16
+ keta = 0.04769481
+ pvoff = 2.6840621e-15
+ dsub = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ peta0 = 5.5000000000000005e-21
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ pnfactor = 0
+ wketa = -8.167253e-9
+ pvth0 = -3.640382e-15
+ wnfactor = 0.0
+ voff = -0.1259132
+ drout = 0.0
+ ldif = 9e-8
+ tpbsw = 0.001572025
+ kt1l = 0.0
+ prwb = 0.0
+ pub1 = 5.158311e-32
+ prwg = 0.0
+ puc1 = -2.0035212e-23
+ eta0 = 5e-5
+ cjswg = 4.221e-10
+ pvag = 0.0
+ etab = -5e-5
+ vsat = 151306.8
+ mjswg = 0.3683619
+ wint = 5e-9
+ pute = -4.378173e-14
+ vth0 = -0.4480035
+ rdsw = 530.0
+ lnfactor = 0.0
+ wvoff = -1.590053e-9
+ wkt1 = 3.574256e-9
+ wkt2 = 2.0011981e-9
+ lint = 1.4999999e-8
+ wmax = 5e-7
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ wmin = 2.2e-7
+ lkt1 = -1.0417262e-8
+ lkt2 = -1.6001408e-9
+ weta0 = 0
+ nfactor = 1.0
+ lmax = 1e-5
+ pscbe1 = 180397700.0
+ pscbe2 = 5e-7
+ wvsat = 0.0
+ lmin = 1.2e-6
+ lpclm = 2.6005691e-7
+ wvth0 = 9.70648e-9
+ lpdiblc2 = 5.201136e-9
+ ags = 0.02
+ nqsmod = 0
+ )

.model pch_mc_15 pmos (
+ level = 49
+ ute = -0.5904401
+ wk1 = 4.182789e-8
+ wk2 = -2.2085489e-8
+ beta0 = 22.67827
+ wln = 1.0
+ wu0 = -3.987341e-10
+ pkt1 = -8.599671e-15
+ pkt2 = 1.9347028e-16
+ lpdiblc2 = 3.696429e-9
+ keta = 0.0004484208
+ wua = -1.9008923e-16
+ leta0 = 3.697228e-11
+ wub = 8.369847e-27
+ wuc = 5.370726e-18
+ wwl = 0.0
+ wwn = 1.0
+ letab = -3.696428e-11
+ xti = 3
+ mobmod = 1
+ lvsat = -0.007392816
+ dsub = 0.0
+ lvth0 = -1.5532533e-8
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ delta = 0.01
+ lcit = 2.2622144e-10
+ dvt0w = 0.0
+ dvt1w = 0.0
+ dvt2w = 0.0
+ voff = -0.1186655
+ ldif = 9e-8
+ kt1l = 0.0
+ prwb = 0.0
+ pub1 = -1.2589071e-33
+ prwg = 0.0
+ puc1 = 4.27717e-24
+ eta0 = 1.7857146e-5
+ pvag = 0.0
+ etab = -1.7857146e-5
+ vsat = 146428.52
+ wint = 5e-9
+ pute = -8.783067e-15
+ vth0 = -0.4385042
+ rdsw = 530.0
+ pketa = -5.090041e-15
+ wkt1 = 1.3269771e-8
+ wkt2 = 1.4140165e-9
+ lint = 1.4999999e-8
+ wmax = 5e-7
+ tcjswg = 0.0004130718
+ wmin = 2.2e-7
+ lkt1 = 1.1386779e-8
+ lkt2 = -8.841858e-10
+ lmax = 1.2e-6
+ lmin = 5e-7
+ tcjsw = 0.0004130718
+ nfactor = 1.0
+ pvoff = 3.95383e-15
+ wub1 = 4.292976e-26
+ cdscb = 0.0
+ wuc1 = -3.165437e-17
+ cdscd = 0.0
+ peta0 = 5.5000000000000005e-21
+ hdif = 2e-7
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.0017857139
+ pdiblcb = 0.01
+ lub1 = -9.299159e-27
+ wketa = 1.1519229e-8
+ luc1 = 4.434689e-18
+ pvth0 = 7.623086e-16
+ wute = -1.9135335e-8
+ mjsw = 0.3683619
+ drout = 0.0
+ tpbsw = 0.001572025
+ lute = -1.2362289e-9
+ cjswg = 4.221e-10
+ binunit = 2
+ mjswg = 0.3683619
+ ags = 0.02
+ cdsc = 0.0
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ wvoff = -2.6941984e-9
+ cit = -0.00029671428
+ cgdo = 3.28e-10
+ pscbe1 = 349999900.0
+ pscbe2 = 5e-7
+ dlc = 2e-9
+ cgso = 3.28e-10
+ k3b = 0.0
+ weta0 = 0
+ dwb = 0.0
+ dwg = 0.0
+ wvsat = 0.0
+ lpclm = 1.4785714e-7
+ wvth0 = 5.878054e-9
+ nqsmod = 0
+ a0 = 1.1508681
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ tpbswg = 0.001572025
+ cjsw = 2.481e-10
+ noimod = 2
+ at = 10000.0
+ cf = 0
+ cj = 0.001121
+ ef = 1.064
+ k1 = 0.510219
+ k2 = 0.05410628
+ k3 = 0.0
+ em = 30000000.0
+ js = 2.5e-7
+ ll = 0.0
+ noia = 9.5e+18
+ mj = 0.4476
+ noib = 100000.0
+ noic = 1.4e-12
+ lw = 0.0
+ u0 = 0.009203287
+ pb = 0.895226
+ w0 = 0.0
+ rd = 0
+ rs = 0
+ ua = 1.0922192e-9
+ ub = 2.0536515e-20
+ uc = -2.183638e-10
+ la0 = 1.2687106e-7
+ wl = 0.0
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -2e-8
+ ww = 0.0
+ xw = 0.0
+ jsw = 1.2e-12
+ version = 3.24
+ kt1 = -0.2426738
+ lk1 = -6.473878e-9
+ kt2 = -0.027530843
+ lk2 = -5.853628e-10
+ llc = -0.039
+ lln = -1
+ pnfactor = 0
+ lu0 = 3.614737e-10
+ tnom = 25.0
+ lua = 1.6252487e-16
+ lub = 3.353441e-26
+ luc = 5.502275e-18
+ nch = 3.9e+17
+ wnfactor = 0.0
+ lwl = 0.0
+ lwn = 1.0
+ pa0 = 5.971399e-14
+ nlx = 0.0
+ toxm = 4.08e-9
+ lketa = 8.708591e-9
+ pk1 = -1.0521005e-14
+ pk2 = 5.669729e-15
+ pbsw = 0.895226
+ pclm = 0.6714286
+ pu0 = -1.384194e-16
+ xpart = 1
+ prt = 0
+ pua = -5.973716e-23
+ pub = -9.521269e-33
+ puc = -8.311478e-24
+ rsh = 7.2
+ lnfactor = 0.0
+ tcj = 0.0009739001
+ ua1 = 1.224e-9
+ ub1 = -1.4562286e-18
+ uc1 = 1.3909653e-10
+ pbswg = 0.895226
+ capmod = 3
+ tpb = 0.001572025
+ tox = 4.08e-9
+ wa0 = -1.0502199e-7
+ lvoff = -1.0723419e-8
+ )

.model pch_mc_16 pmos (
+ level = 49
+ cdsc = 0.0
+ binunit = 2
+ pketa = 7.45672e-16
+ lnfactor = 0.0
+ tcjswg = 0.0004130718
+ cgdo = 3.28e-10
+ wpclm = 4.634222e-9
+ cgso = 3.28e-10
+ tcjsw = 0.0004130718
+ lpdiblc2 = 1.8281252e-9
+ cjsw = 2.481e-10
+ pvoff = 1.4541431e-15
+ noia = 9.5e+18
+ noib = 100000.0
+ noic = 1.4e-12
+ wcdscd = -1.4183201e-11
+ ags = 0.03625
+ cdscb = 0.0
+ cdscd = -6.449223e-5
+ peta0 = 5.5000000000000005e-21
+ cit = 8.534377e-5
+ tnom = 25.0
+ wketa = -1.4490222e-9
+ pvth0 = -2.8414808e-16
+ version = 3.24
+ dlc = 2e-9
+ drout = 0.0
+ pcdscd = 6.382441e-18
+ tpbsw = 0.001572025
+ k3b = 0.0
+ toxm = 4.08e-9
+ dwb = 0.0
+ dwg = 0.0
+ pbsw = 0.895226
+ pclm = 0.9648299
+ cjswg = 4.221e-10
+ mjswg = 0.3683619
+ alpha0 = 0.0
+ alpha1 = 6.8730453846
+ wvoff = 2.8606606e-9
+ pscbe1 = 350000000.0
+ pscbe2 = 5e-7
+ la0 = 7.233052e-9
+ jsw = 1.2e-12
+ kt1 = -0.2130934
+ lk1 = 1.3789155e-8
+ kt2 = -0.03589084
+ lk2 = -3.106946e-9
+ llc = -0.039
+ weta0 = 0
+ lln = -1
+ lu0 = -3.566262e-10
+ nqsmod = 0
+ lua = -2.6402067e-16
+ lub = 2.6345733e-25
+ luc = 3.340897e-17
+ nch = 3.9e+17
+ wvsat = 0.0
+ tpbswg = 0.001572025
+ lwl = 0.0
+ lwn = 1.0
+ noimod = 2
+ lpclm = 1.5826547e-8
+ pa0 = -6.072043e-15
+ wvth0 = 8.203513e-9
+ nlx = 0.0
+ pkt1 = -9.758805e-16
+ pkt2 = -1.0643102e-15
+ keta = 0.03159368
+ pk1 = 4.122718e-15
+ pk2 = -2.3103772e-15
+ dsub = 0.0
+ pu0 = 1.3574996e-16
+ prt = 0
+ pua = 6.304761e-23
+ pub = -7.522618e-32
+ puc = -8.758834e-24
+ lags = -7.312499e-9
+ dvt0 = 0.0
+ dvt1 = 0.0
+ dvt2 = 0.0
+ rsh = 7.2
+ tcj = 0.0009739001
+ ua1 = 1.224e-9
+ ub1 = -1.4433942e-18
+ uc1 = 2.0396977e-10
+ tpb = 0.001572025
+ tox = 4.08e-9
+ lcit = 5.429531e-11
+ voff = -0.1287204
+ wa0 = 4.116919e-8
+ lcdscd = 2.9021494e-11
+ ldif = 9e-8
+ ute = -0.5893072
+ wk1 = 9.286284e-9
+ kt1l = 0.0
+ wk2 = -4.351921e-9
+ prwb = 0.0
+ pub1 = 1.9106841e-32
+ prwg = 0.0
+ lketa = -5.306775e-9
+ puc1 = 6.153712e-24
+ wln = 1.0
+ wu0 = -1.0079994e-9
+ eta0 = -0.0004687502
+ wua = -4.629443e-16
+ pvag = 0.0
+ wub = 1.5438073e-25
+ wuc = 6.364847e-18
+ etab = 0.0006718753
+ xpart = 1
+ wwl = 0.0
+ wwn = 1.0
+ vsat = 130812.55
+ xti = 3
+ wint = 5e-9
+ pute = 5.968411e-15
+ vth0 = -0.4513863
+ capmod = 3
+ rdsw = 530.0
+ wkt1 = -3.671987e-9
+ wkt2 = 4.209085e-9
+ pbswg = 0.895226
+ lint = 1.4999999e-8
+ wmax = 5e-7
+ wmin = 2.2e-7
+ lvoff = -6.198719e-9
+ lkt1 = -1.9244071e-9
+ lkt2 = 2.877812e-9
+ lmax = 5e-7
+ beta0 = 22.67827
+ lmin = 1.8e-7
+ mobmod = 1
+ leta0 = 2.5594558000000004e-10
+ letab = -3.473438e-10
+ lvsat = -0.0003656336
+ nfactor = 1.0
+ lvth0 = -9.735581e-9
+ ppclm = -2.0853998e-15
+ wub1 = -2.3274574e-27
+ wuc1 = -3.582447e-17
+ delta = 0.01
+ hdif = 2e-7
+ a0 = 1.4167303
+ a1 = 0.0
+ a2 = 0.4
+ b0 = 0.0
+ b1 = 0.0
+ pnfactor = 0
+ lub1 = -1.5074642e-26
+ luc1 = -2.4758267e-17
+ at = 10000.0
+ cf = 0
+ cj = 0.001121
+ ef = 1.064
+ k1 = 0.46519
+ dvt0w = 0.0
+ k2 = 0.0597098
+ k3 = 0.0
+ em = 30000000.0
+ wnfactor = 0.0
+ wute = -5.191639e-8
+ dvt1w = 0.0
+ dvt2w = 0.0
+ mjsw = 0.3683619
+ js = 2.5e-7
+ pdiblc1 = 1e-6
+ pdiblc2 = 0.005937499
+ ll = 0.0
+ mj = 0.4476
+ lw = 0.0
+ u0 = 0.010799064
+ pb = 0.895226
+ w0 = 0.0
+ rd = 0
+ pdiblcb = 0.01
+ rs = 0
+ ua = 2.0400983e-9
+ ub = -4.904033e-19
+ uc = -2.8037866e-10
+ wl = 0.0
+ wr = 1.0
+ xj = 1.7000001e-7
+ xl = -2e-8
+ ww = 0.0
+ lute = -1.7460413e-9
+ xw = 0.0
+ )

